chr5	1192522	+	chr5	1191303	+	.	24	0	3147401_1	42.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=3147401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:1191303(-)-5:1192522(+)__5_1176001_1201001D;SPAN=1219;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:135 GQ:42.8 PL:[42.8, 0.0, 283.7] SR:0 DR:24 LR:-42.65 LO:53.02);ALT=]chr5:1192522]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1465909	+	chr5	1464635	+	.	39	3	3148990_1	50.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TGCACACTTTCAA;MAPQ=60;MATEID=3148990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_1445501_1470501_20C;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:42 DP:325 GQ:50.7 PL:[50.7, 0.0, 737.3] SR:3 DR:39 LR:-50.59 LO:86.42);ALT=]chr5:1465909]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1968413	+	chr5	1971584	+	.	98	40	3152303_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAATAAAGAAAATTGTGG;MAPQ=60;MATEID=3152303_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_1960001_1985001_366C;SPAN=3171;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:135 DP:326 GQ:99 PL:[357.4, 0.0, 433.3] SR:40 DR:98 LR:-357.3 LO:357.7);ALT=G[chr5:1971584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	2138484	-	chr14	76733257	+	.	3	17	3153906_1	47.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCTTTCCTTTCCTTTCCTTTCCTTTC;MAPQ=60;MATEID=3153906_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_2131501_2156501_536C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:30 GQ:24.8 PL:[47.9, 0.0, 24.8] SR:17 DR:3 LR:-48.39 LO:48.39);ALT=[chr14:76733257[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	77304244	-	chr14	77310625	+	.	90	88	8618214_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=8618214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_77297501_77322501_462C;SPAN=6381;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:155 DP:210 GQ:55.3 PL:[454.7, 0.0, 55.3] SR:88 DR:90 LR:-473.0 LO:473.0);ALT=[chr14:77310625[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
