chr5	159263388	+	chr5	159275383	+	ACATGCATATA	0	37	3880572_1	99.0	.	EVDNC=ASSMB;INSERTION=ACATGCATATA;MAPQ=60;MATEID=3880572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_159274501_159299501_105C;SPAN=11995;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:52 GQ:15.8 PL:[108.2, 0.0, 15.8] SR:37 DR:0 LR:-111.7 LO:111.7);ALT=T[chr5:159275383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	159444293	+	chr5	159445305	-	.	0	4	3881079_1	0	.	EVDNC=ASSMB;HOMSEQ=AATAAATTTCTATTATTTATAA;MAPQ=60;MATEID=3881079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_159421501_159446501_59C;SPAN=1012;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:126 GQ:20.7 PL:[0.0, 20.7, 346.5] SR:4 DR:0 LR:20.93 LO:5.71);ALT=T]chr5:159445305];VARTYPE=BND:INV-hh;JOINTYPE=hh
