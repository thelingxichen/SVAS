chr21	26934569	+	chr21	26942146	+	.	6	4	7142329_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7142329_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_26925501_26950501_20C;SPAN=7577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:4 DR:6 LR:-7.543 LO:19.68);ALT=G[chr21:26942146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	26934573	+	chr21	26946202	+	.	10	0	7142330_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7142330_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:26934573(+)-21:26946202(-)__21_26925501_26950501D;SPAN=11629;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:0 DR:10 LR:-10.79 LO:20.31);ALT=C[chr21:26946202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	26942235	+	chr21	26946204	+	.	0	11	7142349_1	13.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7142349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_26925501_26950501_106C;SPAN=3969;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:11 DR:0 LR:-13.28 LO:22.64);ALT=T[chr21:26946204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	27097661	+	chr21	27101941	+	.	0	59	7142832_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7142832_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_27097001_27122001_92C;SPAN=4280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:93 GQ:54.2 PL:[169.7, 0.0, 54.2] SR:59 DR:0 LR:-172.7 LO:172.7);ALT=C[chr21:27101941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	27097701	+	chr21	27107163	+	.	28	0	7142834_1	57.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7142834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:27097701(+)-21:27107163(-)__21_27097001_27122001D;SPAN=9462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:130 GQ:57.2 PL:[57.2, 0.0, 258.5] SR:0 DR:28 LR:-57.21 LO:64.48);ALT=C[chr21:27107163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	27102152	+	chr21	27107162	+	.	57	0	7142842_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7142842_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:27102152(+)-21:27107162(-)__21_27097001_27122001D;SPAN=5010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:129 GQ:99 PL:[153.2, 0.0, 159.8] SR:0 DR:57 LR:-153.2 LO:153.2);ALT=A[chr21:27107162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	28020683	-	chr21	28021726	+	.	33	23	7145479_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7145479_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_21_28003501_28028501_205C;SECONDARY;SPAN=1043;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:78 GQ:41.6 PL:[147.2, 0.0, 41.6] SR:23 DR:33 LR:-150.5 LO:150.5);ALT=[chr21:28021726[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
