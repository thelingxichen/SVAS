chrX	152506377	-	chrX	152634502	+	.	17	21	11428835_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=GCCACCACACCTGGCTAATTTTTTTGTATTTTTAGTAGAGA;MAPQ=57;MATEID=11428835_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=AGAG;SCTG=c_23_152610501_152635501_22C;SECONDARY;SPAN=128125;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:38 DP:23 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:21 DR:17 LR:-112.2 LO:112.2);ALT=[chrX:152634502[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
