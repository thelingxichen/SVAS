chr2	130940026	+	chr2	130948042	+	.	22	12	993241_1	61.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=993241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_130928001_130953001_6C;SPAN=8016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:141 GQ:61.1 PL:[61.1, 0.0, 278.9] SR:12 DR:22 LR:-60.83 LO:68.9);ALT=G[chr2:130948042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	130954939	+	chr2	130957404	+	.	26	22	993387_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=CACACCTGTA;MAPQ=23;MATEID=993387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_130952501_130977501_7C;SPAN=2465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:63 GQ:39.2 PL:[111.8, 0.0, 39.2] SR:22 DR:26 LR:-113.4 LO:113.4);ALT=A[chr2:130957404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	131100573	+	chr2	131102946	+	.	11	0	993676_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=993676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:131100573(+)-2:131102946(-)__2_131099501_131124501D;SPAN=2373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:0 DR:11 LR:-11.39 LO:22.24);ALT=G[chr2:131102946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	131100767	+	chr2	131102200	+	.	5	29	993680_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=993680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_131099501_131124501_303C;SPAN=1433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:101 GQ:85.1 PL:[85.1, 0.0, 157.7] SR:29 DR:5 LR:-84.87 LO:86.14);ALT=G[chr2:131102200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
