chr5	117096153	+	chr5	117260703	+	.	12	0	2562621_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2562621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:117096153(+)-5:117260703(-)__5_117257001_117282001D;SPAN=164550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:19 GQ:11.3 PL:[34.4, 0.0, 11.3] SR:0 DR:12 LR:-35.09 LO:35.09);ALT=T[chr5:117260703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
