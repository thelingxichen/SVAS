chr13	65342433	+	chr13	65344424	+	.	33	31	5532172_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATTTTT;MAPQ=60;MATEID=5532172_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_13_65341501_65366501_267C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:48 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:31 DR:33 LR:-148.5 LO:148.5);ALT=T[chr13:65344424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
