chr10	132909062	+	chr10	132912780	+	.	114	46	6607370_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTCA;MAPQ=60;MATEID=6607370_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_132912501_132937501_193C;SPAN=3718;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:141 DP:16 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:46 DR:114 LR:-415.9 LO:415.9);ALT=A[chr10:132912780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	133522773	+	chr10	133519935	+	.	8	0	6609416_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6609416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:133519935(-)-10:133522773(+)__10_133500501_133525501D;SPAN=2838;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:222 GQ:33.4 PL:[0.0, 33.4, 604.0] SR:0 DR:8 LR:33.74 LO:11.86);ALT=]chr10:133522773]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134367081	+	chr10	134366070	+	.	19	0	6612760_1	19.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6612760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134366070(-)-10:134367081(+)__10_134358001_134383001D;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:160 GQ:19.3 PL:[19.3, 0.0, 369.2] SR:0 DR:19 LR:-19.37 LO:38.35);ALT=]chr10:134367081]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134387874	+	chr10	134386371	+	.	45	0	6612948_1	98.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6612948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134386371(-)-10:134387874(+)__10_134382501_134407501D;SPAN=1503;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:184 GQ:98.9 PL:[98.9, 0.0, 346.4] SR:0 DR:45 LR:-98.7 LO:106.5);ALT=]chr10:134387874]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134534060	+	chr10	134532009	+	.	11	0	6613319_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6613319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134532009(-)-10:134534060(+)__10_134529501_134554501D;SPAN=2051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:161 GQ:7 PL:[0.0, 7.0, 402.6] SR:0 DR:11 LR:7.308 LO:19.43);ALT=]chr10:134534060]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134745437	+	chr10	134743975	+	.	10	0	6614103_1	0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6614103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134743975(-)-10:134745437(+)__10_134725501_134750501D;SPAN=1462;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:163 GQ:10.9 PL:[0.0, 10.9, 415.9] SR:0 DR:10 LR:11.15 LO:17.18);ALT=]chr10:134745437]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134793926	+	chr10	134795018	-	.	4	2	6614196_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAGGC;MAPQ=60;MATEID=6614196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_134774501_134799501_155C;SPAN=1092;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:158 GQ:29.5 PL:[0.0, 29.5, 442.3] SR:2 DR:4 LR:29.6 LO:5.317);ALT=G]chr10:134795018];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	135104816	+	chr10	135105935	+	.	145	6	6615510_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTCCGTGTCCCCCATGTCCCTCCGTGTCCCCCATGTCCCTCCGTGTCCCTGTGTCCCGGGGAGCCCTACCTGTA;MAPQ=60;MATEID=6615510_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_10_135093001_135118001_196C;SPAN=1119;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:150 DP:8 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:6 DR:145 LR:-445.6 LO:445.6);ALT=A[chr10:135105935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
