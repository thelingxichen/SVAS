chr4	59944565	+	chr4	59950602	+	.	27	29	1988265_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTGT;MAPQ=60;MATEID=1988265_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_4_59927001_59952001_294C;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:66 GQ:8.6 PL:[150.5, 0.0, 8.6] SR:29 DR:27 LR:-157.8 LO:157.8);ALT=T[chr4:59950602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
