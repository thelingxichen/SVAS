chr9	66276429	+	chr14	28269626	+	.	0	21	8405829_1	47.0	.	EVDNC=ASSMB;HOMSEQ=GCAAAATA;MAPQ=53;MATEID=8405829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_28248501_28273501_448C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:80 GQ:47.6 PL:[47.6, 0.0, 146.6] SR:21 DR:0 LR:-47.65 LO:50.45);ALT=A[chr14:28269626[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	66844464	+	chr9	66842853	+	.	8	0	5867267_1	0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=5867267_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:66842853(-)-9:66844464(+)__9_66836001_66861001D;SPAN=1611;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:115 GQ:4.5 PL:[0.0, 4.5, 287.1] SR:0 DR:8 LR:4.748 LO:14.2);ALT=]chr9:66844464]A;VARTYPE=BND:DUP-th;JOINTYPE=th
