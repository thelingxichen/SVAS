chr13	113762168	+	chr13	113763575	+	.	8	0	8346188_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=8346188_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:113762168(+)-13:113763575(-)__13_113753501_113778501D;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:179 GQ:22 PL:[0.0, 22.0, 478.6] SR:0 DR:8 LR:22.09 LO:12.62);ALT=C[chr13:113763575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113796771	-	chr13	113799300	+	.	8	0	8346085_1	0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=8346085_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:113796771(-)-13:113799300(-)__13_113778001_113803001D;SPAN=2529;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:192 GQ:25.3 PL:[0.0, 25.3, 514.9] SR:0 DR:8 LR:25.61 LO:12.37);ALT=[chr13:113799300[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	114000379	+	chr13	114001595	+	.	29	0	8347761_1	74.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=8347761_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:114000379(+)-13:114001595(-)__13_113998501_114023501D;SPAN=1216;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:78 GQ:74.6 PL:[74.6, 0.0, 114.2] SR:0 DR:29 LR:-74.6 LO:75.06);ALT=A[chr13:114001595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114000542	+	chr13	114001993	+	.	17	0	8347774_1	29.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=8347774_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:114000542(+)-13:114001993(-)__13_113998501_114023501D;SPAN=1451;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:100 GQ:29 PL:[29.0, 0.0, 213.8] SR:0 DR:17 LR:-29.02 LO:37.19);ALT=A[chr13:114001993[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114771156	+	chr13	114772822	+	.	8	0	8351671_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=8351671_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:114771156(+)-13:114772822(-)__13_114758001_114783001D;SPAN=1666;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:152 GQ:14.5 PL:[0.0, 14.5, 396.0] SR:0 DR:8 LR:14.77 LO:13.2);ALT=A[chr13:114772822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
