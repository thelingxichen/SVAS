chr1	114402132	+	chr1	114414269	+	.	8	0	270697_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=270697_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:114402132(+)-1:114414269(-)__1_114390501_114415501D;SPAN=12137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=G[chr1:114414269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	114645955	-	chr1	114654368	+	.	0	45	271121_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GTGC;MAPQ=60;MATEID=271121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_114635501_114660501_81C;SPAN=8413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:45 DR:0 LR:-141.9 LO:141.9);ALT=[chr1:114654368[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	115256601	+	chr1	115258670	+	.	0	9	271987_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=271987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115248001_115273001_220C;SPAN=2069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:9 DR:0 LR:-15.08 LO:19.6);ALT=T[chr1:115258670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115263339	+	chr1	115266503	+	.	3	26	272005_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=272005_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115248001_115273001_80C;SPAN=3164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:72 GQ:69.8 PL:[69.8, 0.0, 102.8] SR:26 DR:3 LR:-69.62 LO:70.02);ALT=C[chr1:115266503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115263375	+	chr1	115267841	+	.	18	0	272006_1	43.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=272006_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:115263375(+)-1:115267841(-)__1_115248001_115273001D;SPAN=4466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:0 DR:18 LR:-43.7 LO:44.82);ALT=C[chr1:115267841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115266625	+	chr1	115267842	+	.	4	15	272014_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=272014_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_115248001_115273001_119C;SPAN=1217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:61 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:15 DR:4 LR:-36.29 LO:38.43);ALT=T[chr1:115267842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115266625	+	chr1	115268832	+	GAGTGTGTTTTGTTCACTTTTTCTGCACTGACTTTGTTGCCTTTGCCTTTGGACAAGCTATACTCGACCATGTCCCCCAGTTCCAGGCTATCAACATCACCAGAGAACTCA	6	28	272015_1	92.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GAGTGTGTTTTGTTCACTTTTTCTGCACTGACTTTGTTGCCTTTGCCTTTGGACAAGCTATACTCGACCATGTCCCCCAGTTCCAGGCTATCAACATCACCAGAGAACTCA;MAPQ=60;MATEID=272015_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_115248001_115273001_119C;SPAN=2207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:51 GQ:29.3 PL:[92.0, 0.0, 29.3] SR:28 DR:6 LR:-93.4 LO:93.4);ALT=T[chr1:115268832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115269713	+	chr1	115272878	+	.	7	9	272060_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=272060_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115272501_115297501_159C;SPAN=3165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:35 GQ:30.2 PL:[30.2, 0.0, 53.3] SR:9 DR:7 LR:-30.13 LO:30.52);ALT=T[chr1:115272878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115273270	+	chr1	115275224	+	.	12	6	272063_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=272063_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115272501_115297501_242C;SPAN=1954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:54 GQ:41.6 PL:[41.6, 0.0, 87.8] SR:6 DR:12 LR:-41.49 LO:42.46);ALT=C[chr1:115275224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115279476	+	chr1	115280583	+	.	2	3	272077_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=272077_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_115272501_115297501_161C;SPAN=1107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:55 GQ:1.5 PL:[0.0, 1.5, 135.3] SR:3 DR:2 LR:1.697 LO:7.178);ALT=C[chr1:115280583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115280695	+	chr1	115282313	+	.	0	9	272081_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=272081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115272501_115297501_229C;SPAN=1618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:55 GQ:14.9 PL:[14.9, 0.0, 117.2] SR:9 DR:0 LR:-14.81 LO:19.52);ALT=T[chr1:115282313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115292831	+	chr1	115300544	+	.	137	0	272140_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=272140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:115292831(+)-1:115300544(-)__1_115297001_115322001D;SPAN=7713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:61 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:0 DR:137 LR:-406.0 LO:406.0);ALT=A[chr1:115300544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115604854	+	chr1	115615525	+	.	0	11	272597_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=272597_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115615501_115640501_178C;SPAN=10671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:35 GQ:26.9 PL:[26.9, 0.0, 56.6] SR:11 DR:0 LR:-26.83 LO:27.46);ALT=C[chr1:115615525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115604901	+	chr1	115632022	+	.	8	0	272598_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=272598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:115604901(+)-1:115632022(-)__1_115615501_115640501D;SPAN=27121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:0 DR:8 LR:-19.91 LO:20.23);ALT=T[chr1:115632022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	115615629	+	chr1	115631985	+	.	9	5	272600_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=272600_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_115615501_115640501_135C;SPAN=16356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:5 DR:9 LR:-20.55 LO:23.07);ALT=C[chr1:115631985[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	116184707	+	chr1	116193896	+	.	9	3	273293_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=273293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_116179001_116204001_190C;SPAN=9189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:3 DR:9 LR:-16.75 LO:21.78);ALT=G[chr1:116193896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	116916087	+	chr1	116926634	+	.	8	0	274417_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=274417_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:116916087(+)-1:116926634(-)__1_116914001_116939001D;SPAN=10547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=G[chr1:116926634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	116916147	+	chr1	116927404	+	TGGACGTGATAAGTATGAGCCTGCAGCTGTTTCAGAACAAGGTGATAAAAAGGGCAAAAAGGGCAAAAAAGACAGGGACATGGATGAACTGAAGAAAGAAGTTTCTAT	0	11	274419_1	23.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=TGGACGTGATAAGTATGAGCCTGCAGCTGTTTCAGAACAAGGTGATAAAAAGGGCAAAAAGGGCAAAAAAGACAGGGACATGGATGAACTGAAGAAAGAAGTTTCTAT;MAPQ=60;MATEID=274419_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_116914001_116939001_251C;SPAN=11257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:47 GQ:23.6 PL:[23.6, 0.0, 89.6] SR:11 DR:0 LR:-23.58 LO:25.79);ALT=T[chr1:116927404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	117076733	+	chr11	3013483	+	.	6	2	274629_1	18.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=12;MATEID=274629_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_1_117061001_117086001_213C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:2 DR:6 LR:-18.55 LO:19.42);ALT=T[chr11:3013483[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	117087220	+	chr1	117113552	+	.	12	0	274686_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=274686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:117087220(+)-1:117113552(-)__1_117110001_117135001D;SPAN=26332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:27 GQ:32.3 PL:[32.3, 0.0, 32.3] SR:0 DR:12 LR:-32.3 LO:32.3);ALT=A[chr1:117113552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	117603037	+	chr1	117605008	+	.	10	0	275537_1	19.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=275537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:117603037(+)-1:117605008(-)__1_117600001_117625001D;SPAN=1971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:52 GQ:19.1 PL:[19.1, 0.0, 104.9] SR:0 DR:10 LR:-18.92 LO:22.47);ALT=T[chr1:117605008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	117945063	+	chr1	117948169	+	.	4	2	276025_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=276025_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_117943001_117968001_58C;SPAN=3106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:49 GQ:0 PL:[0.0, 0.0, 118.8] SR:2 DR:4 LR:0.0713 LO:7.387);ALT=G[chr1:117948169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	117948268	+	chr1	117957334	+	.	3	7	276029_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=276029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_117943001_117968001_263C;SPAN=9066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:54 GQ:18.5 PL:[18.5, 0.0, 110.9] SR:7 DR:3 LR:-18.38 LO:22.29);ALT=G[chr1:117957334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	117957453	+	chr1	117963190	+	.	2	7	276040_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=276040_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_117943001_117968001_124C;SPAN=5737;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:53 GQ:8.9 PL:[8.9, 0.0, 117.8] SR:7 DR:2 LR:-8.748 LO:14.48);ALT=G[chr1:117963190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	118148775	+	chr1	118165461	+	.	22	3	276395_1	65.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=276395_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_118163501_118188501_148C;SPAN=16686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:28 GQ:2.3 PL:[65.0, 0.0, 2.3] SR:3 DR:22 LR:-68.45 LO:68.45);ALT=G[chr1:118165461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	205709	+	chr11	207335	+	.	10	0	4727268_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4727268_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:205709(+)-11:207335(-)__11_196001_221001D;SPAN=1626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:0 DR:10 LR:-12.96 LO:20.79);ALT=C[chr11:207335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	237093	+	chr11	244038	+	.	12	0	4727380_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4727380_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:237093(+)-11:244038(-)__11_220501_245501D;SPAN=6945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:83 GQ:17.3 PL:[17.3, 0.0, 182.3] SR:0 DR:12 LR:-17.13 LO:25.33);ALT=G[chr11:244038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	237146	+	chr11	238998	+	.	34	24	4727382_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=4727382_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_220501_245501_322C;SPAN=1852;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:86 GQ:89 PL:[118.7, 0.0, 89.0] SR:24 DR:34 LR:-118.9 LO:118.9);ALT=T[chr11:238998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	410030	+	chr11	414823	+	.	0	16	4728674_1	31.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4728674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_392001_417001_297C;SPAN=4793;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:79 GQ:31.4 PL:[31.4, 0.0, 160.1] SR:16 DR:0 LR:-31.41 LO:36.36);ALT=G[chr11:414823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	500657	+	chr11	502061	+	.	22	48	4728767_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4728767_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_490001_515001_239C;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:102 GQ:55.1 PL:[190.4, 0.0, 55.1] SR:48 DR:22 LR:-194.2 LO:194.2);ALT=G[chr11:502061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	500693	+	chr11	507133	+	.	19	0	4728768_1	41.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4728768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:500693(+)-11:507133(-)__11_490001_515001D;SPAN=6440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:79 GQ:41.3 PL:[41.3, 0.0, 150.2] SR:0 DR:19 LR:-41.32 LO:44.8);ALT=A[chr11:507133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	500695	+	chr11	504425	+	.	9	0	4728769_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4728769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:500695(+)-11:504425(-)__11_490001_515001D;SPAN=3730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:100 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.617 LO:17.02);ALT=C[chr11:504425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	502218	+	chr11	504426	+	.	14	0	4728777_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4728777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:502218(+)-11:504426(-)__11_490001_515001D;SPAN=2208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:114 GQ:15.5 PL:[15.5, 0.0, 259.7] SR:0 DR:14 LR:-15.33 LO:28.48);ALT=G[chr11:504426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	502251	+	chr11	507113	+	.	42	6	4728778_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4728778_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_490001_515001_217C;SPAN=4862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:72 GQ:50 PL:[122.6, 0.0, 50.0] SR:6 DR:42 LR:-124.0 LO:124.0);ALT=T[chr11:507113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	502289	+	chr11	504838	+	.	11	0	4728780_1	19.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4728780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:502289(+)-11:504838(-)__11_490001_515001D;SPAN=2549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:0 DR:11 LR:-19.51 LO:24.29);ALT=C[chr11:504838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	736900	+	chr11	3917255	+	.	18	0	4729955_1	48.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4729955_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:736900(+)-11:3917255(-)__11_735001_760001D;SPAN=3180355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:39 GQ:45.5 PL:[48.8, 0.0, 45.5] SR:0 DR:18 LR:-48.86 LO:48.86);ALT=G[chr11:3917255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3917414	+	chr11	737067	+	.	37	25	4729956_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCAAAGTGCTGGGATTACAGGCG;MAPQ=60;MATEID=4729956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_735001_760001_113C;SPAN=3180347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:29 GQ:15 PL:[165.0, 15.0, 0.0] SR:25 DR:37 LR:-165.0 LO:165.0);ALT=]chr11:3917414]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	747578	+	chr11	755878	+	.	0	64	4730001_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4730001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_735001_760001_243C;SPAN=8300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:181 GQ:99 PL:[162.5, 0.0, 274.7] SR:64 DR:0 LR:-162.2 LO:163.9);ALT=G[chr11:755878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	747591	+	chr11	758948	+	.	19	0	4730002_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4730002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:747591(+)-11:758948(-)__11_735001_760001D;SPAN=11357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:126 GQ:28.7 PL:[28.7, 0.0, 276.2] SR:0 DR:19 LR:-28.58 LO:40.48);ALT=C[chr11:758948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	756004	+	chr11	760120	+	CACAAGAGGACCAGATTAAAAATGCTATTGATAAACTTTTTGTGTTGTTTGGAGCAGAAATACTAAAGAAGATTCCGGGCCGAGTATCCACAGAAGTAGACGCA	5	140	4730030_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CACAAGAGGACCAGATTAAAAATGCTATTGATAAACTTTTTGTGTTGTTTGGAGCAGAAATACTAAAGAAGATTCCGGGCCGAGTATCCACAGAAGTAGACGCA;MAPQ=60;MATEID=4730030_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_735001_760001_403C;SPAN=4116;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:128 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:140 DR:5 LR:-425.8 LO:425.8);ALT=T[chr11:760120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	759058	+	chr11	760120	+	.	8	47	4730044_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=4730044_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCTC;SCTG=c_11_735001_760001_403C;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:61 GQ:12.9 PL:[171.6, 12.9, 0.0] SR:47 DR:8 LR:-171.4 LO:171.4);ALT=G[chr11:760120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	760254	+	chr11	763344	+	.	14	23	4729626_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4729626_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_759501_784501_175C;SPAN=3090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:86 GQ:82.4 PL:[82.4, 0.0, 125.3] SR:23 DR:14 LR:-82.33 LO:82.84);ALT=G[chr11:763344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	763520	+	chr11	764813	+	GGTAAAGAGTGTCACTAAAATCTACAACTACTACAAGAAGTTTAGCTACAAAACCATTGTCATGGGCGCCTCCTTCCGCAACACGGGCGAGATCAAAGCACTGGCCGGCTGTGACTTCCTCACCATCTCACCCAAGCTCCTGGGAGAGCTGCTGCAGGACAACGCCAAGCTGGTGCCTGTGCTCTCAGCCAAGGCGGCCCAAGCCAGTGACCTGGAAAAAATCCACCTGGATGAGAAGTCTTTCCGTTGGTTGCACAACGAGGACCAGATGGCTGTGGAGAAGCTCTCTGACGGGATCCGCAAGTTTGCCGCTGATGCAGTGAAGCTGGAGCGGATGCTGACA	0	286	4729640_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GGTAAAGAGTGTCACTAAAATCTACAACTACTACAAGAAGTTTAGCTACAAAACCATTGTCATGGGCGCCTCCTTCCGCAACACGGGCGAGATCAAAGCACTGGCCGGCTGTGACTTCCTCACCATCTCACCCAAGCTCCTGGGAGAGCTGCTGCAGGACAACGCCAAGCTGGTGCCTGTGCTCTCAGCCAAGGCGGCCCAAGCCAGTGACCTGGAAAAAATCCACCTGGATGAGAAGTCTTTCCGTTGGTTGCACAACGAGGACCAGATGGCTGTGGAGAAGCTCTCTGACGGGATCCGCAAGTTTGCCGCTGATGCAGTGAAGCTGGAGCGGATGCTGACA;MAPQ=60;MATEID=4729640_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_759501_784501_97C;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:286 DP:140 GQ:77.3 PL:[848.3, 77.3, 0.0] SR:286 DR:0 LR:-848.3 LO:848.3);ALT=G[chr11:764813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	810084	+	chr11	812532	+	.	41	0	4729798_1	16.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4729798_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:810084(+)-11:812532(-)__11_808501_833501D;SPAN=2448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:440 GQ:16.2 PL:[16.2, 0.0, 1053.0] SR:0 DR:41 LR:-16.13 LO:78.18);ALT=G[chr11:812532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	819910	+	chr11	821627	+	.	7	11	4729840_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGAG;MAPQ=60;MATEID=4729840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_808501_833501_24C;SPAN=1717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:11 DR:7 LR:-20.92 LO:26.38);ALT=G[chr11:821627[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	833079	+	chr11	836060	+	.	72	0	4729721_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4729721_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:833079(+)-11:836060(-)__11_833001_858001D;SPAN=2981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:56 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:0 DR:72 LR:-211.3 LO:211.3);ALT=G[chr11:836060[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	840481	+	chr11	842413	+	.	98	32	4729746_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4729746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_833001_858001_71C;SPAN=1932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:117 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:32 DR:98 LR:-346.6 LO:346.6);ALT=C[chr11:842413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	903113	+	chr11	904706	+	.	0	32	4729929_1	74.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4729929_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_882001_907001_155C;SPAN=1593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:115 GQ:74.6 PL:[74.6, 0.0, 203.3] SR:32 DR:0 LR:-74.48 LO:77.84);ALT=T[chr11:904706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	903159	+	chr11	910773	+	.	23	0	4730263_1	65.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4730263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:903159(+)-11:910773(-)__11_906501_931501D;SPAN=7614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:37 GQ:23 PL:[65.9, 0.0, 23.0] SR:0 DR:23 LR:-66.98 LO:66.98);ALT=G[chr11:910773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	904883	+	chr11	910774	+	.	29	0	4730265_1	85.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4730265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:904883(+)-11:910774(-)__11_906501_931501D;SPAN=5891;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:39 GQ:9.2 PL:[85.1, 0.0, 9.2] SR:0 DR:29 LR:-88.68 LO:88.68);ALT=C[chr11:910774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1119598	+	chr11	1118254	+	.	27	1	4730830_1	64.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AGTG;MAPQ=60;MATEID=4730830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1102501_1127501_61C;SECONDARY;SPAN=1344;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:103 GQ:64.7 PL:[64.7, 0.0, 183.5] SR:1 DR:27 LR:-64.52 LO:67.77);ALT=]chr11:1119598]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	1290025	-	chr12	108935074	+	.	3	3	4731218_1	2.0	.	DISC_MAPQ=8;EVDNC=ASDIS;HOMSEQ=TTGGGAGGCTGAGGCAGGAGAATCGCTTGAA;MAPQ=42;MATEID=4731218_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_1274001_1299001_1C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:51 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:3 DR:3 LR:-2.688 LO:9.65);ALT=[chr12:108935074[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	1317025	+	chr11	1330693	+	.	0	11	4731318_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=4731318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1323001_1348001_47C;SPAN=13668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:34 GQ:27.2 PL:[27.2, 0.0, 53.6] SR:11 DR:0 LR:-27.1 LO:27.63);ALT=C[chr11:1330693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1643100	-	chr11	71249252	+	.	8	0	4732324_1	16.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4732324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:1643100(-)-11:71249252(-)__11_1641501_1666501D;SPAN=69606152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=[chr11:71249252[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	1776260	+	chr11	1778553	+	.	2	5	4732759_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4732759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1764001_1789001_280C;SPAN=2293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:5 DR:2 LR:-2.788 LO:13.35);ALT=T[chr11:1778553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1778787	+	chr11	1780196	+	.	0	7	4732764_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=4732764_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1764001_1789001_302C;SPAN=1409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:70 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:7 DR:0 LR:-4.142 LO:13.57);ALT=C[chr11:1780196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1780869	+	chr11	1782538	+	.	4	88	4732772_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4732772_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_1764001_1789001_162C;SPAN=1669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:138 GQ:74.9 PL:[259.7, 0.0, 74.9] SR:88 DR:4 LR:-265.3 LO:265.3);ALT=C[chr11:1782538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1780869	+	chr11	1785021	+	GTCCATGTAGTTCTTGAGCACCTCGGGAATGGGCCCCTCGGTCACGGCTGGCACCGCCTGGGAGTACTTTGAGACGGGGCCTTTGGCAATCAGGTCCTCCACAGAGCCCCCAACCTCCGACATGGTCCGGCGGATGGACGTGAACTTGTGCAGCGGGAT	89	122	4732773_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=GTCCATGTAGTTCTTGAGCACCTCGGGAATGGGCCCCTCGGTCACGGCTGGCACCGCCTGGGAGTACTTTGAGACGGGGCCTTTGGCAATCAGGTCCTCCACAGAGCCCCCAACCTCCGACATGGTCCGGCGGATGGACGTGAACTTGTGCAGCGGGAT;MAPQ=60;MATEID=4732773_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_1764001_1789001_162C;SPAN=4152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:93 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:122 DR:89 LR:-458.8 LO:458.8);ALT=C[chr11:1785021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1782701	+	chr11	1785021	+	.	138	28	4732777_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=4732777_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_1764001_1789001_162C;SPAN=2320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:92 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:28 DR:138 LR:-429.1 LO:429.1);ALT=G[chr11:1785021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1874428	+	chr11	1901316	+	.	102	3	4733094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4733094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1862001_1887001_344C;SPAN=26888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:61 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:3 DR:102 LR:-310.3 LO:310.3);ALT=G[chr11:1901316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1901454	+	chr11	1902662	+	.	0	118	4732977_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4732977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1886501_1911501_21C;SPAN=1208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:118 DP:223 GQ:99 PL:[329.3, 0.0, 210.5] SR:118 DR:0 LR:-330.5 LO:330.5);ALT=T[chr11:1902662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1901455	+	chr11	1904649	+	.	2	6	4732978_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4732978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1886501_1911501_252C;SPAN=3194;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:164 GQ:17.8 PL:[0.0, 17.8, 432.4] SR:6 DR:2 LR:18.02 LO:12.93);ALT=G[chr11:1904649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1902827	+	chr11	1904645	+	.	10	24	4732982_1	84.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACAGG;MAPQ=60;MATEID=4732982_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_1886501_1911501_46C;SPAN=1818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:92 GQ:84.2 PL:[84.2, 0.0, 137.0] SR:24 DR:10 LR:-84.01 LO:84.76);ALT=G[chr11:1904645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1905811	+	chr11	1907960	+	.	9	43	4733001_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4733001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1886501_1911501_317C;SPAN=2149;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:126 GQ:99 PL:[131.0, 0.0, 173.9] SR:43 DR:9 LR:-130.9 LO:131.3);ALT=G[chr11:1907960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1908806	+	chr11	1913002	+	.	28	12	4733284_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4733284_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1911001_1936001_14C;SPAN=4196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:57 GQ:24.2 PL:[113.3, 0.0, 24.2] SR:12 DR:28 LR:-116.5 LO:116.5);ALT=G[chr11:1913002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1910839	+	chr11	1913002	+	.	54	6	4733285_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4733285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1911001_1936001_90C;SPAN=2163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:57 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:6 DR:54 LR:-168.3 LO:168.3);ALT=G[chr11:1913002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1915274	+	chr11	1936956	+	ATG	96	13	4733453_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=ATG;MAPQ=60;MATEID=4733453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1935501_1960501_133C;SPAN=21682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:85 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:13 DR:96 LR:-307.0 LO:307.0);ALT=G[chr11:1936956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1918400	+	chr11	1923818	+	.	10	0	4733326_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:1918400(+)-11:1923818(-)__11_1911001_1936001D;SPAN=5418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=A[chr11:1923818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1918402	+	chr11	1924332	+	.	12	0	4733327_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4733327_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:1918402(+)-11:1924332(-)__11_1911001_1936001D;SPAN=5930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:92 GQ:14.9 PL:[14.9, 0.0, 206.3] SR:0 DR:12 LR:-14.69 LO:24.74);ALT=T[chr11:1924332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1968611	+	chr11	1972129	+	.	33	8	4733595_1	87.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=4733595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1960001_1985001_110C;SPAN=3518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:128 GQ:87.5 PL:[87.5, 0.0, 222.8] SR:8 DR:33 LR:-87.46 LO:90.74);ALT=T[chr11:1972129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1968660	+	chr11	1977484	+	.	10	0	4733597_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733597_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:1968660(+)-11:1977484(-)__11_1960001_1985001D;SPAN=8824;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:0 DR:10 LR:-10.79 LO:20.31);ALT=A[chr11:1977484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1968663	+	chr11	1973389	+	.	34	0	4733599_1	74.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733599_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:1968663(+)-11:1973389(-)__11_1960001_1985001D;SPAN=4726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:139 GQ:74.6 PL:[74.6, 0.0, 262.7] SR:0 DR:34 LR:-74.58 LO:80.46);ALT=A[chr11:1973389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1972251	+	chr11	1973357	+	.	7	81	4733608_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4733608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1960001_1985001_176C;SPAN=1106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:84 DP:112 GQ:22.7 PL:[247.1, 0.0, 22.7] SR:81 DR:7 LR:-257.5 LO:257.5);ALT=A[chr11:1973357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	1974086	+	chr11	1977485	+	.	4	53	4733614_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4733614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1960001_1985001_160C;SPAN=3399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:112 GQ:99 PL:[158.0, 0.0, 111.8] SR:53 DR:4 LR:-158.2 LO:158.2);ALT=G[chr11:1977485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2079880	+	chr11	2076953	+	.	8	0	4733899_1	2.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4733899_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2076953(-)-11:2079880(+)__11_2058001_2083001D;SPAN=2927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=]chr11:2079880]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	2083082	+	chr11	2079023	+	.	17	0	4733904_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733904_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2079023(-)-11:2083082(+)__11_2058001_2083001D;SPAN=4059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:52 GQ:42.2 PL:[42.2, 0.0, 81.8] SR:0 DR:17 LR:-42.03 LO:42.8);ALT=]chr11:2083082]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	2083093	+	chr11	2081944	+	.	26	0	4733917_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2081944(-)-11:2083093(+)__11_2058001_2083001D;SPAN=1149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:45 GQ:34.1 PL:[73.7, 0.0, 34.1] SR:0 DR:26 LR:-74.35 LO:74.35);ALT=]chr11:2083093]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	2084549	+	chr11	2082478	+	.	43	0	4733702_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4733702_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2082478(-)-11:2084549(+)__11_2082501_2107501D;SPAN=2071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:77 GQ:65 PL:[121.1, 0.0, 65.0] SR:0 DR:43 LR:-122.0 LO:122.0);ALT=]chr11:2084549]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	2319153	+	chr11	2320657	+	.	0	17	4734533_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4734533_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_2303001_2328001_246C;SPAN=1504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:71 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:17 DR:0 LR:-36.88 LO:40.05);ALT=T[chr11:2320657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2320974	+	chr11	2323039	+	.	10	0	4734539_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4734539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2320974(+)-11:2323039(-)__11_2303001_2328001D;SPAN=2065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:0 DR:10 LR:-13.5 LO:20.92);ALT=C[chr11:2323039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2323500	+	chr11	2325335	+	.	17	0	4734545_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4734545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2323500(+)-11:2325335(-)__11_2303001_2328001D;SPAN=1835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:76 GQ:35.6 PL:[35.6, 0.0, 147.8] SR:0 DR:17 LR:-35.53 LO:39.47);ALT=G[chr11:2325335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2324188	+	chr11	2325336	+	.	0	24	4734548_1	56.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4734548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_2303001_2328001_164C;SPAN=1148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:85 GQ:56.3 PL:[56.3, 0.0, 148.7] SR:24 DR:0 LR:-56.2 LO:58.56);ALT=G[chr11:2325336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2422079	+	chr11	2423522	+	.	16	0	4734615_1	32.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4734615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2422079(+)-11:2423522(-)__11_2401001_2426001D;SPAN=1443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:76 GQ:32.3 PL:[32.3, 0.0, 151.1] SR:0 DR:16 LR:-32.23 LO:36.67);ALT=G[chr11:2423522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2997380	+	chr11	3013482	+	.	8	0	4736269_1	21.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=4736269_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2997380(+)-11:3013482(-)__11_3013501_3038501D;SPAN=16102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:21.5 PL:[21.5, 0.0, 21.5] SR:0 DR:8 LR:-21.53 LO:21.53);ALT=T[chr11:3013482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3147788	+	chr11	3150242	+	.	6	16	4736770_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4736770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_3136001_3161001_251C;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:16 DR:6 LR:-42.57 LO:43.16);ALT=G[chr11:3150242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3147840	+	chr11	3186445	+	.	8	0	4736919_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4736919_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:3147840(+)-11:3186445(-)__11_3185001_3210001D;SPAN=38605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:21.5 PL:[21.5, 0.0, 21.5] SR:0 DR:8 LR:-21.53 LO:21.53);ALT=T[chr11:3186445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3150405	+	chr11	3186445	+	.	11	0	4736920_1	31.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4736920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:3150405(+)-11:3186445(-)__11_3185001_3210001D;SPAN=36040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:18 GQ:11.6 PL:[31.4, 0.0, 11.6] SR:0 DR:11 LR:-31.89 LO:31.89);ALT=A[chr11:3186445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3416445	+	chr11	3615515	+	.	12	0	4737877_1	36.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=4737877_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:3416445(+)-11:3615515(-)__11_3601501_3626501D;SPAN=199070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:13 GQ:3.3 PL:[36.3, 3.3, 0.0] SR:0 DR:12 LR:-36.31 LO:36.31);ALT=A[chr11:3615515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3800487	+	chr11	3803272	+	.	0	13	4739079_1	19.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4739079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_3797501_3822501_390C;SPAN=2785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:88 GQ:19.1 PL:[19.1, 0.0, 194.0] SR:13 DR:0 LR:-19.07 LO:27.57);ALT=T[chr11:3803272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3803376	+	chr11	3818630	+	.	0	8	4739094_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4739094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_3797501_3822501_266C;SPAN=15254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:77 GQ:5.6 PL:[5.6, 0.0, 180.5] SR:8 DR:0 LR:-5.547 LO:15.65);ALT=C[chr11:3818630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3849439	+	chr11	3862122	+	.	164	4	4739006_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=4739006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_3846501_3871501_359C;SPAN=12683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:165 DP:145 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:4 DR:164 LR:-488.5 LO:488.5);ALT=G[chr11:3862122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3908980	+	chr11	3909989	-	.	8	0	4739288_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4739288_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:3908980(+)-11:3909989(+)__11_3895501_3920501D;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:80 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:0 DR:8 LR:-4.734 LO:15.51);ALT=C]chr11:3909989];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	4116261	+	chr11	4123221	+	.	0	9	4740028_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4740028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_4091501_4116501_236C;SPAN=6960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:9 DR:0 LR:-20.5 LO:21.66);ALT=G[chr11:4123221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	4779578	+	chr11	4778427	+	.	4	2	4741798_1	0	.	DISC_MAPQ=51;EVDNC=ASDIS;MAPQ=60;MATEID=4741798_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_4777501_4802501_230C;SPAN=1151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:86 GQ:6.6 PL:[0.0, 6.6, 221.1] SR:2 DR:4 LR:6.795 LO:8.471);ALT=]chr11:4779578]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	5711129	+	chr11	5717395	+	.	21	5	4744175_1	54.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4744175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_5708501_5733501_243C;SPAN=6266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:92 GQ:54.5 PL:[54.5, 0.0, 166.7] SR:5 DR:21 LR:-54.3 LO:57.58);ALT=G[chr11:5717395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	6623447	+	chr11	6624633	+	.	0	6	4746530_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4746530_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_6615001_6640001_77C;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:6 DR:0 LR:3.764 LO:10.62);ALT=T[chr11:6624633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	6625108	+	chr11	6629274	+	.	13	0	4746537_1	18.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4746537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:6625108(+)-11:6629274(-)__11_6615001_6640001D;SPAN=4166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:91 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.26 LO:27.36);ALT=G[chr11:6629274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	6625591	+	chr11	6629275	+	.	9	18	4746538_1	61.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4746538_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGGG;SCTG=c_11_6615001_6640001_335C;SPAN=3684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:92 GQ:61.1 PL:[61.1, 0.0, 160.1] SR:18 DR:9 LR:-60.9 LO:63.46);ALT=G[chr11:6629275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	6639007	+	chr11	6640426	+	.	18	2	4746583_1	54.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4746583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_6615001_6640001_1C;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:42 GQ:44.9 PL:[54.8, 0.0, 44.9] SR:2 DR:18 LR:-54.67 LO:54.67);ALT=C[chr11:6640426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	16960731	-	chr11	16961895	+	.	8	0	4774335_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4774335_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:16960731(-)-11:16961895(-)__11_16954001_16979001D;SPAN=1164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=[chr11:16961895[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	17097178	+	chr11	17099164	+	.	53	0	4774938_1	90.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=4774938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:17097178(+)-11:17099164(-)__11_17076501_17101501D;SPAN=1986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:314 GQ:90.1 PL:[90.1, 0.0, 671.0] SR:0 DR:53 LR:-89.88 LO:115.8);ALT=G[chr11:17099164[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17298688	+	chr11	17316870	+	.	46	0	4775825_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4775825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:17298688(+)-11:17316870(-)__11_17297001_17322001D;SPAN=18182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:93 GQ:97.1 PL:[126.8, 0.0, 97.1] SR:0 DR:46 LR:-126.8 LO:126.8);ALT=C[chr11:17316870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17298718	+	chr11	17304332	+	.	88	0	4775826_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4775826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:17298718(+)-11:17304332(-)__11_17297001_17322001D;SPAN=5614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:94 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:0 DR:88 LR:-277.3 LO:277.3);ALT=T[chr11:17304332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17304490	+	chr11	17316871	+	.	9	66	4775851_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4775851_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_17297001_17322001_67C;SPAN=12381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:74 DP:104 GQ:34.7 PL:[216.2, 0.0, 34.7] SR:66 DR:9 LR:-223.4 LO:223.4);ALT=C[chr11:17316871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17317758	+	chr11	17323289	+	.	0	17	4775896_1	45.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4775896_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_17297001_17322001_347C;SPAN=5531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:39 GQ:45.5 PL:[45.5, 0.0, 48.8] SR:17 DR:0 LR:-45.55 LO:45.56);ALT=G[chr11:17323289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17323417	+	chr11	17331117	+	.	0	81	4775978_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4775978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_17321501_17346501_135C;SPAN=7700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:104 GQ:11.6 PL:[239.3, 0.0, 11.6] SR:81 DR:0 LR:-251.3 LO:251.3);ALT=G[chr11:17331117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	17331223	+	chr11	17332371	+	.	0	34	4775999_1	90.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4775999_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_17321501_17346501_166C;SPAN=1148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:82 GQ:90.2 PL:[90.2, 0.0, 106.7] SR:34 DR:0 LR:-90.02 LO:90.12);ALT=G[chr11:17332371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	18124895	+	chr11	18127454	+	.	0	8	4777917_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4777917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_18105501_18130501_32C;SPAN=2559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:111 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:8 DR:0 LR:3.665 LO:14.32);ALT=T[chr11:18127454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	18210596	-	chr12	110318131	+	.	15	0	5334339_1	42.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=5334339_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:18210596(-)-12:110318131(-)__12_110299001_110324001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:26 GQ:19.4 PL:[42.5, 0.0, 19.4] SR:0 DR:15 LR:-42.88 LO:42.88);ALT=[chr12:110318131[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	18416183	+	chr11	18418365	+	.	68	9	4779172_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4779172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_18399501_18424501_377C;SPAN=2182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:92 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:9 DR:68 LR:-346.6 LO:346.6);ALT=G[chr11:18418365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	18427155	+	chr11	18428669	+	.	14	0	4779225_1	22.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=4779225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:18427155(+)-11:18428669(-)__11_18424001_18449001D;SPAN=1514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:88 GQ:22.4 PL:[22.4, 0.0, 190.7] SR:0 DR:14 LR:-22.37 LO:30.18);ALT=T[chr11:18428669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	18541152	+	chr11	18548322	+	.	4	3	4779314_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4779314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_18546501_18571501_284C;SPAN=7170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:50 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:3 DR:4 LR:-2.959 LO:9.695);ALT=T[chr11:18548322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71159931	+	chr11	71162733	+	.	6	5	4909566_1	3.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4909566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_71148001_71173001_216C;SPAN=2802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:73 GQ:3.5 PL:[3.5, 0.0, 171.8] SR:5 DR:6 LR:-3.33 LO:13.44);ALT=G[chr11:71162733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71164370	+	chr11	71169472	+	.	16	0	4909571_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4909571_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:71164370(+)-11:71169472(-)__11_71148001_71173001D;SPAN=5102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:88 GQ:29 PL:[29.0, 0.0, 184.1] SR:0 DR:16 LR:-28.97 LO:35.52);ALT=T[chr11:71169472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71164429	+	chr11	71166156	+	.	16	18	4909572_1	59.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=4909572_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_11_71148001_71173001_6C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:87 GQ:59 PL:[59.0, 0.0, 151.4] SR:18 DR:16 LR:-58.96 LO:61.23);ALT=T[chr11:71166156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71169591	+	chr11	71174478	+	.	0	9	4909584_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4909584_2;MATENM=1;NM=1;NUMPARTS=4;SCTG=c_11_71148001_71173001_6C;SPAN=4887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:9 DR:0 LR:-17.52 LO:20.4);ALT=G[chr11:71174478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71209576	+	chr11	71212345	+	.	2	4	4909837_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=4909837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_71197001_71222001_248C;SPAN=2769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:68 GQ:1.4 PL:[1.4, 0.0, 163.1] SR:4 DR:2 LR:-1.383 LO:11.29);ALT=T[chr11:71212345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71809955	+	chr11	71814227	+	.	71	0	4911931_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4911931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:71809955(+)-11:71814227(-)__11_71809501_71834501D;SPAN=4272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:111 GQ:62.6 PL:[204.5, 0.0, 62.6] SR:0 DR:71 LR:-208.3 LO:208.3);ALT=A[chr11:71814227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71810304	+	chr11	71814228	+	.	118	33	4911933_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4911933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_71809501_71834501_228C;SPAN=3924;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:131 DP:137 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:33 DR:118 LR:-406.0 LO:406.0);ALT=T[chr11:71814228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	71822543	+	chr11	71823696	+	.	30	11	4911965_1	91.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4911965_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_71809501_71834501_218C;SPAN=1153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:102 GQ:91.4 PL:[91.4, 0.0, 154.1] SR:11 DR:30 LR:-91.2 LO:92.14);ALT=C[chr11:71823696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	72525560	+	chr11	72528799	+	.	16	0	4913691_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4913691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:72525560(+)-11:72528799(-)__11_72520001_72545001D;SPAN=3239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:77 GQ:32 PL:[32.0, 0.0, 154.1] SR:0 DR:16 LR:-31.96 LO:36.56);ALT=C[chr11:72528799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	72525608	+	chr11	72527773	+	.	34	20	4913692_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4913692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_72520001_72545001_287C;SPAN=2165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:81 GQ:87.2 PL:[107.0, 0.0, 87.2] SR:20 DR:34 LR:-106.9 LO:106.9);ALT=T[chr11:72527773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73087555	+	chr11	73101589	+	.	13	0	4915010_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4915010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:73087555(+)-11:73101589(-)__11_73083501_73108501D;SPAN=14034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:77 GQ:22.1 PL:[22.1, 0.0, 164.0] SR:0 DR:13 LR:-22.05 LO:28.39);ALT=C[chr11:73101589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73584440	+	chr11	73587802	+	.	99	8	4916857_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4916857_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_73573501_73598501_66C;SPAN=3362;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:87 GQ:27 PL:[297.0, 27.0, 0.0] SR:8 DR:99 LR:-297.1 LO:297.1);ALT=C[chr11:73587802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73686167	+	chr11	73687686	+	CTTTGTAGAAGGCTCGGGGCCCCTCCTTCTGGAGCATGGTAAGGGCACAGTGGCCAGCGCTACTGTACTGGCCCAGGGCAGAGTTCATGTATCTCGTCTTGACCACGTCTACAGGGGAGGCGATGACAGTGGTGCAGAAGCCTGCCCCAAAGGCAGAAGTGAAGTGGCAAGGGAGGTCAT	2	12	4917271_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTTTGTAGAAGGCTCGGGGCCCCTCCTTCTGGAGCATGGTAAGGGCACAGTGGCCAGCGCTACTGTACTGGCCCAGGGCAGAGTTCATGTATCTCGTCTTGACCACGTCTACAGGGGAGGCGATGACAGTGGTGCAGAAGCCTGCCCCAAAGGCAGAAGTGAAGTGGCAAGGGAGGTCAT;MAPQ=60;MATEID=4917271_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_73671501_73696501_278C;SPAN=1519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:12 DR:2 LR:-21.19 LO:26.47);ALT=C[chr11:73687686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73689523	+	chr11	73692521	+	.	5	52	4917281_1	99.0	.	DISC_MAPQ=48;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4917281_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_73671501_73696501_119C;SPAN=2998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:128 GQ:99 PL:[146.9, 0.0, 163.4] SR:52 DR:5 LR:-146.9 LO:146.9);ALT=C[chr11:73692521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73689523	+	chr11	73693765	+	CGGCTTTGTAAGGTCTCACGGTGAGGCCTCCAAGATCAAGCTTCTCTAAAGGTGTCCCGTTCTTCAAAGCTGCCAGTGGCTATCATGGCCCGATCCCCTTGGTTTTCCATAGAAAATGGGTGGGAGACGAAACACCTAATGGTCATACTATGTGT	46	92	4917282_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CGGCTTTGTAAGGTCTCACGGTGAGGCCTCCAAGATCAAGCTTCTCTAAAGGTGTCCCGTTCTTCAAAGCTGCCAGTGGCTATCATGGCCCGATCCCCTTGGTTTTCCATAGAAAATGGGTGGGAGACGAAACACCTAATGGTCATACTATGTGT;MAPQ=60;MATEID=4917282_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_73671501_73696501_119C;SPAN=4242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:129 GQ:24.9 PL:[363.0, 24.9, 0.0] SR:92 DR:46 LR:-366.8 LO:366.8);ALT=C[chr11:73693765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	73692678	+	chr11	73693765	+	.	118	35	4917290_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=4917290_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_11_73671501_73696501_119C;SPAN=1087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:149 GQ:13.9 PL:[389.4, 13.9, 0.0] SR:35 DR:118 LR:-402.6 LO:402.6);ALT=C[chr11:73693765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108079745	+	chr12	108082391	+	.	20	0	5327965_1	42.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5327965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:108079745(+)-12:108082391(-)__12_108069501_108094501D;SPAN=2646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:87 GQ:42.5 PL:[42.5, 0.0, 167.9] SR:0 DR:20 LR:-42.45 LO:46.71);ALT=C[chr12:108082391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108079750	+	chr12	108086588	+	AGAGCTGAGTAAAGAAGAAGTAAAACGCCTCATTGCTGAGGCAAAGGAGAAATTGCAAGAAGAAGGTGGTGGCAGTGATGAAGAGGAGACAGGCAGTCCTTCAGAAGATGGCATGCAGAGTGCACGCACCCAGGCACGCCCAAGAGAGCCCCTGGAGGATGGTGACCCAGAGGATGACAGGACGCTTGATGATGATGAGCTGGCTGAGTACGACTTAGATAAATATGATGAGGAAGGTGACC	0	19	5327967_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AGAGCTGAGTAAAGAAGAAGTAAAACGCCTCATTGCTGAGGCAAAGGAGAAATTGCAAGAAGAAGGTGGTGGCAGTGATGAAGAGGAGACAGGCAGTCCTTCAGAAGATGGCATGCAGAGTGCACGCACCCAGGCACGCCCAAGAGAGCCCCTGGAGGATGGTGACCCAGAGGATGACAGGACGCTTGATGATGATGAGCTGGCTGAGTACGACTTAGATAAATATGATGAGGAAGGTGACC;MAPQ=60;MATEID=5327967_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_108069501_108094501_14C;SPAN=6838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:72 GQ:43.4 PL:[43.4, 0.0, 129.2] SR:19 DR:0 LR:-43.21 LO:45.7);ALT=T[chr12:108086588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108086873	+	chr12	108090250	+	.	0	11	5327982_1	17.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5327982_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_108069501_108094501_159C;SPAN=3377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:11 DR:0 LR:-17.89 LO:23.8);ALT=G[chr12:108090250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108956481	+	chr12	108959094	+	.	18	0	5330345_1	37.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5330345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:108956481(+)-12:108959094(-)__12_108951501_108976501D;SPAN=2613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:80 GQ:37.7 PL:[37.7, 0.0, 156.5] SR:0 DR:18 LR:-37.74 LO:41.84);ALT=T[chr12:108959094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108956514	+	chr12	108958053	+	.	28	19	5330346_1	97.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5330346_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_108951501_108976501_342C;SPAN=1539;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:79 GQ:94.1 PL:[97.4, 0.0, 94.1] SR:19 DR:28 LR:-97.44 LO:97.44);ALT=T[chr12:108958053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	108959209	+	chr12	108960965	+	.	0	10	5330358_1	12.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=5330358_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_108951501_108976501_194C;SPAN=1756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:10 DR:0 LR:-12.69 LO:20.72);ALT=T[chr12:108960965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	109018117	+	chr12	109027513	+	.	22	0	5330423_1	61.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5330423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:109018117(+)-12:109027513(-)__12_109025001_109050001D;SPAN=9396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:42 GQ:38.3 PL:[61.4, 0.0, 38.3] SR:0 DR:22 LR:-61.46 LO:61.46);ALT=T[chr12:109027513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	109095078	+	chr12	109125233	+	.	8	0	5330684_1	16.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5330684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:109095078(+)-12:109125233(-)__12_109123001_109148001D;SPAN=30155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=C[chr12:109125233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110006714	+	chr12	110011234	+	.	12	0	5333274_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5333274_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110006714(+)-12:110011234(-)__12_110005001_110030001D;SPAN=4520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:0 DR:12 LR:-17.67 LO:25.46);ALT=C[chr12:110011234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110338231	+	chr12	110340832	+	.	12	9	5334306_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5334306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110323501_110348501_337C;SPAN=2601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:89 GQ:28.7 PL:[28.7, 0.0, 187.1] SR:9 DR:12 LR:-28.7 LO:35.43);ALT=T[chr12:110340832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110427609	+	chr12	110429432	+	.	0	12	5334708_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5334708_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110421501_110446501_73C;SPAN=1823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:12 DR:0 LR:-18.21 LO:25.61);ALT=T[chr12:110429432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110429566	+	chr12	110433978	+	.	18	8	5334715_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5334715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110421501_110446501_102C;SPAN=4412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:92 GQ:41.3 PL:[41.3, 0.0, 179.9] SR:8 DR:18 LR:-41.1 LO:46.15);ALT=C[chr12:110433978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110466395	+	chr12	110486168	+	.	12	9	5334831_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5334831_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110470501_110495501_295C;SPAN=19773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:9 DR:12 LR:-35.16 LO:36.62);ALT=C[chr12:110486168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110480456	+	chr12	110486232	+	.	11	0	5334860_1	8.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5334860_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110480456(+)-12:110486232(-)__12_110470501_110495501D;SPAN=5776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:105 GQ:8 PL:[8.0, 0.0, 245.6] SR:0 DR:11 LR:-7.864 LO:21.56);ALT=T[chr12:110486232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110834302	+	chr12	110841409	+	.	11	0	5336560_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5336560_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110834302(+)-12:110841409(-)__12_110813501_110838501D;SPAN=7107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=A[chr12:110841409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110874503	+	chr12	110888059	+	.	12	0	5336592_1	20.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=5336592_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110874503(+)-12:110888059(-)__12_110887001_110912001D;SPAN=13556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:73 GQ:20 PL:[20.0, 0.0, 155.3] SR:0 DR:12 LR:-19.83 LO:26.06);ALT=A[chr12:110888059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110874988	+	chr12	110888063	+	.	8	0	5336593_1	2.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5336593_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110874988(+)-12:110888063(-)__12_110887001_110912001D;SPAN=13075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=G[chr12:110888063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110883357	+	chr12	110888059	+	.	97	35	5336594_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=13;MATEID=5336594_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110887001_110912001_322C;SPAN=4702;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:73 GQ:27 PL:[297.0, 27.0, 0.0] SR:35 DR:97 LR:-297.1 LO:297.1);ALT=C[chr12:110888059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110897668	+	chr12	110902911	+	.	0	35	5336626_1	91.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5336626_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110887001_110912001_380C;SPAN=5243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:90 GQ:91.1 PL:[91.1, 0.0, 127.4] SR:35 DR:0 LR:-91.15 LO:91.48);ALT=C[chr12:110902911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110897718	+	chr12	110905960	+	.	29	0	5336628_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5336628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110897718(+)-12:110905960(-)__12_110887001_110912001D;SPAN=8242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:82 GQ:73.7 PL:[73.7, 0.0, 123.2] SR:0 DR:29 LR:-73.51 LO:74.26);ALT=T[chr12:110905960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110903050	+	chr12	110905960	+	.	28	0	5336652_1	72.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5336652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110903050(+)-12:110905960(-)__12_110887001_110912001D;SPAN=2910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:73 GQ:72.8 PL:[72.8, 0.0, 102.5] SR:0 DR:28 LR:-72.65 LO:72.97);ALT=G[chr12:110905960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110906797	+	chr12	110922879	+	.	12	0	5336669_1	32.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5336669_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110906797(+)-12:110922879(-)__12_110887001_110912001D;SPAN=16082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:25 GQ:26.3 PL:[32.9, 0.0, 26.3] SR:0 DR:12 LR:-32.86 LO:32.86);ALT=G[chr12:110922879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110931038	+	chr12	110933817	+	.	10	43	5336320_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5336320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_110911501_110936501_213C;SPAN=2779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:101 GQ:99 PL:[128.0, 0.0, 114.8] SR:43 DR:10 LR:-127.8 LO:127.8);ALT=T[chr12:110933817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110931085	+	chr12	110939852	+	.	27	0	5336349_1	68.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5336349_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110931085(+)-12:110939852(-)__12_110936001_110961001D;SPAN=8767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:75 GQ:68.9 PL:[68.9, 0.0, 111.8] SR:0 DR:27 LR:-68.81 LO:69.4);ALT=T[chr12:110939852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110934034	+	chr12	110939815	+	.	69	0	5336352_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5336352_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110934034(+)-12:110939815(-)__12_110936001_110961001D;SPAN=5781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:40 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:0 DR:69 LR:-204.7 LO:204.7);ALT=G[chr12:110939815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	110937361	+	chr12	110939852	+	.	9	0	5336357_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5336357_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110937361(+)-12:110939852(-)__12_110936001_110961001D;SPAN=2491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:114 GQ:0.9 PL:[0.0, 0.9, 277.2] SR:0 DR:9 LR:1.176 LO:16.48);ALT=A[chr12:110939852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	111162569	+	chr12	111168330	+	.	2	3	5337131_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTAC;MAPQ=60;MATEID=5337131_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_111156501_111181501_279C;SPAN=5761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:75 GQ:6.9 PL:[0.0, 6.9, 194.7] SR:3 DR:2 LR:7.115 LO:6.623);ALT=C[chr12:111168330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	111169708	+	chr12	111180458	+	.	0	45	5337152_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5337152_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_111156501_111181501_70C;SPAN=10750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:88 GQ:88.4 PL:[124.7, 0.0, 88.4] SR:45 DR:0 LR:-125.0 LO:125.0);ALT=T[chr12:111180458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
