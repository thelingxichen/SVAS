chr12	22538191	+	chr13	45143367	+	.	25	0	7466498_1	58.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7466498_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:22538191(+)-13:45143367(-)__12_22515501_22540501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:91 GQ:58.1 PL:[58.1, 0.0, 160.4] SR:0 DR:25 LR:-57.87 LO:60.65);ALT=G[chr13:45143367[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	45143518	+	chr12	22538392	+	.	35	0	7466502_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=7466502_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:22538392(-)-13:45143518(+)__12_22515501_22540501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:51 GQ:19.4 PL:[101.9, 0.0, 19.4] SR:0 DR:35 LR:-104.6 LO:104.6);ALT=]chr13:45143518]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	22817754	+	chr12	22747188	+	.	60	17	7468278_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=7468278_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_22809501_22834501_245C;SPAN=70566;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:65 DP:111 GQ:82.4 PL:[184.7, 0.0, 82.4] SR:17 DR:60 LR:-186.5 LO:186.5);ALT=]chr12:22817754]T;VARTYPE=BND:DUP-th;JOINTYPE=th
