chr13	77236139	+	chr13	77238282	+	.	54	49	8164968_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGT;MAPQ=60;MATEID=8164968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_77224001_77249001_323C;SPAN=2143;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:76 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:49 DR:54 LR:-247.6 LO:247.6);ALT=T[chr13:77238282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	77573912	+	chr13	77389680	+	TTTTTCCTT	7	2	8166097_1	8.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TTTTTCCTT;MAPQ=60;MATEID=8166097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_77567001_77592001_315C;SPAN=184232;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:56 GQ:8 PL:[8.0, 0.0, 126.8] SR:2 DR:7 LR:-7.935 LO:14.3);ALT=]chr13:77573912]T;VARTYPE=BND:DUP-th;JOINTYPE=th
