chr4	78178805	+	chr4	79036036	-	.	20	0	2763125_1	53.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2763125_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:78178805(+)-4:79036036(+)__4_79012501_79037501D;SPAN=857231;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:47 GQ:53.3 PL:[53.3, 0.0, 59.9] SR:0 DR:20 LR:-53.29 LO:53.31);ALT=A]chr4:79036036];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	78179108	-	chr4	79035835	+	.	14	0	2763126_1	35.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=2763126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:78179108(-)-4:79035835(-)__4_79012501_79037501D;SPAN=856727;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:40 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:0 DR:14 LR:-35.38 LO:35.77);ALT=[chr4:79035835[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	79269134	+	chr4	79275196	+	.	86	28	2763514_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAGCTTCAAGATA;MAPQ=60;MATEID=2763514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_79257501_79282501_139C;SPAN=6062;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:168 GQ:99 PL:[274.7, 0.0, 132.8] SR:28 DR:86 LR:-277.3 LO:277.3);ALT=A[chr4:79275196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
