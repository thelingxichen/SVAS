chr3	197530842	-	chr3	197531958	+	.	11	0	2601715_1	2.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2601715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:197530842(-)-3:197531958(-)__3_197519001_197544001D;SPAN=1116;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:124 GQ:2.9 PL:[2.9, 0.0, 296.6] SR:0 DR:11 LR:-2.716 LO:20.73);ALT=[chr3:197531958[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
