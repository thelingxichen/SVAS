chr11	75112778	+	chr11	75115062	+	.	3	5	4921333_1	0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=29;MATEID=4921333_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_75092501_75117501_339C;SPAN=2284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:152 GQ:14.5 PL:[0.0, 14.5, 396.0] SR:5 DR:3 LR:14.77 LO:13.2);ALT=G[chr11:75115062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	75273365	+	chr11	75277358	+	.	3	2	4921687_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4921687_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_75264001_75289001_58C;SPAN=3993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:2 DR:3 LR:5.711 LO:8.577);ALT=G[chr11:75277358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	75526569	+	chr11	75562925	+	.	11	11	4922217_1	44.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4922217_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_75558001_75583001_372C;SPAN=36356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:11 DR:11 LR:-44.2 LO:44.37);ALT=G[chr11:75562925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	75591084	+	chr11	75622996	+	ATTCATGCCCGAAACCAAAATGAAATAATTTTTGGGCTGAATGATGGATACTATGGTGCTCCATTTGAACATA	2	17	4922367_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTCATGCCCGAAACCAAAATGAAATAATTTTTGGGCTGAATGATGGATACTATGGTGCTCCATTTGAACATA;MAPQ=60;MATEID=4922367_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_75582501_75607501_307C;SPAN=31912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:38 GQ:39.2 PL:[52.4, 0.0, 39.2] SR:17 DR:2 LR:-52.52 LO:52.52);ALT=G[chr11:75622996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
