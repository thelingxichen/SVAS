chr5	166383887	+	chr12	61302378	+	.	2	6	3908570_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATATATATATGTGTATATATATATA;MAPQ=60;MATEID=3908570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_166379501_166404501_370C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:11 GQ:3.8 PL:[20.3, 0.0, 3.8] SR:6 DR:2 LR:-20.51 LO:20.51);ALT=A[chr12:61302378[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	129465168	+	chr8	129471267	+	.	99	49	5692964_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CCAGCTTGTGTTTTT;MAPQ=60;MATEID=5692964_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_129458001_129483001_174C;SPAN=6099;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:126 DP:1021 GQ:99 PL:[139.7, 0.0, 2338.0] SR:49 DR:99 LR:-139.3 LO:256.6);ALT=T[chr8:129471267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	129762521	+	chr8	129766027	+	.	41	32	5694424_1	99.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=31;MATEID=5694424_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_8_129752001_129777001_64C;SPAN=3506;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:56 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:32 DR:41 LR:-194.7 LO:194.7);ALT=T[chr8:129766027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	130149176	+	chr12	60402590	-	.	23	29	5695657_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5695657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_130144001_130169001_40C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:29 DR:23 LR:-118.8 LO:118.8);ALT=T]chr12:60402590];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	60521845	+	chr12	60525052	+	TTTCTGTCC	129	91	7648145_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TTTCTGTCC;MAPQ=60;MATEID=7648145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_60515001_60540001_56C;SPAN=3207;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:179 DP:67 GQ:48.4 PL:[531.4, 48.4, 0.0] SR:91 DR:129 LR:-531.4 LO:531.4);ALT=A[chr12:60525052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
