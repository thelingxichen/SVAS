chr6	135363292	+	chr6	135375887	+	.	8	0	3037747_1	5.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3037747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:135363292(+)-6:135375887(-)__6_135362501_135387501D;SPAN=12595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:0 DR:8 LR:-5.276 LO:15.61);ALT=T[chr6:135375887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
