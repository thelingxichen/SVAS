chr1	95541860	-	chr1	95542934	+	.	8	0	425585_1	8.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=425585_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:95541860(-)-1:95542934(-)__1_95525501_95550501D;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:0 DR:8 LR:-8.798 LO:16.28);ALT=[chr1:95542934[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
