chr11	110150482	+	chr11	110167192	+	.	0	7	5000341_1	13.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5000341_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_110127501_110152501_161C;SPAN=16710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:36 GQ:13.4 PL:[13.4, 0.0, 72.8] SR:7 DR:0 LR:-13.35 LO:15.77);ALT=C[chr11:110167192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
