chr1	241677013	+	chr1	241680482	+	.	0	10	632959_1	6.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=632959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_241668001_241693001_297C;SPAN=3469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:10 DR:0 LR:-6.73 LO:19.53);ALT=T[chr1:241680482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	241680617	+	chr1	241682890	+	.	19	13	632970_1	57.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=632970_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_241668001_241693001_116C;SPAN=2273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:94 GQ:57.2 PL:[57.2, 0.0, 169.4] SR:13 DR:19 LR:-57.06 LO:60.23);ALT=C[chr1:241682890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
