chr8	61320517	-	chr8	61321517	+	.	9	0	3881613_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3881613_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:61320517(-)-8:61321517(-)__8_61299001_61324001D;SPAN=1000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=[chr8:61321517[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	61429815	+	chr8	61471408	+	.	0	23	3882053_1	62.0	.	EVDNC=ASSMB;HOMSEQ=CAGGTG;MAPQ=60;MATEID=3882053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_61470501_61495501_135C;SPAN=41593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:50 GQ:59 PL:[62.3, 0.0, 59.0] SR:23 DR:0 LR:-62.38 LO:62.38);ALT=G[chr8:61471408[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	61471484	+	chr8	61496766	+	GTAGAGTTCGGTGCTCGAATGATAACTATTGATGGGAAACAGATAAAACTTCAGATATGGGATAC	3	31	3882060_1	96.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GTAGAGTTCGGTGCTCGAATGATAACTATTGATGGGAAACAGATAAAACTTCAGATATGGGATAC;MAPQ=60;MATEID=3882060_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_61470501_61495501_294C;SPAN=25282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:46 GQ:14 PL:[96.5, 0.0, 14.0] SR:31 DR:3 LR:-99.86 LO:99.86);ALT=T[chr8:61496766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	61496850	+	chr8	61504415	+	AGAGATACATTCAACCACTTGACAACCTGGTTAGAAGATGCCCGCCAGCATTCCAATTCCAACATGGTCATTATGCTTATTGGAAATAAA	0	24	3882236_1	57.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGAGATACATTCAACCACTTGACAACCTGGTTAGAAGATGCCCGCCAGCATTCCAATTCCAACATGGTCATTATGCTTATTGGAAATAAA;MAPQ=60;MATEID=3882236_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_61495001_61520001_271C;SPAN=7565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:82 GQ:57.2 PL:[57.2, 0.0, 139.7] SR:24 DR:0 LR:-57.01 LO:59.01);ALT=G[chr8:61504415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	61531208	+	chr8	61533231	+	.	0	10	3882340_1	11.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3882340_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_61519501_61544501_160C;SPAN=2023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:0 LR:-11.34 LO:20.42);ALT=G[chr8:61533231[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
