chr9	90858996	+	chr9	90860964	+	.	124	58	4321638_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTATGTACCTTTT;MAPQ=60;MATEID=4321638_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_90846001_90871001_272C;SPAN=1968;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:44 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:58 DR:124 LR:-432.4 LO:432.4);ALT=T[chr9:90860964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	91003459	+	chr9	91041298	+	.	9	0	4322337_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4322337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:91003459(+)-9:91041298(-)__9_90993001_91018001D;SPAN=37839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:6 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=G[chr9:91041298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	91926267	+	chr9	91930084	+	.	40	38	4325178_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4325178_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_91924001_91949001_326C;SPAN=3817;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:87 GQ:9.5 PL:[200.9, 0.0, 9.5] SR:38 DR:40 LR:-211.2 LO:211.2);ALT=G[chr9:91930084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	91933528	+	chr9	91934565	+	.	34	7	4325206_1	93.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4325206_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_91924001_91949001_361C;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:93 GQ:93.8 PL:[93.8, 0.0, 130.1] SR:7 DR:34 LR:-93.64 LO:94.0);ALT=G[chr9:91934565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
