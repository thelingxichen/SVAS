chr2	146862621	+	chr2	146876863	+	.	0	111	1405239_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=1405239_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_2_146853001_146878001_79C;SPAN=14242;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:42 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:111 DR:0 LR:-326.8 LO:326.8);ALT=T[chr2:146876863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
