chr3	119431705	+	chr21	30382812	+	.	25	70	10743787_1	99.0	.	DISC_MAPQ=11;EVDNC=ASDIS;HOMSEQ=TCCCAGCTACTTGGGAGGCTGAG;MAPQ=32;MATEID=10743787_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_30380001_30405001_438C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:63 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:70 DR:25 LR:-241.0 LO:241.0);ALT=G[chr21:30382812[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
