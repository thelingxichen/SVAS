chr21	9834344	+	chr21	9835501	+	.	0	63	7102480_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GA;MAPQ=60;MATEID=7102480_2;MATENM=3;NM=3;NUMPARTS=2;SCTG=c_21_9824501_9849501_567C;SPAN=1157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:244 GQ:99 PL:[142.0, 0.0, 449.0] SR:63 DR:0 LR:-141.9 LO:150.8);ALT=A[chr21:9835501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	10815200	+	chr21	10810640	+	.	12	0	7108949_1	0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7108949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:10810640(-)-21:10815200(+)__21_10804501_10829501D;SPAN=4560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:249 GQ:27.7 PL:[0.0, 27.7, 660.1] SR:0 DR:12 LR:27.85 LO:19.33);ALT=]chr21:10815200]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	11122404	+	chrX	858670	+	.	2	33	7112222_1	0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=GGCCATTATTCTGTCTCCCACATGGG;MAPQ=19;MATEID=7112222_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_21_11098501_11123501_378C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:35 DP:444 GQ:4.4 PL:[0.0, 4.4, 1086.0] SR:33 DR:2 LR:4.756 LO:64.08);ALT=G[chrX:858670[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chrX	545941	+	chrX	544617	+	.	10	0	7346516_1	17.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=7346516_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:544617(-)-23:545941(+)__23_539001_564001D;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=]chrX:545941]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	901072	+	chrX	899396	+	.	27	0	7347442_1	76.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=7347442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:899396(-)-23:901072(+)__23_882001_907001D;SPAN=1676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:46 GQ:33.8 PL:[76.7, 0.0, 33.8] SR:0 DR:27 LR:-77.51 LO:77.51);ALT=]chrX:901072]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	1340220	+	chrX	1337548	+	.	16	0	7348034_1	34.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=7348034_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1337548(-)-23:1340220(+)__23_1323001_1348001D;SPAN=2672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:67 GQ:34.7 PL:[34.7, 0.0, 127.1] SR:0 DR:16 LR:-34.66 LO:37.67);ALT=]chrX:1340220]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	1338719	+	chrX	1337635	+	.	11	0	7348035_1	20.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7348035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1337635(-)-23:1338719(+)__23_1323001_1348001D;SPAN=1084;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:58 GQ:20.6 PL:[20.6, 0.0, 119.6] SR:0 DR:11 LR:-20.6 LO:24.64);ALT=]chrX:1338719]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	1360542	+	chrX	1551603	+	.	3	11	7348092_1	35.0	.	DISC_MAPQ=26;EVDNC=TSI_L;HOMSEQ=TCCCAGCTACTCGGGAGGCTGAGGCAGGAGAATCGCTTGAACCC;MAPQ=60;MATEID=7348092_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_23_1347501_1372501_81C;SPAN=191061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:38 GQ:35.9 PL:[35.9, 0.0, 55.7] SR:11 DR:3 LR:-35.92 LO:36.17);ALT=C[chrX:1551603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1387810	+	chrX	1401569	+	.	8	0	7348812_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7348812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1387810(+)-23:1401569(-)__23_1372001_1397001D;SPAN=13759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=G[chrX:1401569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1387817	+	chrX	1393643	+	.	15	0	7348814_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7348814_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1387817(+)-23:1393643(-)__23_1372001_1397001D;SPAN=5826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:0 DR:15 LR:-34.89 LO:36.48);ALT=C[chrX:1393643[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1401672	+	chrX	1404670	+	.	0	10	7348186_1	19.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7348186_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1396501_1421501_275C;SPAN=2998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:50 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:10 DR:0 LR:-19.46 LO:22.66);ALT=G[chrX:1404670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1453443	+	chrX	1450040	+	.	29	8	7348364_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;HOMSEQ=GCCACTGCACTCCAGCCTGGGTGACAGAGGAAGACTCCATCTCAAAAAAAAAAAAAAAA;MAPQ=60;MATEID=7348364_2;MATENM=4;NM=6;NUMPARTS=2;SCTG=c_23_1445501_1470501_102C;SPAN=3403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:53 GQ:18.8 PL:[107.9, 0.0, 18.8] SR:8 DR:29 LR:-111.1 LO:111.1);ALT=]chrX:1453443]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	1455819	+	chrX	1460619	+	.	0	24	7348399_1	60.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7348399_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_1445501_1470501_80C;SPAN=4800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:71 GQ:60.2 PL:[60.2, 0.0, 109.7] SR:24 DR:0 LR:-59.99 LO:60.86);ALT=G[chrX:1460619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1455830	+	chrX	1464206	+	.	20	0	7348400_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7348400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1455830(+)-23:1464206(-)__23_1445501_1470501D;SPAN=8376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:66 GQ:48.2 PL:[48.2, 0.0, 110.9] SR:0 DR:20 LR:-48.14 LO:49.55);ALT=C[chrX:1464206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1460722	+	chrX	1467323	+	ATCCAAACCCACCAATCACGAACCTAAGGATGAAAGCAAAGGCTCAGCAGTTGACCTGGGACCTTAACAGAAATGTGACCGATATCGAGTGTGTTAAAGACGCCGACTATTCTATGCC	0	32	7348412_1	89.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATCCAAACCCACCAATCACGAACCTAAGGATGAAAGCAAAGGCTCAGCAGTTGACCTGGGACCTTAACAGAAATGTGACCGATATCGAGTGTGTTAAAGACGCCGACTATTCTATGCC;MAPQ=60;MATEID=7348412_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_1445501_1470501_320C;SPAN=6601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:59 GQ:53.3 PL:[89.6, 0.0, 53.3] SR:32 DR:0 LR:-90.14 LO:90.14);ALT=G[chrX:1467323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1479407	+	chrX	1478336	+	.	13	0	7348135_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7348135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1478336(-)-23:1479407(+)__23_1470001_1495001D;SPAN=1071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:45 GQ:30.8 PL:[30.8, 0.0, 77.0] SR:0 DR:13 LR:-30.72 LO:31.88);ALT=]chrX:1479407]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	1487597	+	chrX	1495998	+	.	8	0	7348283_1	23.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7348283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1487597(+)-23:1495998(-)__23_1494501_1519501D;SPAN=8401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:5 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=T[chrX:1495998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1499999	+	chrX	1501283	+	.	0	7	7348293_1	7.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7348293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1494501_1519501_155C;SPAN=1284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:59 GQ:7.1 PL:[7.1, 0.0, 135.8] SR:7 DR:0 LR:-7.123 LO:14.13);ALT=T[chrX:1501283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1506313	+	chrX	1508133	+	.	10	17	7348312_1	64.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=7348312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1494501_1519501_59C;SPAN=1820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:56 GQ:64.1 PL:[64.1, 0.0, 70.7] SR:17 DR:10 LR:-64.05 LO:64.08);ALT=C[chrX:1508133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1508623	+	chrX	1510790	+	.	0	102	7348317_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=7348317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1494501_1519501_51C;SPAN=2167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:220 GQ:99 PL:[277.1, 0.0, 257.3] SR:102 DR:0 LR:-277.1 LO:277.1);ALT=G[chrX:1510790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1561211	+	chrX	1571640	+	.	0	17	7348841_1	50.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=7348841_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1568001_1593001_130C;SPAN=10429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:22 GQ:0.8 PL:[50.3, 0.0, 0.8] SR:17 DR:0 LR:-52.61 LO:52.61);ALT=C[chrX:1571640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1710652	+	chrX	1712335	+	.	8	0	7349200_1	15.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7349200_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1710652(+)-23:1712335(-)__23_1690501_1715501D;SPAN=1683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=G[chrX:1712335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1713119	+	chrX	1714274	+	.	5	5	7349204_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGGT;MAPQ=60;MATEID=7349204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_1690501_1715501_170C;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:5 DR:5 LR:-17.25 LO:20.3);ALT=T[chrX:1714274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1842602	-	chrX	1843673	+	.	8	0	7349760_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7349760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1842602(-)-23:1843673(-)__23_1837501_1862501D;SPAN=1071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:0 DR:8 LR:-9.34 LO:16.4);ALT=[chrX:1843673[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	2527523	+	chrX	2530191	+	GCTGACTTTGACTTAGCGATGCCTTTCCTGATGGAGGAAACA	14	15	7351005_1	59.0	.	DISC_MAPQ=46;EVDNC=TSI_G;HOMSEQ=GTGA;INSERTION=GCTGACTTTGACTTAGCGATGCCTTTCCTGATGGAGGAAACA;MAPQ=60;MATEID=7351005_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_2523501_2548501_122C;SPAN=2668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:48 GQ:56.3 PL:[59.6, 0.0, 56.3] SR:15 DR:14 LR:-59.62 LO:59.62);ALT=G[chrX:2530191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2527523	+	chrX	2529036	+	.	4	7	7351004_1	14.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=7351004_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_23_2523501_2548501_122C;SPAN=1513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:7 DR:4 LR:-14.76 LO:17.85);ALT=G[chrX:2529036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2527545	+	chrX	2533855	+	.	10	0	7351006_1	17.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=7351006_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:2527545(+)-23:2533855(-)__23_2523501_2548501D;SPAN=6310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:0 DR:10 LR:-17.57 LO:22.03);ALT=G[chrX:2533855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2530261	+	chrX	2533856	+	.	0	12	7351012_1	24.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7351012_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_2523501_2548501_214C;SPAN=3595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:12 DR:0 LR:-24.71 LO:27.71);ALT=T[chrX:2533856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2609468	+	chrX	2635645	+	ATGGTGGTTTCGATTTATCCGATGCCCTTCCT	51	19	7351434_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATGGTGGTTTCGATTTATCCGATGCCCTTCCT;MAPQ=60;MATEID=7351434_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_2597001_2622001_57C;SPAN=26177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:70 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:19 DR:51 LR:-208.0 LO:208.0);ALT=G[chrX:2635645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2638468	+	chrX	2640667	+	.	2	86	7351523_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGTA;MAPQ=60;MATEID=7351523_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_2621501_2646501_259C;SPAN=2199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:141 GQ:94.1 PL:[245.9, 0.0, 94.1] SR:86 DR:2 LR:-249.2 LO:249.2);ALT=A[chrX:2640667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2640716	+	chrX	2656240	+	AAAAGGAGGCAGTGATGGTGGAGGCAGCCACAGGAAAGAAGGGGAAGAGGCCGACGCCCCAGGCGTGATCCCCGGGATTGTGGGGGCTGTCGTGGTCGCCGTGGCTGGAGCCATCTCTAGCTTCATTGCTTACCAGAAAAAGAAGCTATGCTTCAAAGAAAAT	3	80	7351529_1	99.0	.	DISC_MAPQ=43;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AAAAGGAGGCAGTGATGGTGGAGGCAGCCACAGGAAAGAAGGGGAAGAGGCCGACGCCCCAGGCGTGATCCCCGGGATTGTGGGGGCTGTCGTGGTCGCCGTGGCTGGAGCCATCTCTAGCTTCATTGCTTACCAGAAAAAGAAGCTATGCTTCAAAGAAAAT;MAPQ=60;MATEID=7351529_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_2621501_2646501_265C;SPAN=15524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:55 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:80 DR:3 LR:-237.7 LO:237.7);ALT=G[chrX:2656240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2644414	+	chrX	2656240	+	.	3	19	7351562_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=7351562_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_23_2646001_2671001_9C;SPAN=11826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:39 GQ:42.2 PL:[52.1, 0.0, 42.2] SR:19 DR:3 LR:-52.2 LO:52.2);ALT=G[chrX:2656240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2644465	+	chrX	2658817	+	.	14	0	7351563_1	37.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7351563_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:2644465(+)-23:2658817(-)__23_2646001_2671001D;SPAN=14352;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:34 GQ:37.1 PL:[37.1, 0.0, 43.7] SR:0 DR:14 LR:-37.0 LO:37.05);ALT=A[chrX:2658817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2656297	+	chrX	2658819	+	.	14	17	7351583_1	84.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=7351583_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_23_2646001_2671001_9C;SPAN=2522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:65 GQ:71.6 PL:[84.8, 0.0, 71.6] SR:17 DR:14 LR:-84.77 LO:84.77);ALT=G[chrX:2658819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2840067	+	chrX	2843657	+	.	0	7	7351933_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7351933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_2842001_2867001_299C;SPAN=3590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:20 GQ:17.6 PL:[17.6, 0.0, 30.8] SR:7 DR:0 LR:-17.69 LO:17.88);ALT=T[chrX:2843657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2843810	+	chrX	2847272	+	.	9	1	7351937_1	17.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=CCTGG;MAPQ=19;MATEID=7351937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_2842001_2867001_201C;SPAN=3462;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:1 DR:9 LR:-17.25 LO:20.3);ALT=G[chrX:2847272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	3351470	-	chrY	7431135	+	.	17	11	7563710_1	66.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTAAGGTCATG;MAPQ=45;MATEID=7563710_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_24_7423501_7448501_5C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:9 GQ:6 PL:[66.0, 6.0, 0.0] SR:11 DR:17 LR:-66.02 LO:66.02);ALT=[chrY:7431135[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
