chr17	76282255	+	chr17	76283431	+	.	57	23	9827894_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCAGCCTGGCCAACATGGT;MAPQ=60;MATEID=9827894_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_76268501_76293501_55C;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:25 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:23 DR:57 LR:-221.2 LO:221.2);ALT=T[chr17:76283431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
