chr10	114136208	+	chr10	114154675	+	.	0	7	4692686_1	14.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=4692686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_114145501_114170501_187C;SPAN=18467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:34 GQ:14 PL:[14.0, 0.0, 66.8] SR:7 DR:0 LR:-13.9 LO:15.96);ALT=T[chr10:114154675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	114205410	+	chr10	114206461	+	.	10	12	4692739_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4692739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_114194501_114219501_184C;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:55 GQ:47.9 PL:[47.9, 0.0, 84.2] SR:12 DR:10 LR:-47.82 LO:48.41);ALT=T[chr10:114206461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	114207225	+	chr10	114220282	+	.	3	5	4692763_1	20.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4692763_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_114219001_114244001_80C;SPAN=13057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:5 DR:3 LR:-19.91 LO:20.23);ALT=G[chr10:114220282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
