chr1	32738250	+	chr1	46281894	+	.	2	34	231253_1	92.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=AGAGAGAGAGAGAGAGAGAGAG;MAPQ=60;MATEID=231253_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46280501_46305501_65C;SPAN=13543644;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:74 GQ:85.7 PL:[92.3, 0.0, 85.7] SR:34 DR:2 LR:-92.19 LO:92.19);ALT=G[chr1:46281894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33270900	+	chr8	125445125	+	.	0	9	5674648_1	16.0	.	EVDNC=ASSMB;HOMSEQ=GAGAGGGAGAGAGGGAGAG;MAPQ=60;MATEID=5674648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_125440001_125465001_21C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:9 DR:0 LR:-16.16 LO:19.94);ALT=G[chr8:125445125[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	33476428	+	chr2	32048478	+	.	11	0	170267_1	15.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=170267_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:33476428(+)-2:32048478(-)__1_33467001_33492001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:0 DR:11 LR:-15.45 LO:23.15);ALT=T[chr2:32048478[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	34471261	-	chr1	34473077	+	.	10	0	174575_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=174575_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:34471261(-)-1:34473077(-)__1_34447001_34472001D;SPAN=1816;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:66 GQ:15.2 PL:[15.2, 0.0, 143.9] SR:0 DR:10 LR:-15.13 LO:21.33);ALT=[chr1:34473077[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	77859321	+	chr1	35007076	+	.	9	0	177283_1	21.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=177283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:35007076(-)-10:77859321(+)__1_34986001_35011001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:29 GQ:21.8 PL:[21.8, 0.0, 48.2] SR:0 DR:9 LR:-21.85 LO:22.41);ALT=]chr10:77859321]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	46195367	+	chr1	46123932	+	.	85	34	231844_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTTT;MAPQ=60;MATEID=231844_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46182501_46207501_386C;SPAN=71435;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:73 GQ:27 PL:[297.0, 27.0, 0.0] SR:34 DR:85 LR:-297.1 LO:297.1);ALT=]chr1:46195367]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	17459958	+	chr1	46673196	+	.	10	61	10193454_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;HOMSEQ=TTTTCTTTCTTTCTTTCTTTCTTT;MAPQ=3;MATEID=10193454_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_19_17444001_17469001_202C;SPAN=-1;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:61 DP:33 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:61 DR:10 LR:-178.2 LO:178.2);ALT=]chr19:17459958]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	87051452	+	chr13	96262340	-	.	27	0	8243528_1	12.0	.	DISC_MAPQ=22;EVDNC=TSI_L;HOMSEQ=CACACACACACACACACACACACACACACAC;MAPQ=60;MATEID=8243528_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACACACACACACACACACACACACACACA;SCTG=c_13_96260501_96285501_137C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:97 GQ:12.6 PL:[12.6, 0.0, 58.1] SR:0 DR:27 LR:-11.46 LO:14.86);ALT=C]chr13:96262340];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr13	49371052	+	chr1	87512434	+	.	33	0	401572_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=401572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:87512434(-)-13:49371052(+)__1_87489501_87514501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:33 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:0 DR:33 LR:-99.02 LO:99.02);ALT=]chr13:49371052]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	101237235	+	chr12	6407650	+	.	30	132	7360941_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=7360941_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_12_6394501_6419501_132C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:140 DP:48 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:132 DR:30 LR:-415.9 LO:415.9);ALT=A[chr12:6407650[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	155713283	+	chr20	44237876	+	ACGAGACT	0	8	10568415_1	1.0	.	EVDNC=ASSMB;INSERTION=ACGAGACT;MAPQ=60;MATEID=10568415_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_44222501_44247501_11C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:8 DR:0 LR:-1.212 LO:14.96);ALT=G[chr20:44237876[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	155749846	-	chr1	155750998	+	.	8	0	563835_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=563835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155749846(-)-1:155750998(-)__1_155746501_155771501D;SPAN=1152;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:139 GQ:11.1 PL:[0.0, 11.1, 359.7] SR:0 DR:8 LR:11.25 LO:13.52);ALT=[chr1:155750998[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	156526723	+	chr1	156528936	+	.	139	66	568044_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAATTGAGTAGCTCAGC;MAPQ=60;MATEID=568044_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_1_156506001_156531001_249C;SPAN=2213;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:168 DP:40 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:66 DR:139 LR:-498.4 LO:498.4);ALT=C[chr1:156528936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156705379	+	chr14	61033233	+	.	12	0	569583_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=569583_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156705379(+)-14:61033233(-)__1_156702001_156727001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:12 DP:11 GQ:3 PL:[33.0, 3.0, 0.0] SR:0 DR:12 LR:-33.01 LO:33.01);ALT=T[chr14:61033233[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	200577714	-	chr1	200579528	+	.	8	1	748458_1	0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CTCAGGAG;MAPQ=49;MATEID=748458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_200557001_200582001_396C;SPAN=1814;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:175 GQ:17.5 PL:[0.0, 17.5, 458.8] SR:1 DR:8 LR:17.7 LO:14.76);ALT=[chr1:200579528[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	200693890	-	chr12	7108122	+	.	10	0	7364967_1	18.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=7364967_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:200693890(-)-12:7108122(-)__12_7105001_7130001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:0 DR:10 LR:-18.65 LO:22.38);ALT=[chr12:7108122[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	201452924	+	chr1	201450401	+	.	9	73	752453_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGGGC;MAPQ=60;MATEID=752453_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_201439001_201464001_296C;SPAN=2523;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:74 DP:310 GQ:99 PL:[160.3, 0.0, 592.7] SR:73 DR:9 LR:-160.3 LO:174.2);ALT=]chr1:201452924]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	203040565	+	chrX	52961551	+	.	4	40	760370_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCCGCCTCGGCCTCCCAAAGTGC;MAPQ=60;MATEID=760370_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_203031501_203056501_184C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:40 DR:4 LR:-128.7 LO:128.7);ALT=C[chrX:52961551[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	236549103	+	chr1	236551330	+	.	45	27	866535_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TAATAATTTGAAAGTTA;MAPQ=60;MATEID=866535_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_236547501_236572501_205C;SPAN=2227;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:14 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:27 DR:45 LR:-178.2 LO:178.2);ALT=A[chr1:236551330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	237449857	-	chr5	35747707	+	TGGTATATGATA	12	40	3368285_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TGGTATATGATA;MAPQ=60;MATEID=3368285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_35745501_35770501_86C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:77 GQ:61.7 PL:[124.4, 0.0, 61.7] SR:40 DR:12 LR:-125.5 LO:125.5);ALT=[chr5:35747707[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	38570669	+	chr1	242480401	+	.	0	8	6209223_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CTGGGT;MAPQ=60;MATEID=6209223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_38563001_38588001_376C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:8 DR:0 LR:-9.882 LO:16.52);ALT=]chr10:38570669]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	243127797	+	chr1	243129216	+	.	38	59	879143_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=GCCTCCCAAAGTGCTGGGATTACAGG;MAPQ=60;MATEID=879143_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_1_243113501_243138501_303C;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:13 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:59 DR:38 LR:-257.5 LO:257.5);ALT=G[chr1:243129216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	245784989	+	chr1	245826805	+	.	72	25	884813_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=884813_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_245759501_245784501_350C;SPAN=41816;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:0 GQ:24 PL:[264.0, 24.0, 0.0] SR:25 DR:72 LR:-264.1 LO:264.1);ALT=G[chr1:245826805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246402504	+	chr11	93394098	+	.	7	19	7104531_1	16.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TAAC;MAPQ=60;MATEID=7104531_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_93394001_93419001_361C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:197 GQ:16 PL:[16.0, 0.0, 461.6] SR:19 DR:7 LR:-15.95 LO:41.34);ALT=C[chr11:93394098[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	247254725	+	chr1	247260676	+	.	35	32	887837_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=A;MAPQ=26;MATEID=887837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_247229501_247254501_66C;SPAN=5951;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:0 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:32 DR:35 LR:-171.6 LO:171.6);ALT=A[chr1:247260676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	247850475	+	chr1	247856516	+	.	57	49	889935_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GAAAAGAAAGATC;MAPQ=60;MATEID=889935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_247842001_247867001_83C;SPAN=6041;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:28 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:49 DR:57 LR:-260.8 LO:260.8);ALT=C[chr1:247856516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	248051492	+	chr1	248057639	+	.	0	48	890052_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GCATGTATTTATTT;MAPQ=60;MATEID=890052_2;MATENM=5;NM=2;NUMPARTS=2;SCTG=c_1_248038001_248063001_112C;SPAN=6147;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:18 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:48 DR:0 LR:-141.9 LO:141.9);ALT=T[chr1:248057639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	189904	+	chr2	11984	+	.	8	0	6618601_1	0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6618601_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:11984(-)-11:189904(+)__11_171501_196501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:206 GQ:29.2 PL:[0.0, 29.2, 557.8] SR:0 DR:8 LR:29.4 LO:12.13);ALT=]chr11:189904]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	145554076	+	chr2	13428658	+	.	18	28	917360_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=ATATATATATATCCATATATATATATATCCATATATATATAT;MAPQ=19;MATEID=917360_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_13426001_13451001_269C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:34 DP:14 GQ:9 PL:[99.0, 9.0, 0.0] SR:28 DR:18 LR:-99.02 LO:99.02);ALT=]chr5:145554076]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	13534878	-	chr15	20609634	+	.	86	0	8759683_1	99.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=8759683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:13534878(-)-15:20609634(-)__15_20604501_20629501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:86 DP:192 GQ:99 PL:[232.1, 0.0, 232.1] SR:0 DR:86 LR:-231.9 LO:231.9);ALT=[chr15:20609634[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	13535069	+	chr15	20609518	-	.	30	0	8759685_1	34.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=8759685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:13535069(+)-15:20609518(+)__15_20604501_20629501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:238 GQ:34.6 PL:[34.6, 0.0, 542.9] SR:0 DR:30 LR:-34.55 LO:61.38);ALT=T]chr15:20609518];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chrX	56782687	+	chr2	31727422	+	.	12	5	11186115_1	37.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=TTAATGGGTGCAGCACACCAGCATGGCACATGTATACATATGTAACTAACCTGC;MAPQ=60;MATEID=11186115_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_23_56766501_56791501_173C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:70 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:5 DR:12 LR:-37.15 LO:40.17);ALT=]chrX:56782687]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	31816805	+	chr4	52742341	+	.	2	21	953551_1	66.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CAACAATGATAGACTGGATCAAGAAAATGCGGCACATATACA;MAPQ=60;MATEID=953551_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_31801001_31826001_126C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:23 DP:15 GQ:6 PL:[66.0, 6.0, 0.0] SR:21 DR:2 LR:-66.02 LO:66.02);ALT=A[chr4:52742341[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	32048486	+	chr12	53344194	-	.	3	23	7614893_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTGACTCTAAAATCATCAGCAG;MAPQ=60;MATEID=7614893_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_12_53336501_53361501_378C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:59 GQ:69.8 PL:[69.8, 0.0, 73.1] SR:23 DR:3 LR:-69.84 LO:69.85);ALT=G]chr12:53344194];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	34523656	+	chr2	34525720	+	.	59	49	959505_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=959505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_34520501_34545501_178C;SPAN=2064;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:18 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:49 DR:59 LR:-244.3 LO:244.3);ALT=G[chr2:34525720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39529128	+	chr2	34577789	+	.	10	0	10289780_1	22.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=10289780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:34577789(-)-19:39529128(+)__19_39518501_39543501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:41 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-21.9 LO:23.65);ALT=]chr19:39529128]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	34732900	+	chr6	78560888	+	.	11	38	959924_1	99.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=ACTTTTACACTGTTGGTGGGACTGTAAACTAGTTCAA;MAPQ=60;MATEID=959924_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_34716501_34741501_120C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:46 DP:12 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:38 DR:11 LR:-135.3 LO:135.3);ALT=A[chr6:78560888[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	34797628	+	chr2	34801577	+	.	67	43	960664_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAAATTATTATGTTTT;MAPQ=60;MATEID=960664_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_34790001_34815001_106C;SPAN=3949;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:31 GQ:24 PL:[264.0, 24.0, 0.0] SR:43 DR:67 LR:-264.1 LO:264.1);ALT=T[chr2:34801577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	35154964	-	chr12	114891197	+	.	16	0	960442_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=960442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:35154964(-)-12:114891197(-)__2_35133001_35158001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:26 GQ:16.1 PL:[45.8, 0.0, 16.1] SR:0 DR:16 LR:-46.47 LO:46.47);ALT=[chr12:114891197[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	98465797	+	chr2	35879336	+	.	10	0	5935138_1	2.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5935138_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:35879336(-)-9:98465797(+)__9_98441001_98466001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:113 GQ:2.6 PL:[2.6, 0.0, 269.9] SR:0 DR:10 LR:-2.396 LO:18.83);ALT=]chr9:98465797]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	35879355	+	chr9	98459861	+	GA	29	39	5935140_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GA;MAPQ=60;MATEID=5935140_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_98441001_98466001_230C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:52 DP:43 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:39 DR:29 LR:-151.8 LO:151.8);ALT=A[chr9:98459861[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	35976017	+	chr2	35997129	+	.	32	0	961928_1	92.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=961928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:35976017(+)-2:35997129(-)__2_35966001_35991001D;SPAN=21112;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:32 DP:8 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=C[chr2:35997129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	36892138	+	chr2	36893356	-	.	8	0	963437_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=963437_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:36892138(+)-2:36893356(+)__2_36872501_36897501D;SPAN=1218;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=G]chr2:36893356];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	37439980	-	chr10	12791579	+	.	9	32	6094665_1	99.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6094665_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_12789001_12814001_8C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:54 GQ:15.2 PL:[114.2, 0.0, 15.2] SR:32 DR:9 LR:-118.2 LO:118.2);ALT=[chr10:12791579[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr18	47337315	+	chr2	41973164	+	.	28	39	10015848_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;MAPQ=51;MATEID=10015848_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_47334001_47359001_171C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:62 DP:20 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:39 DR:28 LR:-181.5 LO:181.5);ALT=]chr18:47337315]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	42346259	+	chr2	42347319	+	TGTA	80	57	975230_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTA;MAPQ=60;MATEID=975230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_42336001_42361001_67C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:35 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:57 DR:80 LR:-333.4 LO:333.4);ALT=C[chr2:42347319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42775951	-	chr6	26807953	+	.	8	13	4093295_1	39.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=TATATATATATATATATAT;MAPQ=42;MATEID=4093295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_26803001_26828001_286C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:14 DP:9 GQ:3.6 PL:[39.6, 3.6, 0.0] SR:13 DR:8 LR:-39.61 LO:39.61);ALT=[chr6:26807953[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	125432159	+	chr2	71266069	+	.	10	0	1079314_1	15.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=1079314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:71266069(-)-3:125432159(+)__2_71246001_71271001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:66 GQ:15.2 PL:[15.2, 0.0, 143.9] SR:0 DR:10 LR:-15.13 LO:21.33);ALT=]chr3:125432159]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	21687096	+	chr2	115833867	+	.	37	56	1278196_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=1278196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_115811501_115836501_352C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:67 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:56 DR:37 LR:-241.0 LO:241.0);ALT=]chr19:21687096]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	116751295	+	chr2	116752836	-	.	8	0	1281409_1	0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=1281409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:116751295(+)-2:116752836(+)__2_116742501_116767501D;SPAN=1541;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:160 GQ:16.9 PL:[0.0, 16.9, 422.5] SR:0 DR:8 LR:16.94 LO:13.02);ALT=G]chr2:116752836];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	116974340	-	chr2	116981887	+	ACT	95	94	1282267_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ACT;MAPQ=60;MATEID=1282267_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_72C;SPAN=7547;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:183 DP:194 GQ:52.3 PL:[574.3, 52.3, 0.0] SR:94 DR:95 LR:-574.3 LO:574.3);ALT=[chr2:116981887[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	116974634	+	chr2	116978304	+	.	115	128	1282271_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1282271_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_379C;SPAN=3670;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:195 DP:131 GQ:52.6 PL:[577.6, 52.6, 0.0] SR:128 DR:115 LR:-577.6 LO:577.6);ALT=T[chr2:116978304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	116978299	+	chr2	116982310	-	.	99	82	1282293_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATA;MAPQ=60;MATEID=1282293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_384C;SPAN=4011;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:158 DP:96 GQ:42.7 PL:[468.7, 42.7, 0.0] SR:82 DR:99 LR:-468.7 LO:468.7);ALT=A]chr2:116982310];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	117797364	+	chr5	43904163	+	.	11	35	3402355_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAAAA;MAPQ=60;MATEID=3402355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_43904001_43929001_18C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:72 GQ:73.1 PL:[99.5, 0.0, 73.1] SR:35 DR:11 LR:-99.5 LO:99.5);ALT=A[chr5:43904163[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	118035938	+	chr7	52744989	+	.	2	21	4812393_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATATATATATA;MAPQ=60;MATEID=4812393_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_52724001_52749001_164C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:41 GQ:35.3 PL:[61.7, 0.0, 35.3] SR:21 DR:2 LR:-61.81 LO:61.81);ALT=A[chr7:52744989[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	102085249	+	chr2	120149146	+	GCACCTCAGCCTCCTGACCAGCTGGGATTACAGACATTCACCACAGAGCCTGGCTAATT	4	70	2803798_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;INSERTION=GCACCTCAGCCTCCTGACCAGCTGGGATTACAGACATTCACCACAGAGCCTGGCTAATT;MAPQ=60;MATEID=2803798_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_4_102067001_102092001_26C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:25 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:70 DR:4 LR:-214.6 LO:214.6);ALT=]chr4:102085249]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	144594741	+	chr14	58392234	+	.	3	9	1397172_1	30.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=AGGGAGGGAGGGAGGGAGGGAGGGAGGGAGG;MAPQ=18;MATEID=1397172_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_144574501_144599501_324C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:23 GQ:23.6 PL:[30.2, 0.0, 23.6] SR:9 DR:3 LR:-30.1 LO:30.1);ALT=G[chr14:58392234[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	156528004	-	chr9	32074060	+	ACAACTCAATA	16	37	1442054_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ACAACTCAATA;MAPQ=60;MATEID=1442054_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_156506001_156531001_130C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:63 GQ:19.4 PL:[131.6, 0.0, 19.4] SR:37 DR:16 LR:-136.0 LO:136.0);ALT=[chr9:32074060[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	156528145	+	chr7	81674028	+	.	18	0	5004205_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5004205_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:156528145(+)-7:81674028(-)__7_81658501_81683501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:56 GQ:44.3 PL:[44.3, 0.0, 90.5] SR:0 DR:18 LR:-44.25 LO:45.16);ALT=C[chr7:81674028[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	166014695	+	chr2	166016745	+	.	65	57	1478569_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=1478569_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_166012001_166037001_100C;SPAN=2050;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:108 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:57 DR:65 LR:-319.6 LO:319.6);ALT=G[chr2:166016745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	166888737	+	chr18	47205588	-	.	7	93	1482155_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACACACACACACACACACACACACA;MAPQ=60;MATEID=1482155_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_166869501_166894501_307C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:112 GQ:23.4 PL:[316.8, 23.4, 0.0] SR:93 DR:7 LR:-317.9 LO:317.9);ALT=A]chr18:47205588];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	167844961	+	chr2	167851209	+	.	117	57	1486242_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAACTTTA;MAPQ=60;MATEID=1486242_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_167825001_167850001_285C;SPAN=6248;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:154 DP:18 GQ:41.5 PL:[455.5, 41.5, 0.0] SR:57 DR:117 LR:-455.5 LO:455.5);ALT=A[chr2:167851209[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	168732575	+	chr22	43588630	-	.	3	3	10900302_1	14.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TATATATATATACGTATATATATATATATACGTGTATATATATATA;MAPQ=50;MATEID=10900302_2;MATENM=2;NM=1;NUMPARTS=3;SCTG=c_22_43585501_43610501_124C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:5 DP:7 GQ:1.4 PL:[14.6, 0.0, 1.4] SR:3 DR:3 LR:-15.11 LO:15.11);ALT=A]chr22:43588630];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	184345149	-	chr16	78078573	+	.	9	0	1553695_1	13.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1553695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:184345149(-)-16:78078573(-)__2_184338001_184363001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:61 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.18 LO:19.08);ALT=[chr16:78078573[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	184569178	+	chr2	184572010	-	.	57	61	1554454_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1554454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_184558501_184583501_152C;SPAN=2832;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:114 GQ:17.4 PL:[310.2, 17.4, 0.0] SR:61 DR:57 LR:-315.3 LO:315.3);ALT=C]chr2:184572010];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	184569193	-	chr2	184571029	+	.	66	44	1554455_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCCTG;MAPQ=60;MATEID=1554455_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_184558501_184583501_345C;SPAN=1836;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:89 DP:129 GQ:54.2 PL:[258.8, 0.0, 54.2] SR:44 DR:66 LR:-266.4 LO:266.4);ALT=[chr2:184571029[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	184584620	-	chrX	48822177	+	.	12	0	11149701_1	29.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=11149701_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:184584620(-)-23:48822177(-)__23_48804001_48829001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=[chrX:48822177[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	195455806	+	chr2	188649900	+	.	29	39	1569923_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGCCTCCCAAAGTGCTGGGATTACAGGCGTGAGCCACCGC;MAPQ=60;MATEID=1569923_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_188625501_188650501_1C;SPAN=6805906;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:62 DP:51 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:39 DR:29 LR:-181.5 LO:181.5);ALT=]chr2:195455806]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	194007524	+	chr18	66610044	-	.	9	0	10050157_1	21.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=10050157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:194007524(+)-18:66610044(+)__18_66591001_66616001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:29 GQ:21.8 PL:[21.8, 0.0, 48.2] SR:0 DR:9 LR:-21.85 LO:22.41);ALT=C]chr18:66610044];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	194689502	+	chr2	194698766	+	.	48	42	1592912_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1592912_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_194677001_194702001_141C;SPAN=9264;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:42 DR:48 LR:-237.7 LO:237.7);ALT=G[chr2:194698766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	98586533	+	chr2	211048737	+	.	2	14	7154297_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CATTGCACT;MAPQ=60;MATEID=7154297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_98563501_98588501_715C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:14 DP:194 GQ:6.1 PL:[0.0, 6.1, 481.9] SR:14 DR:2 LR:6.345 LO:25.07);ALT=]chr11:98586533]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	228252411	-	chr2	228473779	+	.	18	0	1732621_1	38.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=1732621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:228252411(-)-2:228473779(-)__2_228462501_228487501D;SPAN=221368;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:77 GQ:38.6 PL:[38.6, 0.0, 147.5] SR:0 DR:18 LR:-38.56 LO:42.19);ALT=[chr2:228473779[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	228475751	+	chr15	80435841	+	.	29	26	1732718_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CCTGGCCAAGATGGTGAAACC;MAPQ=60;MATEID=1732718_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_228462501_228487501_367C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:47 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:26 DR:29 LR:-138.6 LO:138.6);ALT=C[chr15:80435841[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	229264346	+	chr2	229268337	+	.	61	76	1735632_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=1735632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_229246501_229271501_301C;SPAN=3991;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:110 DP:96 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:76 DR:61 LR:-326.8 LO:326.8);ALT=A[chr2:229268337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9891163	-	chr19	22762790	+	.	17	0	10221698_1	31.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=10221698_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:9891163(-)-19:22762790(-)__19_22760501_22785501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:93 GQ:31.1 PL:[31.1, 0.0, 192.8] SR:0 DR:17 LR:-30.92 LO:37.78);ALT=[chr19:22762790[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	10096014	+	chr3	10038203	+	.	27	0	1835111_1	75.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1835111_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10038203(-)-3:10096014(+)__3_10020501_10045501D;SPAN=57811;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:49 GQ:42.8 PL:[75.8, 0.0, 42.8] SR:0 DR:27 LR:-76.34 LO:76.34);ALT=]chr3:10096014]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	11108285	+	chr3	11111884	+	.	87	35	1840100_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1840100_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_3_11098501_11123501_215C;SECONDARY;SPAN=3599;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:88 GQ:27 PL:[297.0, 27.0, 0.0] SR:35 DR:87 LR:-297.1 LO:297.1);ALT=T[chr3:11111884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	11645733	+	chr3	11646735	+	TCA	0	47	1842927_1	99.0	.	EVDNC=ASSMB;INSERTION=TCA;MAPQ=60;MATEID=1842927_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_11637501_11662501_225C;SPAN=1002;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:62 GQ:9.8 PL:[138.5, 0.0, 9.8] SR:47 DR:0 LR:-144.6 LO:144.6);ALT=A[chr3:11646735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	11955918	+	chr3	12913421	+	.	38	0	1843939_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1843939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:11955918(+)-3:12913421(-)__3_11931501_11956501D;SPAN=957503;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:38 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:0 DR:38 LR:-112.2 LO:112.2);ALT=T[chr3:12913421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	12715197	-	chr4	147210876	+	GAAAAAAGTGTA	13	54	1848242_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=GAAAAAAGTGTA;MAPQ=60;MATEID=1848242_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_12691001_12716001_491C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:18 GQ:18 PL:[198.0, 18.0, 0.0] SR:54 DR:13 LR:-198.0 LO:198.0);ALT=[chr4:147210876[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	13911208	+	chr3	13910199	+	.	8	0	1853125_1	10.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1853125_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:13910199(-)-3:13911208(+)__3_13891501_13916501D;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=]chr3:13911208]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	6962624	+	chr3	75463422	+	.	10	0	4523781_1	15.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=4523781_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:75463422(-)-7:6962624(+)__7_6958001_6983001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:0 DR:10 LR:-15.67 LO:21.47);ALT=]chr7:6962624]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	9666441	+	chr3	75606396	+	.	12	0	2118077_1	25.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=2118077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:75606396(-)-4:9666441(+)__3_75582501_75607501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=]chr4:9666441]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	3587475	+	chr3	75614077	+	.	10	0	2116751_1	9.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2116751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:75614077(-)-11:3587475(+)__3_75607001_75632001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:0 DR:10 LR:-9.711 LO:20.09);ALT=]chr11:3587475]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	125408095	+	chr3	125404879	+	.	0	51	2298700_1	99.0	.	EVDNC=ASSMB;HOMSEQ=T;MAPQ=60;MATEID=2298700_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_125391001_125416001_363C;SPAN=3216;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:142 GQ:99 PL:[130.1, 0.0, 212.6] SR:51 DR:0 LR:-129.9 LO:131.0);ALT=]chr3:125408095]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	125472587	+	chr3	125450122	+	.	14	0	2299196_1	24.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2299196_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:125450122(-)-3:125472587(+)__3_125440001_125465001D;SPAN=22465;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:80 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:0 DR:14 LR:-24.54 LO:30.82);ALT=]chr3:125472587]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	3454586	+	chr3	125624695	+	.	4	3	6625619_1	1.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=CCATCCTC;MAPQ=60;MATEID=6625619_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_3454501_3479501_276C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:5 DP:56 GQ:1.4 PL:[1.4, 0.0, 133.4] SR:3 DR:4 LR:-1.333 LO:9.437);ALT=]chr11:3454586]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	125672309	+	chr3	125676376	+	.	50	0	2300725_1	99.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=2300725_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:125672309(+)-3:125676376(-)__3_125660501_125685501D;SPAN=4067;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:70 GQ:23.9 PL:[146.0, 0.0, 23.9] SR:0 DR:50 LR:-151.1 LO:151.1);ALT=G[chr3:125676376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	135260733	-	chr6	43257761	+	.	2	34	2340726_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=ATATATATACACACACACACATATATA;MAPQ=20;MATEID=2340726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_135240001_135265001_333C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:34 DP:40 GQ:4.2 PL:[105.6, 4.2, 0.0] SR:34 DR:2 LR:-108.9 LO:108.9);ALT=[chr6:43257761[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	136021013	+	chr3	136026200	+	A	81	61	2343975_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=2343975_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_136024001_136049001_219C;SPAN=5187;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:118 DP:42 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:61 DR:81 LR:-349.9 LO:349.9);ALT=C[chr3:136026200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	144734789	+	chr9	98994270	-	.	10	0	2381710_1	9.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2381710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:144734789(+)-9:98994270(+)__3_144721501_144746501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:0 DR:10 LR:-9.44 LO:20.03);ALT=C]chr9:98994270];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr20	16875043	+	chr3	159596233	+	.	7	18	2441232_1	62.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TGCACTCCAGCCTGGGCGACAGAGTGAGACTCTGTCTCAAAAAATAAAAATA;MAPQ=42;MATEID=2441232_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_159593001_159618001_23C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:73 GQ:62.9 PL:[62.9, 0.0, 112.4] SR:18 DR:7 LR:-62.75 LO:63.57);ALT=]chr20:16875043]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	160438239	+	chr3	160232333	+	.	8	0	2444857_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2444857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:160232333(-)-3:160438239(+)__3_160426001_160451001D;SPAN=205906;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:0 DR:8 LR:-8.527 LO:16.22);ALT=]chr3:160438239]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	166540660	+	chr9	89203834	+	.	8	0	5916622_1	12.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=5916622_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:166540660(+)-9:89203834(-)__9_89180001_89205001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=A[chr9:89203834[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	166840449	+	chr3	166791338	+	TCCT	54	43	2468149_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCCT;MAPQ=60;MATEID=2468149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_166820501_166845501_274C;SPAN=49111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:53 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:43 DR:54 LR:-241.0 LO:241.0);ALT=]chr3:166840449]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	194398724	+	chr3	194400290	+	.	47	0	2583402_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2583402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:194398724(+)-3:194400290(-)__3_194383001_194408001D;SPAN=1566;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:71 GQ:33.8 PL:[136.1, 0.0, 33.8] SR:0 DR:47 LR:-139.1 LO:139.1);ALT=C[chr3:194400290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	194543294	+	chr3	194546257	+	.	63	49	2584510_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=2584510_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_194530001_194555001_357C;SPAN=2963;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:122 GQ:3 PL:[300.3, 3.0, 0.0] SR:49 DR:63 LR:-315.7 LO:315.7);ALT=G[chr3:194546257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	194546431	+	chr3	194543310	+	.	34	56	2584511_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2584511_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_3_194530001_194555001_273C;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:83 DP:116 GQ:38 PL:[242.6, 0.0, 38.0] SR:56 DR:34 LR:-251.0 LO:251.0);ALT=]chr3:194546431]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	195194116	+	chr20	3349267	+	.	9	0	2587616_1	20.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2587616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195194116(+)-20:3349267(-)__3_195191501_195216501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=T[chr20:3349267[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	3582302	+	chr4	3579696	+	.	9	0	2613948_1	7.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=2613948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3579696(-)-4:3582302(+)__4_3577001_3602001D;SPAN=2606;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:0 DR:9 LR:-6.951 LO:17.74);ALT=]chr4:3582302]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	3931722	-	chr4	4005043	+	.	22	0	2615367_1	63.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2615367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3931722(-)-4:4005043(-)__4_3993501_4018501D;SPAN=73321;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:34 GQ:17.3 PL:[63.5, 0.0, 17.3] SR:0 DR:22 LR:-64.73 LO:64.73);ALT=[chr4:4005043[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	4006796	+	chr4	9641379	-	.	15	0	2615400_1	42.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=2615400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:4006796(+)-4:9641379(+)__4_3993501_4018501D;SPAN=5634583;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:14 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=T]chr4:9641379];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	4014946	-	chr4	9633060	+	.	41	0	2629795_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2629795_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:4014946(-)-4:9633060(-)__4_9628501_9653501D;SPAN=5618114;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:7 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=[chr4:9633060[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	4265580	-	chrX	13693567	+	GTTGTGCTGAGCCAAGATCGCACCACTGCACTCCAGCCTGGGCAACCAGAGCGAAACTCTGTC	7	79	10980261_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=GTTGTGCTGAGCCAAGATCGCACCACTGCACTCCAGCCTGGGCAACCAGAGCGAAACTCTGTC;MAPQ=60;MATEID=10980261_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_23_13671001_13696001_34C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:38 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:79 DR:7 LR:-237.7 LO:237.7);ALT=[chrX:13693567[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	9457225	+	chr4	9481542	+	.	41	0	2627932_1	99.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2627932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:9457225(+)-4:9481542(-)__4_9481501_9506501D;SPAN=24317;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:18 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=A[chr4:9481542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	9494936	+	chr4	9492754	+	.	15	36	2627967_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GATGCGGGGAGTAAGAGCCAGCCCCTC;MAPQ=60;MATEID=2627967_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_9481501_9506501_343C;SPAN=2182;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:49 DP:45 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:36 DR:15 LR:-145.2 LO:145.2);ALT=]chr4:9494936]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	10211267	+	chr4	10234568	+	.	81	57	2630662_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTTCAA;MAPQ=60;MATEID=2630662_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_10192001_10217001_152C;SPAN=23301;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:108 DP:9 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:57 DR:81 LR:-320.2 LO:320.2);ALT=A[chr4:10234568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	30377377	+	chr13	49892594	-	.	10	27	8059984_1	34.0	.	DISC_MAPQ=0;EVDNC=TSI_L;HOMSEQ=A;MAPQ=60;MATEID=8059984_2;MATENM=13;NM=0;NUMPARTS=3;REPSEQ=AAAAGAAAAG;SCTG=c_13_49882001_49907001_36C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:30 DP:16 GQ:7.5 PL:[34.5, 7.5, 0.0] SR:27 DR:10 LR:-34.53 LO:34.53);ALT=T]chr13:49892594];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	30474825	+	chr12	71022112	-	.	22	0	7720066_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7720066_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:30474825(+)-12:71022112(+)__12_71001001_71026001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:121 GQ:40.1 PL:[40.1, 0.0, 251.3] SR:0 DR:22 LR:-39.84 LO:48.84);ALT=G]chr12:71022112];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	61663773	+	chr4	36216927	+	.	0	40	3469637_1	99.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=3469637_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_61642001_61667001_78C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:90 GQ:99 PL:[107.6, 0.0, 110.9] SR:40 DR:0 LR:-107.7 LO:107.7);ALT=]chr5:61663773]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	36224538	+	chr5	35606222	-	.	55	39	2681598_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=2681598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_36211001_36236001_20C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:39 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:39 DR:55 LR:-224.5 LO:224.5);ALT=A]chr5:35606222];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	44795699	+	chr5	72498253	-	ATTTTTTA	18	30	3529070_1	94.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=T;INSERTION=ATTTTTTA;MAPQ=60;MATEID=3529070_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTTTT;SCTG=c_5_72495501_72520501_48C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:85 GQ:57.8 PL:[94.2, 0.0, 57.8] SR:30 DR:18 LR:-94.57 LO:94.57);ALT=T]chr5:72498253];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	72498253	+	chr4	44795702	+	GCCCTACTTTTATTAAATATACACCTATTTTATTGTTTTTGATGCTATTGTAAATAGTATTGCTTTATTAATTTTGTCTTTTTTTCTAGTATATAGAAATACAATTGATTTTATTATATTTAACTTATTTTTTA	13	71	3529071_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=T;INSERTION=GCCCTACTTTTATTAAATATACACCTATTTTATTGTTTTTGATGCTATTGTAAATAGTATTGCTTTATTAATTTTGTCTTTTTTTCTAGTATATAGAAATACAATTGATTTTATTATATTTAACTTATTTTTTA;MAPQ=60;MATEID=3529071_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_5_72495501_72520501_48C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:85 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:71 DR:13 LR:-250.9 LO:250.9);ALT=]chr5:72498253]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	45554647	+	chr4	45545415	+	.	8	0	2701840_1	11.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2701840_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:45545415(-)-4:45554647(+)__4_45521001_45546001D;SPAN=9232;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=]chr4:45554647]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	46055996	+	chr4	46058203	+	A	0	43	2703802_1	99.0	.	EVDNC=ASSMB;INSERTION=A;MAPQ=60;MATEID=2703802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_46035501_46060501_180C;SPAN=2207;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:43 DP:139 GQ:99 PL:[104.3, 0.0, 233.0] SR:43 DR:0 LR:-104.3 LO:107.0);ALT=T[chr4:46058203[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	46202797	+	chr4	46205027	+	.	122	104	2703958_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=2703958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_46182501_46207501_188C;SPAN=2230;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:179 DP:37 GQ:48.4 PL:[531.4, 48.4, 0.0] SR:104 DR:122 LR:-531.4 LO:531.4);ALT=C[chr4:46205027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	46740313	+	chr4	46987218	+	.	57	57	2706277_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=2706277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_46966501_46991501_4C;SPAN=246905;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:33 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:57 DR:57 LR:-277.3 LO:277.3);ALT=A[chr4:46987218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	47262254	+	chr4	100270984	+	.	32	0	2800050_1	92.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=2800050_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:47262254(+)-4:100270984(-)__4_100254001_100279001D;SPAN=53008730;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:47 GQ:20.3 PL:[92.9, 0.0, 20.3] SR:0 DR:32 LR:-95.43 LO:95.43);ALT=G[chr4:100270984[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	100224580	+	chr6	79723785	+	.	8	14	2799625_1	45.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=39;MATEID=2799625_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_100205001_100230001_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:28 GQ:22.1 PL:[45.2, 0.0, 22.1] SR:14 DR:8 LR:-45.63 LO:45.63);ALT=A[chr6:79723785[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	100699496	+	chr4	105044838	+	.	88	54	2813168_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=32;MATEID=2813168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_105031501_105056501_402C;SPAN=4345342;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:72 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:54 DR:88 LR:-340.0 LO:340.0);ALT=T[chr4:105044838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	102336327	+	chr20	47019890	+	.	19	40	10587593_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=CTTCCTTCCTTCCTTCCTTCCTTC;MAPQ=60;MATEID=10587593_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_47015501_47040501_36C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:54 DP:43 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:40 DR:19 LR:-158.4 LO:158.4);ALT=G[chr20:47019890[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	106196607	+	chr4	103050633	+	.	91	66	2819630_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2819630_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_106183001_106208001_135C;SPAN=3145974;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:127 DP:89 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:66 DR:91 LR:-376.3 LO:376.3);ALT=]chr4:106196607]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	104140510	+	chr4	104135594	+	.	4	3	2809809_1	0	.	DISC_MAPQ=39;EVDNC=ASDIS;MAPQ=60;MATEID=2809809_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_104125001_104150001_26C;SPAN=4916;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:140 GQ:21.3 PL:[0.0, 21.3, 382.8] SR:3 DR:4 LR:21.42 LO:7.395);ALT=]chr4:104140510]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	106427337	-	chr4	106428472	+	.	9	0	2821312_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2821312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:106427337(-)-4:106428472(-)__4_106403501_106428501D;SPAN=1135;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:131 GQ:5.4 PL:[0.0, 5.4, 326.7] SR:0 DR:9 LR:5.782 LO:15.92);ALT=[chr4:106428472[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	106922710	+	chr4	106538354	+	.	68	59	2823869_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=2823869_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_4_106918001_106943001_332C;SPAN=384356;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:78 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:59 DR:68 LR:-293.8 LO:293.8);ALT=]chr4:106922710]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	107056578	+	chr4	107063363	+	CA	49	41	2824727_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CA;MAPQ=60;MATEID=2824727_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_107040501_107065501_272C;SPAN=6785;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:68 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:41 DR:49 LR:-214.6 LO:214.6);ALT=C[chr4:107063363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107317375	-	chr4	107320346	+	.	28	0	2825811_1	55.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2825811_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107317375(-)-4:107320346(-)__4_107310001_107335001D;SPAN=2971;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:138 GQ:55.1 PL:[55.1, 0.0, 279.5] SR:0 DR:28 LR:-55.04 LO:63.66);ALT=[chr4:107320346[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	107372864	+	chr6	140408919	+	.	61	71	4408438_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4408438_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_140385001_140410001_177C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:97 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:71 DR:61 LR:-310.3 LO:310.3);ALT=C[chr6:140408919[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	107372909	+	chr6	140409425	+	.	63	0	4408742_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4408742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107372909(+)-6:140409425(-)__6_140409501_140434501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:18 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:0 DR:63 LR:-184.8 LO:184.8);ALT=G[chr6:140409425[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	108127828	+	chr4	108131715	+	.	133	72	2827354_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAACATTAGGATTCTCTTT;MAPQ=60;MATEID=2827354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108118501_108143501_80C;SPAN=3887;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:174 DP:34 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:72 DR:133 LR:-514.9 LO:514.9);ALT=T[chr4:108131715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147953942	+	chr20	54914679	-	.	33	38	10639455_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=10639455_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_54904501_54929501_480C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:100 GQ:65.3 PL:[177.5, 0.0, 65.3] SR:38 DR:33 LR:-180.4 LO:180.4);ALT=C]chr20:54914679];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	147953944	-	chr20	54914484	+	.	49	47	10639456_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=10639456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_54904501_54929501_79C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:76 DP:105 GQ:31.1 PL:[222.5, 0.0, 31.1] SR:47 DR:49 LR:-230.6 LO:230.6);ALT=[chr20:54914484[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	10547399	+	chr4	165897428	+	.	8	0	7390174_1	0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=7390174_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:165897428(-)-12:10547399(+)__12_10535001_10560001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:102 GQ:0.9 PL:[0.0, 0.9, 247.5] SR:0 DR:8 LR:1.226 LO:14.63);ALT=]chr12:10547399]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	166002672	+	chr4	166005035	+	.	95	0	3046301_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3046301_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:166002672(+)-4:166005035(-)__4_165987501_166012501D;SPAN=2363;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:12 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:0 DR:95 LR:-280.6 LO:280.6);ALT=A[chr4:166005035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	3657092	+	chr5	3660542	+	.	166	94	3162421_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GACC;MAPQ=60;MATEID=3162421_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_3650501_3675501_61C;SPAN=3450;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:217 DP:97 GQ:58.6 PL:[643.6, 58.6, 0.0] SR:94 DR:166 LR:-643.7 LO:643.7);ALT=C[chr5:3660542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	3694118	+	chrX	11731470	-	.	9	0	10972464_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=10972464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:3694118(+)-23:11731470(+)__23_11711001_11736001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:0 DR:9 LR:-14.0 LO:19.3);ALT=G]chrX:11731470];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr20	22863420	+	chr5	9024438	+	.	10	0	3194398_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=3194398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:9024438(-)-20:22863420(+)__5_9016001_9041001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:121 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.2281 LO:18.52);ALT=]chr20:22863420]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	56485981	-	chr12	6643683	+	.	20	55	7360560_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7360560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6639501_6664501_524C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:73 GQ:3.5 PL:[171.8, 0.0, 3.5] SR:55 DR:20 LR:-181.1 LO:181.1);ALT=[chr12:6643683[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	57323478	+	chr5	57333779	+	.	183	74	3449613_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=3449613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_57330001_57355001_369C;SPAN=10301;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:230 DP:32 GQ:62.2 PL:[683.2, 62.2, 0.0] SR:74 DR:183 LR:-683.3 LO:683.3);ALT=C[chr5:57333779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57680001	+	chr5	57686102	+	.	151	111	3451593_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAACAC;MAPQ=60;MATEID=3451593_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_57673001_57698001_157C;SPAN=6101;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:241 DP:63 GQ:64.9 PL:[712.9, 64.9, 0.0] SR:111 DR:151 LR:-713.0 LO:713.0);ALT=C[chr5:57686102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	58412650	+	chr5	62573925	-	.	12	65	3456997_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=3456997_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_5_58408001_58433001_468C;SPAN=4161275;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:99 GQ:19.4 PL:[220.7, 0.0, 19.4] SR:65 DR:12 LR:-230.7 LO:230.7);ALT=A]chr5:62573925];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	58412680	+	chr5	62911008	-	.	10	0	3477421_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3477421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:58412680(+)-5:62911008(+)__5_62891501_62916501D;SPAN=4498328;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:81 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.07 LO:20.36);ALT=A]chr5:62911008];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	58988176	-	chr7	80802060	+	.	19	0	5000967_1	46.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5000967_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:58988176(-)-7:80802060(-)__7_80801001_80826001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:61 GQ:46.4 PL:[46.4, 0.0, 99.2] SR:0 DR:19 LR:-46.19 LO:47.34);ALT=[chr7:80802060[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	58988321	+	chr7	80801568	-	.	16	0	5000972_1	34.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=5000972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:58988321(+)-7:80801568(+)__7_80801001_80826001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:69 GQ:34.1 PL:[34.1, 0.0, 133.1] SR:0 DR:16 LR:-34.12 LO:37.43);ALT=A]chr7:80801568];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	59623345	+	chr5	59624805	-	.	9	0	3461361_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3461361_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:59623345(+)-5:59624805(+)__5_59608501_59633501D;SPAN=1460;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:129 GQ:5.1 PL:[0.0, 5.1, 323.4] SR:0 DR:9 LR:5.24 LO:15.98);ALT=A]chr5:59624805];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	60001709	+	chr5	60003666	+	.	81	54	3462761_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACTAA;MAPQ=60;MATEID=3462761_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_60000501_60025501_59C;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:79 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:54 DR:81 LR:-326.8 LO:326.8);ALT=A[chr5:60003666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	62573338	+	chr5	62910687	+	.	26	0	3475820_1	63.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=3475820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:62573338(+)-5:62910687(-)__5_62573001_62598001D;SPAN=337349;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:84 GQ:63.2 PL:[63.2, 0.0, 139.1] SR:0 DR:26 LR:-63.07 LO:64.7);ALT=C[chr5:62910687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43751247	+	chr5	63370313	+	.	3	19	3478773_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATATA;MAPQ=60;MATEID=3478773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_63357001_63382001_247C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:19 DP:14 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:19 DR:3 LR:-56.11 LO:56.11);ALT=]chr22:43751247]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	63965726	-	chr7	131553229	+	.	13	21	3481134_1	87.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GATAGATAGATAGATAGATAGA;MAPQ=60;MATEID=3481134_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_63945001_63970001_377C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:80 GQ:87.2 PL:[87.2, 0.0, 107.0] SR:21 DR:13 LR:-87.26 LO:87.37);ALT=[chr7:131553229[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	71121296	+	chr5	73276601	-	.	74	30	3523120_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=3523120_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_71099001_71124001_175C;SPAN=2155305;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:93 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:30 DR:74 LR:-277.3 LO:277.3);ALT=T]chr5:73276601];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	72348054	+	chr5	72349093	-	.	8	0	3527830_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3527830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:72348054(+)-5:72349093(+)__5_72324001_72349001D;SPAN=1039;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:159 GQ:16.6 PL:[0.0, 16.6, 419.2] SR:0 DR:8 LR:16.67 LO:13.04);ALT=G]chr5:72349093];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	72743130	+	chr5	72977752	+	.	14	21	3532084_1	70.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3532084_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_72961001_72986001_10C;SPAN=234622;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:70 GQ:70.1 PL:[70.1, 0.0, 99.8] SR:21 DR:14 LR:-70.16 LO:70.45);ALT=C[chr5:72977752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134119173	+	chr9	133575625	+	.	25	0	3773047_1	74.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3773047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:134119173(+)-9:133575625(-)__5_134113001_134138001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:32 GQ:1.4 PL:[74.0, 0.0, 1.4] SR:0 DR:25 LR:-77.64 LO:77.64);ALT=T[chr9:133575625[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	146394711	+	chr5	146397308	+	TTAGG	0	49	3826228_1	99.0	.	EVDNC=ASSMB;INSERTION=TTAGG;MAPQ=60;MATEID=3826228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_146387501_146412501_379C;SPAN=2597;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:81 GQ:54.2 PL:[140.0, 0.0, 54.2] SR:49 DR:0 LR:-141.7 LO:141.7);ALT=A[chr5:146397308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	146663607	-	chrX	74928699	+	.	3	79	11248408_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TCCAACAGC;MAPQ=60;MATEID=11248408_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_74921001_74946001_393C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:40 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:79 DR:3 LR:-237.7 LO:237.7);ALT=[chrX:74928699[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	147553129	+	chr5	147554643	-	.	65	0	3830699_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3830699_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:147553129(+)-5:147554643(+)__5_147539001_147564001D;SPAN=1514;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:73 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:0 DR:65 LR:-212.9 LO:212.9);ALT=T]chr5:147554643];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	168238968	-	chr11	92072561	+	.	58	55	7082905_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AACA;MAPQ=60;MATEID=7082905_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_92071001_92096001_687C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:91 DP:218 GQ:99 PL:[241.4, 0.0, 287.6] SR:55 DR:58 LR:-241.3 LO:241.6);ALT=[chr11:92072561[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	73565519	+	chr6	42820282	+	.	0	15	8597434_1	25.0	.	EVDNC=ASSMB;HOMSEQ=CCCAGCTACT;MAPQ=60;MATEID=8597434_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73549001_73574001_102C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:88 GQ:25.7 PL:[25.7, 0.0, 187.4] SR:15 DR:0 LR:-25.67 LO:32.83);ALT=]chr14:73565519]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	43532491	-	chr6	43533988	+	.	5	3	4172278_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGGTGTGGTGG;MAPQ=60;MATEID=4172278_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_43512001_43537001_150C;SPAN=1497;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:147 GQ:19.9 PL:[0.0, 19.9, 396.0] SR:3 DR:5 LR:20.02 LO:9.226);ALT=[chr6:43533988[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	43655533	+	chr9	33130549	+	CGTAATTTTTTC	7	32	5815542_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CGTAATTTTTTC;MAPQ=60;MATEID=5815542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33124001_33149001_167C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:37 DP:23 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:32 DR:7 LR:-108.9 LO:108.9);ALT=T[chr9:33130549[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	65336579	+	chr15	56253097	+	.	25	58	8905883_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=8905883_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_56252001_56277001_173C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:56 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:58 DR:25 LR:-184.8 LO:184.8);ALT=T[chr15:56253097[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	66260039	+	chr6	66262022	+	.	135	120	4253415_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TACTATATCTTT;MAPQ=60;MATEID=4253415_2;MATENM=2;NM=6;NUMPARTS=2;SCTG=c_6_66248001_66273001_163C;SPAN=1983;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:204 DP:57 GQ:55 PL:[604.0, 55.0, 0.0] SR:120 DR:135 LR:-604.0 LO:604.0);ALT=T[chr6:66262022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	67040800	+	chr6	67043190	+	AATTAATACATGCCAGATT	0	156	4256179_1	99.0	.	EVDNC=ASSMB;INSERTION=AATTAATACATGCCAGATT;MAPQ=60;MATEID=4256179_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_67032001_67057001_338C;SPAN=2390;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:156 DP:58 GQ:42.1 PL:[462.1, 42.1, 0.0] SR:156 DR:0 LR:-462.1 LO:462.1);ALT=T[chr6:67043190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	69242155	+	chr6	67771676	+	.	42	19	4260669_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=4260669_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_6_67767001_67792001_154C;SPAN=1470479;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:64 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:19 DR:42 LR:-194.7 LO:194.7);ALT=]chr6:69242155]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	67771990	+	chr6	69242387	+	.	11	0	4260677_1	16.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=4260677_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:67771990(+)-6:69242387(-)__6_67767001_67792001D;SPAN=1470397;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:0 DR:11 LR:-15.99 LO:23.29);ALT=C[chr6:69242387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	68101533	+	chr6	68112167	+	.	102	48	4260126_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4260126_2;MATENM=1;NM=3;NUMPARTS=2;SCTG=c_6_68085501_68110501_77C;SPAN=10634;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:142 DP:88 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:48 DR:102 LR:-419.2 LO:419.2);ALT=T[chr6:68112167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	68144663	-	chr6	140607373	+	.	44	28	4410160_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=4410160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_140605501_140630501_527C;SPAN=72462710;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:92 GQ:64.4 PL:[156.8, 0.0, 64.4] SR:28 DR:44 LR:-158.6 LO:158.6);ALT=[chr6:140607373[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	68148896	+	chr6	140538018	-	.	51	33	4409525_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=4409525_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_140532001_140557001_131C;SPAN=72389122;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:99 GQ:19.4 PL:[220.7, 0.0, 19.4] SR:33 DR:51 LR:-230.7 LO:230.7);ALT=A]chr6:140538018];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	68433574	+	chr6	76642373	+	.	52	69	4285239_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=4285239_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_76636001_76661001_356C;SPAN=8208799;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:88 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:69 DR:52 LR:-287.2 LO:287.2);ALT=T[chr6:76642373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	74014515	-	chr6	74015639	+	.	8	0	4272168_1	10.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4272168_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:74014515(-)-6:74015639(-)__6_73990001_74015001D;SPAN=1124;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=[chr6:74015639[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	74476277	+	chr6	133948854	-	.	3	42	4395469_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATATA;MAPQ=60;MATEID=4395469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_133941501_133966501_306C;SPAN=59472577;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:44 DP:20 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:42 DR:3 LR:-128.7 LO:128.7);ALT=T]chr6:133948854];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	74512036	-	chr17	8082371	+	.	2	14	4275214_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTT;MAPQ=60;MATEID=4275214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_74504501_74529501_287C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:36 GQ:43.1 PL:[43.1, 0.0, 43.1] SR:14 DR:2 LR:-43.06 LO:43.06);ALT=[chr17:8082371[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	74592062	+	chr6	74602440	+	.	136	31	4275875_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=4275875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_74602501_74627501_100C;SPAN=10378;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:151 DP:12 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:31 DR:136 LR:-445.6 LO:445.6);ALT=T[chr6:74602440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	74865448	+	chr6	74866585	+	.	119	91	4276847_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAACCAAGTTATT;MAPQ=60;MATEID=4276847_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_6_74847501_74872501_367C;SPAN=1137;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:170 DP:41 GQ:46 PL:[505.0, 46.0, 0.0] SR:91 DR:119 LR:-505.0 LO:505.0);ALT=T[chr6:74866585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	78885753	+	chr6	75799689	+	.	69	56	4298777_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4298777_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_78865501_78890501_154C;SPAN=3086064;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:50 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:56 DR:69 LR:-293.8 LO:293.8);ALT=]chr6:78885753]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	142813858	+	chr6	76428930	+	.	52	21	4422891_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=4422891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_142810501_142835501_28C;SPAN=66384928;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:21 DR:52 LR:-208.0 LO:208.0);ALT=]chr6:142813858]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	141800830	+	chr6	76943995	+	.	44	28	4416765_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4416765_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_141781501_141806501_156C;SPAN=64856835;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:141 GQ:99 PL:[153.5, 0.0, 186.5] SR:28 DR:44 LR:-153.3 LO:153.5);ALT=]chr6:141800830]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	77097496	+	chr6	77102642	+	.	150	64	4288874_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTAT;MAPQ=60;MATEID=4288874_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_6_77101501_77126501_87C;SPAN=5146;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:173 DP:27 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:64 DR:150 LR:-511.6 LO:511.6);ALT=T[chr6:77102642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	81297103	+	chr6	77471429	+	.	0	10	4290846_1	0	.	EVDNC=ASSMB;HOMSEQ=CCCAAATCTCAT;MAPQ=60;MATEID=4290846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_77469001_77494001_267C;SPAN=3825674;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:137 GQ:3.9 PL:[0.0, 3.9, 339.9] SR:10 DR:0 LR:4.107 LO:17.96);ALT=]chr6:81297103]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	78846688	+	chr14	44886697	+	TTCCTGGTCAGTAAGACCTCAAAAGG	17	52	8473833_1	99.0	.	DISC_MAPQ=10;EVDNC=TSI_L;HOMSEQ=TATCTCTAGA;INSERTION=TTCCTGGTCAGTAAGACCTCAAAAGG;MAPQ=38;MATEID=8473833_2;MATENM=0;NM=14;NUMPARTS=5;SCTG=c_14_44884001_44909001_156C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:50 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:52 DR:17 LR:-178.2 LO:178.2);ALT=A[chr14:44886697[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	79448918	+	chr6	79451419	-	.	8	0	4300104_1	10.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=4300104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:79448918(+)-6:79451419(+)__6_79429001_79454001D;SPAN=2501;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=C]chr6:79451419];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	81625982	+	chr6	81630664	+	.	63	37	4304362_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGGACAGAGAGATT;MAPQ=60;MATEID=4304362_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_6_81609501_81634501_268C;SPAN=4682;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:16 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:37 DR:63 LR:-241.0 LO:241.0);ALT=T[chr6:81630664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	133341834	+	chr6	133347886	+	.	69	30	4394569_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTGTGATGTTTT;MAPQ=60;MATEID=4394569_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_133329001_133354001_198C;SPAN=6052;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:59 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:30 DR:69 LR:-260.8 LO:260.8);ALT=T[chr6:133347886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	140176538	-	chr6	140178139	+	.	45	40	4407384_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTG;MAPQ=60;MATEID=4407384_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_140164501_140189501_358C;SPAN=1601;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:76 DP:104 GQ:28.1 PL:[222.8, 0.0, 28.1] SR:40 DR:45 LR:-231.2 LO:231.2);ALT=[chr6:140178139[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	140662555	+	chr6	141794002	+	.	89	31	4410445_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4410445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_140654501_140679501_106C;SPAN=1131447;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:126 GQ:14.1 PL:[333.3, 14.1, 0.0] SR:31 DR:89 LR:-342.5 LO:342.5);ALT=A[chr6:141794002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	142075377	-	chr6	142076383	+	.	10	0	4419208_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4419208_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:142075377(-)-6:142076383(-)__6_142051001_142076001D;SPAN=1006;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=[chr6:142076383[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	142411706	+	chr12	71020308	+	.	10	22	7720078_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGAA;MAPQ=60;MATEID=7720078_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_71001001_71026001_341C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:152 GQ:38.3 PL:[38.3, 0.0, 328.7] SR:22 DR:10 LR:-38.04 LO:51.65);ALT=A[chr12:71020308[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	143114796	+	chr8	125929193	+	.	6	31	4424638_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTCTTTCTTTCTTTCTTTCTTTCTTT;MAPQ=60;MATEID=4424638_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_143104501_143129501_378C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:51 GQ:29.3 PL:[92.0, 0.0, 29.3] SR:31 DR:6 LR:-93.4 LO:93.4);ALT=T[chr8:125929193[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	147138126	+	chr6	147131196	+	.	10	0	4440148_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4440148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:147131196(-)-6:147138126(+)__6_147122501_147147501D;SPAN=6930;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:133 GQ:2.7 PL:[0.0, 2.7, 326.7] SR:0 DR:10 LR:3.023 LO:18.09);ALT=]chr6:147138126]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	147133757	+	chr6	147140449	+	.	16	0	4440159_1	35.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4440159_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:147133757(+)-6:147140449(-)__6_147122501_147147501D;SPAN=6692;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:66 GQ:35 PL:[35.0, 0.0, 124.1] SR:0 DR:16 LR:-34.94 LO:37.79);ALT=G[chr6:147140449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	147961979	+	chr6	148086792	+	CATGTTT	88	24	4443314_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CATGTTT;MAPQ=60;MATEID=4443314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_148078001_148103001_198C;SPAN=124813;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:51 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:24 DR:88 LR:-287.2 LO:287.2);ALT=G[chr6:148086792[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93957164	+	chr6	148199082	+	TAGAAAGAAAGATAGATTTTTTTTTCTTTTTGAGACAGAGTCT	16	124	4443981_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TAGAAAGAAAGATAGATTTTTTTTTCTTTTTGAGACAGAGTCT;MAPQ=60;MATEID=4443981_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_148176001_148201001_365C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:129 DP:32 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:124 DR:16 LR:-382.9 LO:382.9);ALT=]chr11:93957164]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	148268010	+	chr7	66272198	-	.	58	49	4912504_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4912504_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_66248001_66273001_36C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:90 DP:162 GQ:99 PL:[253.4, 0.0, 137.9] SR:49 DR:58 LR:-255.0 LO:255.0);ALT=T]chr7:66272198];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	150101299	+	chr19	39037385	+	.	11	27	10288295_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=AGTTTGAGACCAGCCTGGGCAACATGGTGAGA;MAPQ=47;MATEID=10288295_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_19_39028501_39053501_691C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:46 GQ:7.4 PL:[103.1, 0.0, 7.4] SR:27 DR:11 LR:-107.8 LO:107.8);ALT=A[chr19:39037385[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	150353648	+	chr7	7062371	+	TTGTATTTTTAGTAGATGC	12	78	4522830_1	99.0	.	DISC_MAPQ=3;EVDNC=TSI_G;HOMSEQ=GGGGTTTC;INSERTION=TTGTATTTTTAGTAGATGC;MAPQ=34;MATEID=4522830_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_7_7056001_7081001_168C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:19 GQ:21 PL:[231.0, 21.0, 0.0] SR:78 DR:12 LR:-231.1 LO:231.1);ALT=T[chr7:7062371[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	151510041	-	chr6	151511737	+	.	9	0	4451031_1	12.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4451031_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:151510041(-)-6:151511737(-)__6_151508001_151533001D;SPAN=1696;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=[chr6:151511737[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	151776937	-	chr10	43833073	+	.	13	0	6221363_1	25.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=6221363_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:151776937(-)-10:43833073(-)__10_43830501_43855501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:65 GQ:25.4 PL:[25.4, 0.0, 131.0] SR:0 DR:13 LR:-25.3 LO:29.46);ALT=[chr10:43833073[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	151777087	+	chr10	43832692	-	.	8	0	6221364_1	10.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6221364_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:151777087(+)-10:43832692(+)__10_43830501_43855501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:0 DR:8 LR:-10.69 LO:16.71);ALT=G]chr10:43832692];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	152389994	+	chr6	152392234	+	.	74	62	4452855_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACTGC;MAPQ=60;MATEID=4452855_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_152390001_152415001_196C;SPAN=2240;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:14 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:62 DR:74 LR:-326.8 LO:326.8);ALT=C[chr6:152392234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	153029990	+	chr6	153033790	+	.	53	30	4454008_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCTGAAAGAGTATTTATTT;MAPQ=60;MATEID=4454008_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_153027001_153052001_139C;SPAN=3800;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:30 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:30 DR:53 LR:-208.0 LO:208.0);ALT=T[chr6:153033790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	153958371	+	chr6	153961525	+	.	76	46	4455577_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=ATTT;MAPQ=60;MATEID=4455577_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_153958001_153983001_118C;SPAN=3154;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:18 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:46 DR:76 LR:-293.8 LO:293.8);ALT=T[chr6:153961525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	4610803	-	chr10	77452045	+	.	13	40	4509038_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4509038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_4606001_4631001_349C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:51 DP:39 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:40 DR:13 LR:-148.5 LO:148.5);ALT=[chr10:77452045[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	5621462	+	chr7	5625751	+	.	56	0	4514581_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4514581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:5621462(+)-7:5625751(-)__7_5610501_5635501D;SPAN=4289;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:83 GQ:37.1 PL:[162.5, 0.0, 37.1] SR:0 DR:56 LR:-166.6 LO:166.6);ALT=A[chr7:5625751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	5831459	+	chr19	8538236	+	.	33	40	4516380_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TCGGGAGGCTGAGGCAG;MAPQ=60;MATEID=4516380_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_5831001_5856001_508C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:58 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:40 DR:33 LR:-208.0 LO:208.0);ALT=G[chr19:8538236[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	6140427	+	chr7	6141515	-	.	8	0	4517875_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4517875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:6140427(+)-7:6141515(+)__7_6125001_6150001D;SPAN=1088;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:141 GQ:11.4 PL:[0.0, 11.4, 363.0] SR:0 DR:8 LR:11.79 LO:13.47);ALT=A]chr7:6141515];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	6616912	+	chr9	132621563	-	.	9	34	4520679_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=TTTTATTTTATTTTATTTTATTTTATTTTA;MAPQ=10;MATEID=4520679_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_6615001_6640001_336C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:37 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:34 DR:9 LR:-115.5 LO:115.5);ALT=A]chr9:132621563];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	7583516	+	chr7	10708427	-	.	11	73	4538611_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4538611_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_10706501_10731501_295C;SPAN=3124911;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:74 DP:122 GQ:82.7 PL:[211.4, 0.0, 82.7] SR:73 DR:11 LR:-214.2 LO:214.2);ALT=G]chr7:10708427];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	7595533	+	chr7	9818114	+	.	0	51	4533320_1	99.0	.	EVDNC=ASSMB;HOMSEQ=T;MAPQ=60;MATEID=4533320_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_9800001_9825001_290C;SPAN=2222581;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:84 GQ:56.6 PL:[145.7, 0.0, 56.6] SR:51 DR:0 LR:-147.6 LO:147.6);ALT=T[chr7:9818114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	8374193	-	chr8	49965549	+	.	57	54	4527637_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4527637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_8354501_8379501_149C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:49 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:54 DR:57 LR:-274.0 LO:274.0);ALT=[chr8:49965549[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	10312466	+	chr7	10849105	-	.	47	0	4539666_1	99.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=4539666_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:10312466(+)-7:10849105(+)__7_10829001_10854001D;SPAN=536639;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:130 GQ:99 PL:[119.9, 0.0, 195.8] SR:0 DR:47 LR:-119.9 LO:120.9);ALT=C]chr7:10849105];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	10313274	-	chr7	10848217	+	.	19	0	4539667_1	21.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=4539667_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:10313274(-)-7:10848217(-)__7_10829001_10854001D;SPAN=534943;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:152 GQ:21.8 PL:[21.8, 0.0, 345.2] SR:0 DR:19 LR:-21.54 LO:38.8);ALT=[chr7:10848217[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	16171773	+	chr7	16174073	+	.	210	111	4571066_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4571066_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_16170001_16195001_263C;SPAN=2300;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:278 DP:64 GQ:75.2 PL:[825.2, 75.2, 0.0] SR:111 DR:210 LR:-825.2 LO:825.2);ALT=C[chr7:16174073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139205879	+	chr7	16830728	+	.	8	0	5301619_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5301619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:16830728(-)-7:139205879(+)__7_139184501_139209501D;SPAN=122375151;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=]chr7:139205879]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	17094701	-	chrX	11953198	+	.	52	40	10972950_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=10972950_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_11931501_11956501_228C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:64 GQ:21 PL:[231.0, 21.0, 0.0] SR:40 DR:52 LR:-231.1 LO:231.1);ALT=[chrX:11953198[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	17472367	+	chr7	17415035	+	.	80	31	4578713_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=4578713_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_17468501_17493501_417C;SPAN=57332;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:96 DP:128 GQ:28.1 PL:[282.2, 0.0, 28.1] SR:31 DR:80 LR:-294.3 LO:294.3);ALT=]chr7:17472367]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	17753132	+	chr15	89459015	+	.	5	18	4581233_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GTGTGTATATATATA;MAPQ=28;MATEID=4581233_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=ATATATATAT;SCTG=c_7_17738001_17763001_512C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:36 GQ:3.8 PL:[19.2, 0.0, 3.8] SR:18 DR:5 LR:-19.54 LO:19.54);ALT=A[chr15:89459015[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	32390165	+	chr7	32393113	+	.	130	85	4677626_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTGACTAATATAT;MAPQ=60;MATEID=4677626_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_7_32389001_32414001_374C;SPAN=2948;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:193 DP:55 GQ:52 PL:[571.0, 52.0, 0.0] SR:85 DR:130 LR:-571.0 LO:571.0);ALT=T[chr7:32393113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32974630	-	chr16	7059001	+	.	8	0	4682288_1	5.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=4682288_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:32974630(-)-16:7059001(-)__7_32952501_32977501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:0 DR:8 LR:-5.276 LO:15.61);ALT=[chr16:7059001[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	33177805	+	chr7	33179369	+	AATCTACCAGAAGCTTAACAGGGGCATTCAC	0	79	4684129_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TGAGA;INSERTION=AATCTACCAGAAGCTTAACAGGGGCATTCAC;MAPQ=60;MATEID=4684129_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_33173001_33198001_190C;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:79 DP:178 GQ:99 PL:[212.6, 0.0, 219.2] SR:79 DR:0 LR:-212.6 LO:212.6);ALT=G[chr7:33179369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	33848463	+	chr7	33849610	-	.	8	0	4688427_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4688427_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:33848463(+)-7:33849610(+)__7_33834501_33859501D;SPAN=1147;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:183 GQ:22.9 PL:[0.0, 22.9, 488.5] SR:0 DR:8 LR:23.17 LO:12.54);ALT=G]chr7:33849610];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	4619474	+	chr7	54416133	+	.	15	45	4822148_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTATCTATCTATCTATCTATCT;MAPQ=60;MATEID=4822148_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_7_54414501_54439501_209C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:105 GQ:99 PL:[140.0, 0.0, 113.6] SR:45 DR:15 LR:-140.0 LO:140.0);ALT=]chr8:4619474]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	55286758	+	chr7	55289062	+	.	181	104	4827416_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGCAATGTGCTTTTA;MAPQ=60;MATEID=4827416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_55272001_55297001_43C;SPAN=2304;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:244 DP:66 GQ:65.8 PL:[722.8, 65.8, 0.0] SR:104 DR:181 LR:-722.9 LO:722.9);ALT=A[chr7:55289062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	55858685	-	chr7	62570353	+	.	0	35	4833944_1	79.0	.	EVDNC=ASSMB;HOMSEQ=AGAGACATCTAAAAACAA;MAPQ=60;MATEID=4833944_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_55835501_55860501_874C;SPAN=6711668;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:134 GQ:79.4 PL:[79.4, 0.0, 244.4] SR:35 DR:0 LR:-79.23 LO:84.0);ALT=[chr7:62570353[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	63259415	+	chr7	56846631	+	.	4	5	4873307_1	2.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GTACAGG;MAPQ=60;MATEID=4873307_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_63259001_63284001_300C;SPAN=6412784;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:5 DR:4 LR:-1.804 LO:16.9);ALT=]chr7:63259415]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	63029437	+	chr7	57075502	+	.	19	13	4870255_1	75.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CCTTG;MAPQ=57;MATEID=4870255_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_63014001_63039001_442C;SPAN=5953935;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:112 GQ:75.5 PL:[75.5, 0.0, 194.3] SR:13 DR:19 LR:-75.29 LO:78.28);ALT=]chr7:63029437]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	57551927	+	chr7	57556092	+	CAAATCAAATGGAATGGAATGGAATCGAATCAAATGGAATGGAATGGAATTGAATGGGAGCTGAGATTGTGCCACTGCGCTTCAGTCTGGGTGACAGGGTGAGATACTCTAGAAAGAAAGGAATGGAATGGAATGCAGTGG	30	54	4850972_1	99.0	.	DISC_MAPQ=38;EVDNC=TSI_G;HOMSEQ=AATGGAATGGAGTGGACGAGTGGAGTGGAGTGAAGTGGA;INSERTION=CAAATCAAATGGAATGGAATGGAATCGAATCAAATGGAATGGAATGGAATTGAATGGGAGCTGAGATTGTGCCACTGCGCTTCAGTCTGGGTGACAGGGTGAGATACTCTAGAAAGAAAGGAATGGAATGGAATGCAGTGG;MAPQ=0;MATEID=4850972_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_57550501_57575501_193C;SPAN=4165;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:81 DP:324 GQ:99 PL:[179.8, 0.0, 605.6] SR:54 DR:30 LR:-179.6 LO:192.6);ALT=T[chr7:57556092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	57965809	+	chr7	57975176	+	.	48	39	4854308_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TAGTTTTTATGTGAAGATATT;MAPQ=60;MATEID=4854308_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_57942501_57967501_446C;SPAN=9367;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:13 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:39 DR:48 LR:-247.6 LO:247.6);ALT=T[chr7:57975176[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	61847521	+	chr7	61862657	+	.	42	52	4859830_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=CCAAATGTCCATTCACAGAATGGACAAAAACAGT;MAPQ=42;MATEID=4859830_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_7_61838001_61863001_143C;SPAN=15136;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:82 DP:295 GQ:99 PL:[190.9, 0.0, 524.3] SR:52 DR:42 LR:-190.8 LO:199.4);ALT=T[chr7:61862657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	61848994	+	chr7	61857683	+	CAAATATACA	29	18	4859856_1	81.0	.	DISC_MAPQ=10;EVDNC=ASDIS;INSERTION=CAAATATACA;MAPQ=55;MATEID=4859856_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_61838001_61863001_182C;SPAN=8689;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:43 DP:225 GQ:81.1 PL:[81.1, 0.0, 464.0] SR:18 DR:29 LR:-80.99 LO:96.5);ALT=C[chr7:61857683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	62232307	-	chr7	62237451	+	.	8	0	4862978_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4862978_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:62232307(-)-7:62237451(-)__7_62230001_62255001D;SPAN=5144;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:175 GQ:20.8 PL:[0.0, 20.8, 465.4] SR:0 DR:8 LR:21.0 LO:12.7);ALT=[chr7:62237451[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	67427921	+	chr7	63296509	+	.	87	63	4926391_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=4926391_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_67424001_67449001_280C;SPAN=4131412;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:146 DP:75 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:63 DR:87 LR:-432.4 LO:432.4);ALT=]chr7:67427921]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	63711832	-	chr7	63712854	+	.	8	0	4877757_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4877757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:63711832(-)-7:63712854(-)__7_63700001_63725001D;SPAN=1022;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:175 GQ:20.8 PL:[0.0, 20.8, 465.4] SR:0 DR:8 LR:21.0 LO:12.7);ALT=[chr7:63712854[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	64289989	+	chr19	21129556	+	.	40	0	4882360_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4882360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:64289989(+)-19:21129556(-)__7_64288001_64313001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:102 GQ:99 PL:[104.6, 0.0, 140.9] SR:0 DR:40 LR:-104.4 LO:104.7);ALT=T[chr19:21129556[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	64315824	+	chr7	64318059	+	.	182	64	4881333_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGAATTTTATTTTATC;MAPQ=60;MATEID=4881333_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_64312501_64337501_54C;SPAN=2235;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:219 DP:51 GQ:59.2 PL:[650.2, 59.2, 0.0] SR:64 DR:182 LR:-650.3 LO:650.3);ALT=C[chr7:64318059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64556095	-	chr7	65250670	+	.	6	5	4887285_1	0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=TGAGGTCAGGAGTTTGAGACCAGCCTGGCCAACATGGT;MAPQ=22;MATEID=4887285_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_64533001_64558001_354C;SPAN=694575;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:172 GQ:10 PL:[0.0, 10.0, 435.7] SR:5 DR:6 LR:10.29 LO:19.1);ALT=[chr7:65250670[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	64883443	-	chr12	43291992	+	.	54	0	7569284_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=7569284_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:64883443(-)-12:43291992(-)__12_43267001_43292001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:54 DP:85 GQ:49.7 PL:[155.3, 0.0, 49.7] SR:0 DR:54 LR:-158.1 LO:158.1);ALT=[chr12:43291992[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	65238287	+	chr7	65229716	+	.	34	50	4895101_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;MAPQ=23;MATEID=4895101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65219001_65244001_719C;SPAN=8571;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:69 DP:424 GQ:99 PL:[113.1, 0.0, 915.2] SR:50 DR:34 LR:-112.9 LO:149.5);ALT=]chr7:65238287]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	65575674	-	chr7	65579337	+	.	8	0	4901214_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4901214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:65575674(-)-7:65579337(-)__7_65562001_65587001D;SPAN=3663;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:290 GQ:52.1 PL:[0.0, 52.1, 808.6] SR:0 DR:8 LR:52.16 LO:10.93);ALT=[chr7:65579337[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	65857660	+	chr7	65860104	+	.	25	0	4904598_1	20.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4904598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:65857660(+)-7:65860104(-)__7_65856001_65881001D;SPAN=2444;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:229 GQ:20.5 PL:[20.5, 0.0, 535.4] SR:0 DR:25 LR:-20.48 LO:49.49);ALT=T[chr7:65860104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73382119	+	chr7	66193573	+	.	36	68	4960336_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTCCAC;MAPQ=60;MATEID=4960336_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_73377501_73402501_267C;SPAN=7188546;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:67 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:68 DR:36 LR:-293.8 LO:293.8);ALT=]chr7:73382119]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	66633036	+	chr7	72109262	-	.	31	0	4916132_1	65.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=4916132_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:66633036(+)-7:72109262(+)__7_66615501_66640501D;SPAN=5476226;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:137 GQ:65.3 PL:[65.3, 0.0, 266.6] SR:0 DR:31 LR:-65.21 LO:72.15);ALT=T]chr7:72109262];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	66697505	+	chr7	66699292	+	.	119	91	4917056_1	99.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTGGG;MAPQ=60;MATEID=4917056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_66689001_66714001_526C;SPAN=1787;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:196 DP:122 GQ:52.9 PL:[580.9, 52.9, 0.0] SR:91 DR:119 LR:-580.9 LO:580.9);ALT=G[chr7:66699292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66767222	-	chr7	66769167	+	.	9	0	4919060_1	0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=4919060_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:66767222(-)-7:66769167(-)__7_66762501_66787501D;SPAN=1945;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:246 GQ:36.7 PL:[0.0, 36.7, 670.0] SR:0 DR:9 LR:36.94 LO:13.41);ALT=[chr7:66769167[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	70057958	-	chr21	10706542	+	.	78	26	10698610_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=10698610_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_10706501_10731501_317C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:93 DP:397 GQ:99 PL:[199.5, 0.0, 764.0] SR:26 DR:78 LR:-199.4 LO:218.1);ALT=[chr21:10706542[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	70426185	-	chr7	70438880	+	.	63	61	4941414_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=4941414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_70437501_70462501_254C;SPAN=12695;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:114 DP:45 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:61 DR:63 LR:-336.7 LO:336.7);ALT=[chr7:70438880[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	71211920	+	chr7	71212955	+	.	67	28	4945654_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAAAAGAACC;MAPQ=60;MATEID=4945654_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_71197001_71222001_33C;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:60 GQ:21 PL:[231.0, 21.0, 0.0] SR:28 DR:67 LR:-231.1 LO:231.1);ALT=C[chr7:71212955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	72270265	+	chr7	72275843	+	.	80	29	4951836_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGA;MAPQ=60;MATEID=4951836_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_72275001_72300001_58C;SPAN=5578;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:56 GQ:27 PL:[297.0, 27.0, 0.0] SR:29 DR:80 LR:-297.1 LO:297.1);ALT=A[chr7:72275843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102009660	+	chr7	72355105	+	TATATATATATTTGCTAT	0	25	5091689_1	72.0	.	EVDNC=ASSMB;INSERTION=TATATATATATTTGCTAT;MAPQ=23;MATEID=5091689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_101993501_102018501_62C;SPAN=29654555;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:25 DP:7 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:25 DR:0 LR:-72.62 LO:72.62);ALT=]chr7:102009660]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	73549766	+	chr7	73550967	+	.	29	54	4961001_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTGAGA;MAPQ=60;MATEID=4961001_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_73549001_73574001_263C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:28 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:54 DR:29 LR:-217.9 LO:217.9);ALT=A[chr7:73550967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73828495	+	chr7	73831262	+	.	103	59	4963125_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AGGCCAGGCGCGGTGGCTCACGCCTGTAATCCCAGCACTTTGGGAGGCCGAG;MAPQ=60;MATEID=4963125_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_73818501_73843501_262C;SPAN=2767;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:143 DP:37 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:59 DR:103 LR:-422.5 LO:422.5);ALT=G[chr7:73831262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100185039	+	chr15	52264813	-	.	9	0	8897345_1	22.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=8897345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100185039(+)-15:52264813(+)__15_52258501_52283501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:0 DR:9 LR:-22.12 LO:22.58);ALT=C]chr15:52264813];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	100626435	-	chr7	100627689	+	.	9	0	5085196_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5085196_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100626435(-)-7:100627689(-)__7_100621501_100646501D;SPAN=1254;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:150 GQ:10.9 PL:[0.0, 10.9, 386.1] SR:0 DR:9 LR:10.93 LO:15.37);ALT=[chr7:100627689[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	101001266	+	chr7	101003796	+	.	53	27	5087102_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCAATTTTTGTATTTTT;MAPQ=60;MATEID=5087102_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_7_100989001_101014001_274C;SPAN=2530;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:88 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:27 DR:53 LR:-260.8 LO:260.8);ALT=T[chr7:101003796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101360004	-	chr20	5663475	+	GGCATGATCACAGCTCACTGTAGCCTCGACCTCCTGGGATCAAGAGATGTTCCTGCCTCACCTCCTGAGT	5	97	5089234_1	99.0	.	DISC_MAPQ=18;EVDNC=TSI_L;INSERTION=GGCATGATCACAGCTCACTGTAGCCTCGACCTCCTGGGATCAAGAGATGTTCCTGCCTCACCTCCTGAGT;MAPQ=60;MATEID=5089234_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_7_101356501_101381501_457C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:68 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:97 DR:5 LR:-293.8 LO:293.8);ALT=[chr20:5663475[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	85211624	+	chr7	107829249	+	.	22	30	6992081_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TAAA;MAPQ=60;MATEID=6992081_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_85211001_85236001_218C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:41 DP:75 GQ:65.6 PL:[115.1, 0.0, 65.6] SR:30 DR:22 LR:-115.7 LO:115.7);ALT=]chr11:85211624]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	139451460	+	chr20	36823025	-	.	15	0	10522118_1	17.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=10522118_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:139451460(+)-20:36823025(+)__20_36799001_36824001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:120 GQ:17 PL:[17.0, 0.0, 274.4] SR:0 DR:15 LR:-17.0 LO:30.63);ALT=C]chr20:36823025];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	153757358	+	chr7	153760742	+	.	19	0	5341571_1	38.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=5341571_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:153757358(+)-7:153760742(-)__7_153737501_153762501D;SPAN=3384;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:90 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:0 DR:19 LR:-38.34 LO:43.57);ALT=A[chr7:153760742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	153760751	+	chr7	153757752	+	.	18	0	5341580_1	27.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=5341580_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:153757752(-)-7:153760751(+)__7_153737501_153762501D;SPAN=2999;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:118 GQ:27.5 PL:[27.5, 0.0, 258.5] SR:0 DR:18 LR:-27.45 LO:38.44);ALT=]chr7:153760751]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	99071872	+	chr7	154010815	+	.	16	25	6465134_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CACACACACACACACACACACA;MAPQ=60;MATEID=6465134_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_10_99053501_99078501_301C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:65 GQ:51.8 PL:[104.6, 0.0, 51.8] SR:25 DR:16 LR:-105.4 LO:105.4);ALT=]chr10:99071872]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	154153823	+	chr7	154155071	+	.	153	58	5343096_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAGAAGGAAATA;MAPQ=60;MATEID=5343096_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_154154001_154179001_34C;SPAN=1248;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:186 DP:20 GQ:50.2 PL:[551.2, 50.2, 0.0] SR:58 DR:153 LR:-551.2 LO:551.2);ALT=A[chr7:154155071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	154391960	+	chr7	154399762	+	.	83	0	5344263_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5344263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:154391960(+)-7:154399762(-)__7_154374501_154399501D;SPAN=7802;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:10 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:0 DR:83 LR:-244.3 LO:244.3);ALT=C[chr7:154399762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	155000737	+	chr7	154997565	+	.	10	0	5346024_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5346024_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:154997565(-)-7:155000737(+)__7_154987001_155012001D;SPAN=3172;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:184 GQ:16.6 PL:[0.0, 16.6, 478.6] SR:0 DR:10 LR:16.84 LO:16.64);ALT=]chr7:155000737]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	6833728	+	chr8	6871956	+	.	10	0	5378679_1	18.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=5378679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:6833728(+)-8:6871956(-)__8_6860001_6885001D;SPAN=38228;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:0 DR:10 LR:-18.65 LO:22.38);ALT=A[chr8:6871956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	22414381	+	chr8	7363905	+	TTACATC	13	87	10221089_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;INSERTION=TTACATC;MAPQ=0;MATEID=10221089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_22393001_22418001_240C;SPAN=-1;SUBN=10;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:34 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:87 DR:13 LR:-270.7 LO:270.7);ALT=]chr19:22414381]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	62130611	+	chr8	62132326	-	.	4	3	5485609_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGTTGGTGG;MAPQ=60;MATEID=5485609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_62107501_62132501_292C;SPAN=1715;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:6 DP:72 GQ:0.5 PL:[0.5, 0.0, 172.1] SR:3 DR:4 LR:-0.2994 LO:11.14);ALT=G]chr8:62132326];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	62666696	-	chr19	21890128	+	GATAGGGATAGGGATAGGGATAGGGATAGGGATAGGCATAGGGA	54	115	5486736_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGGGATAGGGATAGGGATAGGGATAGGGATAGGGATAGGGATAGGGATAGGGATAGG;INSERTION=GATAGGGATAGGGATAGGGATAGGGATAGGGATAGGCATAGGGA;MAPQ=60;MATEID=5486736_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_62646501_62671501_322C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:122 DP:44 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:115 DR:54 LR:-359.8 LO:359.8);ALT=[chr19:21890128[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	64318396	+	chr12	32109024	-	.	16	0	7528245_1	34.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=7528245_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:64318396(+)-12:32109024(+)__12_32095001_32120001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:68 GQ:34.4 PL:[34.4, 0.0, 130.1] SR:0 DR:16 LR:-34.39 LO:37.55);ALT=T]chr12:32109024];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	81709320	+	chr20	41696769	+	.	10	0	10550943_1	20.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=10550943_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:81709320(+)-20:41696769(-)__20_41674501_41699501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:0 DR:10 LR:-20.82 LO:23.18);ALT=C[chr20:41696769[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr19	9254189	+	chr8	94654327	+	.	10	0	10145650_1	19.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=10145650_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:94654327(-)-19:9254189(+)__19_9236501_9261501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:52 GQ:19.1 PL:[19.1, 0.0, 104.9] SR:0 DR:10 LR:-18.92 LO:22.47);ALT=]chr19:9254189]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	94654440	+	chr19	9254435	+	.	8	0	10145653_1	10.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=10145653_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:94654440(+)-19:9254435(-)__19_9236501_9261501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=T[chr19:9254435[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	125894597	+	chr8	125895872	-	.	9	0	5677843_1	0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5677843_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:125894597(+)-8:125895872(+)__8_125881001_125906001D;SPAN=1275;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:127 GQ:4.5 PL:[0.0, 4.5, 316.8] SR:0 DR:9 LR:4.698 LO:16.05);ALT=C]chr8:125895872];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	126595129	+	chr8	126601135	+	.	158	64	5680201_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACTCACA;MAPQ=60;MATEID=5680201_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_126591501_126616501_346C;SPAN=6006;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:199 DP:52 GQ:53.8 PL:[590.8, 53.8, 0.0] SR:64 DR:158 LR:-590.8 LO:590.8);ALT=A[chr8:126601135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	32315101	+	chrX	55088086	-	.	9	0	5813702_1	23.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5813702_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:32315101(+)-23:55088086(+)__9_32291001_32316001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:25 GQ:23 PL:[23.0, 0.0, 36.2] SR:0 DR:9 LR:-22.94 LO:23.13);ALT=A]chrX:55088086];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	33621205	+	chr9	33481007	+	.	81	39	5816237_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=5816237_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_9_33614001_33639001_217C;SPAN=140198;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:46 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:39 DR:81 LR:-283.9 LO:283.9);ALT=]chr9:33621205]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	88806038	-	chrX	74928699	+	.	23	14	5915431_1	98.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=TCAACAAAATACTAGCTAACCAAGTCCAACAGC;MAPQ=32;MATEID=5915431_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_88788001_88813001_207C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:51 GQ:22.7 PL:[98.6, 0.0, 22.7] SR:14 DR:23 LR:-100.8 LO:100.8);ALT=[chrX:74928699[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	89154557	+	chr9	89155947	+	TATTGTGGGCCATGCCTTTTGATCATATTAGCTAGCAAGAGCTCCAGGTTTCCTCTCCATAATGAAAATTTTTGAGCCTAACAATAGTCAA	3	101	5916199_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=A;INSERTION=TATTGTGGGCCATGCCTTTTGATCATATTAGCTAGCAAGAGCTCCAGGTTTCCTCTCCATAATGAAAATTTTTGAGCCTAACAATAGTCAA;MAPQ=60;MATEID=5916199_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_89155501_89180501_169C;SPAN=1390;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:101 DP:9 GQ:27 PL:[297.0, 27.0, 0.0] SR:101 DR:3 LR:-297.1 LO:297.1);ALT=T[chr9:89155947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	89201794	+	chr18	40322301	-	.	13	0	10002498_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10002498_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:89201794(+)-18:40322301(+)__18_40302501_40327501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:30 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:0 DR:13 LR:-34.79 LO:34.79);ALT=G]chr18:40322301];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	89206719	-	chr12	6512727	+	.	10	0	7360351_1	16.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7360351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:89206719(-)-12:6512727(-)__12_6492501_6517501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.48 LO:21.7);ALT=[chr12:6512727[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	93179683	+	chr9	90030745	+	.	17	0	5924636_1	47.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=5924636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:90030745(-)-9:93179683(+)__9_93173501_93198501D;SPAN=3148938;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:30 GQ:24.8 PL:[47.9, 0.0, 24.8] SR:0 DR:17 LR:-48.39 LO:48.39);ALT=]chr9:93179683]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	90030923	+	chr9	93179999	+	.	12	0	5924637_1	25.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5924637_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:90030923(+)-9:93179999(-)__9_93173501_93198501D;SPAN=3149076;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=T[chr9:93179999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	90748507	-	chr9	95646288	+	.	13	0	5928806_1	34.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=5928806_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:90748507(-)-9:95646288(-)__9_95623501_95648501D;SPAN=4897781;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:32 GQ:34.4 PL:[34.4, 0.0, 41.0] SR:0 DR:13 LR:-34.24 LO:34.3);ALT=[chr9:95646288[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	90858996	+	chr9	90860964	+	.	79	44	5919750_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTATGTACCTTTT;MAPQ=60;MATEID=5919750_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_90846001_90871001_161C;SPAN=1968;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:28 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:44 DR:79 LR:-293.8 LO:293.8);ALT=T[chr9:90860964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	96470355	+	chr9	96471465	+	.	98	48	5930429_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5930429_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_9_96456501_96481501_210C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:127 DP:21 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:48 DR:98 LR:-376.3 LO:376.3);ALT=C[chr9:96471465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	96500163	+	chr9	96503043	+	.	42	28	5930542_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=ACT;MAPQ=60;MATEID=5930542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_96481001_96506001_233C;SPAN=2880;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:14 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:28 DR:42 LR:-174.9 LO:174.9);ALT=T[chr9:96503043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	98443687	+	chr12	30311079	+	CAGGAGGAACGAACACCTCCAGATGCGCCGCCTTAAGAGCTGTAACACTCACCGAAG	22	248	7515279_1	99.0	.	DISC_MAPQ=4;EVDNC=ASDIS;INSERTION=CAGGAGGAACGAACACCTCCAGATGCGCCGCCTTAAGAGCTGTAACACTCACCGAAG;MAPQ=42;MATEID=7515279_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_30306501_30331501_378C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:261 DP:46 GQ:70.3 PL:[772.3, 70.3, 0.0] SR:248 DR:22 LR:-772.4 LO:772.4);ALT=C[chr12:30311079[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	130917361	+	chr16	9234482	+	.	8	0	9138944_1	18.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=9138944_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:130917361(+)-16:9234482(-)__16_9212001_9237001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=A[chr16:9234482[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	131791289	-	chr9	131793280	+	.	10	0	6009004_1	2.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6009004_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131791289(-)-9:131793280(-)__9_131785501_131810501D;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:113 GQ:2.6 PL:[2.6, 0.0, 269.9] SR:0 DR:10 LR:-2.396 LO:18.83);ALT=[chr9:131793280[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	132026700	+	chr9	132028070	+	.	141	87	6010057_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCTGGGATTACAGGT;MAPQ=60;MATEID=6010057_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132006001_132031001_35C;SPAN=1370;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:197 DP:37 GQ:53.2 PL:[584.2, 53.2, 0.0] SR:87 DR:141 LR:-584.2 LO:584.2);ALT=T[chr9:132028070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132329991	-	chr9	132331171	+	.	10	0	6011454_1	7.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6011454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:132329991(-)-9:132331171(-)__9_132324501_132349501D;SPAN=1180;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:0 DR:10 LR:-7.543 LO:19.68);ALT=[chr9:132331171[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	132829314	+	chr9	132830424	-	.	14	0	6014574_1	16.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6014574_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:132829314(+)-9:132830424(+)__9_132814501_132839501D;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:109 GQ:16.7 PL:[16.7, 0.0, 247.7] SR:0 DR:14 LR:-16.68 LO:28.77);ALT=T]chr9:132830424];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	134638692	-	chr9	134639830	+	.	8	0	6022734_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6022734_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:134638692(-)-9:134639830(-)__9_134627501_134652501D;SPAN=1138;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:136 GQ:10.2 PL:[0.0, 10.2, 349.8] SR:0 DR:8 LR:10.44 LO:13.6);ALT=[chr9:134639830[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	135423182	+	chr9	135421595	+	.	4	8	6026235_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAC;MAPQ=60;MATEID=6026235_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_135411501_135436501_339C;SPAN=1587;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:142 GQ:1.8 PL:[0.0, 1.8, 346.5] SR:8 DR:4 LR:2.16 LO:20.05);ALT=]chr9:135423182]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	135825407	-	chr9	135826467	+	.	2	2	6027972_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GATCCTC;MAPQ=60;MATEID=6027972_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_135803501_135828501_379C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:160 GQ:30.1 PL:[0.0, 30.1, 448.9] SR:2 DR:2 LR:30.14 LO:5.295);ALT=[chr9:135826467[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	136256974	+	chr20	33742105	+	.	8	0	6030845_1	18.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6030845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136256974(+)-20:33742105(-)__9_136244501_136269501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:0 DR:8 LR:-18.55 LO:19.42);ALT=C[chr20:33742105[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	136625194	+	chr9	136626268	+	TGGG	152	110	6031453_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TGGG;MAPQ=60;MATEID=6031453_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_136612001_136637001_30C;SPAN=1074;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:211 DP:44 GQ:56.8 PL:[623.8, 56.8, 0.0] SR:110 DR:152 LR:-623.9 LO:623.9);ALT=G[chr9:136626268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136696117	+	chr11	25269912	+	.	53	0	6673898_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6673898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136696117(+)-11:25269912(-)__11_25259501_25284501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:155 GQ:99 PL:[133.1, 0.0, 242.0] SR:0 DR:53 LR:-133.0 LO:134.7);ALT=A[chr11:25269912[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	12560473	+	chr10	12562974	+	.	52	28	6094205_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTTATTCATTCTT;MAPQ=60;MATEID=6094205_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_10_12544001_12569001_420C;SPAN=2501;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:45 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:28 DR:52 LR:-211.3 LO:211.3);ALT=T[chr10:12562974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	13259268	+	chr10	13260741	+	.	54	26	6096952_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAATGTTAAACCATGGG;MAPQ=60;MATEID=6096952_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_13254501_13279501_344C;SPAN=1473;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:65 DP:89 GQ:25.4 PL:[190.4, 0.0, 25.4] SR:26 DR:54 LR:-197.7 LO:197.7);ALT=G[chr10:13260741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	15957723	+	chr10	15963763	+	.	38	26	6110431_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=GCTGAATTCTCTT;MAPQ=0;MATEID=6110431_2;MATENM=2;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_10_15949501_15974501_243C;SECONDARY;SPAN=6040;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:132 GQ:99 PL:[155.9, 0.0, 162.5] SR:26 DR:38 LR:-155.7 LO:155.7);ALT=T[chr10:15963763[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	15963763	-	chrX	85816922	+	.	6	7	11288553_1	13.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAGAGAATTCAGC;MAPQ=60;MATEID=11288553_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_85799001_85824001_320C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:86 GQ:13.1 PL:[13.1, 0.0, 194.6] SR:7 DR:6 LR:-13.01 LO:22.58);ALT=[chrX:85816922[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	16454892	+	chrX	5708426	+	.	13	0	10946830_1	36.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=10946830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:16454892(+)-23:5708426(-)__23_5708501_5733501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:13 DP:8 GQ:3.3 PL:[36.3, 3.3, 0.0] SR:0 DR:13 LR:-36.31 LO:36.31);ALT=A[chrX:5708426[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	36219661	+	chr10	36221067	+	.	73	52	6198082_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;MAPQ=60;MATEID=6198082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_36211001_36236001_178C;SPAN=1406;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:79 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:52 DR:73 LR:-313.6 LO:313.6);ALT=G[chr10:36221067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25373447	+	chr10	36335211	+	.	2	4	9570937_1	0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TGTC;MAPQ=60;MATEID=9570937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25357501_25382501_83C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:83 GQ:5.7 PL:[0.0, 5.7, 211.2] SR:4 DR:2 LR:5.982 LO:8.55);ALT=]chr17:25373447]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	34535829	+	chr10	37031557	+	.	10	26	10262799_1	94.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GAGGAAGAGGAAGAGGAAGAGGAAGAAGAAGAAGAAGAAGA;MAPQ=60;MATEID=10262799_2;MATENM=8;NM=1;NUMPARTS=2;SCTG=c_19_34520501_34545501_430C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:43 GQ:8.3 PL:[94.1, 0.0, 8.3] SR:26 DR:10 LR:-97.88 LO:97.88);ALT=]chr19:34535829]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	78606897	+	chr10	38285340	+	.	19	0	6375902_1	48.0	.	DISC_MAPQ=5;EVDNC=DSCRD;IMPRECISE;MAPQ=5;MATEID=6375902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38285340(-)-10:78606897(+)__10_78596001_78621001D;SPAN=40321557;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:53 GQ:48.5 PL:[48.5, 0.0, 78.2] SR:0 DR:19 LR:-48.36 LO:48.79);ALT=]chr10:78606897]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38285686	+	chr10	78607478	+	.	27	0	6375903_1	76.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6375903_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38285686(+)-10:78607478(-)__10_78596001_78621001D;SPAN=40321792;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:46 GQ:33.8 PL:[76.7, 0.0, 33.8] SR:0 DR:27 LR:-77.51 LO:77.51);ALT=A[chr10:78607478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	38376500	+	chr10	43055578	-	CCAGGTGCATATTTTCCCCCTCACTTCATTCAGCGCAGCTG	34	45	6207920_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=CCAGGTGCATATTTTCCCCCTCACTTCATTCAGCGCAGCTG;MAPQ=60;MATEID=6207920_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_38367001_38392001_224C;SPAN=4679078;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:53 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:45 DR:34 LR:-211.3 LO:211.3);ALT=C]chr10:43055578];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	38776219	+	chr10	38772625	+	.	10	0	6212257_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6212257_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38772625(-)-10:38776219(+)__10_38759001_38784001D;SPAN=3594;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:164 GQ:11.2 PL:[0.0, 11.2, 419.2] SR:0 DR:10 LR:11.42 LO:17.15);ALT=]chr10:38776219]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38797448	+	chr10	38789722	+	.	12	0	6210829_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6210829_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38789722(-)-10:38797448(+)__10_38783501_38808501D;SPAN=7726;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:12 DP:185 GQ:10.3 PL:[0.0, 10.3, 468.7] SR:0 DR:12 LR:10.51 LO:20.92);ALT=]chr10:38797448]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38875592	+	chr10	38869350	+	.	9	0	6212038_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6212038_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38869350(-)-10:38875592(+)__10_38857001_38882001D;SPAN=6242;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:194 GQ:22.6 PL:[0.0, 22.6, 514.9] SR:0 DR:9 LR:22.85 LO:14.35);ALT=]chr10:38875592]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42357329	+	chr10	42356269	+	.	18	1	6212484_1	0	.	DISC_MAPQ=8;EVDNC=TSI_L;HOMSEQ=ATTCCATTCCATTCCATTCCATTCCATTCC;MAPQ=20;MATEID=6212484_2;MATENM=4;NM=2;NUMPARTS=3;REPSEQ=TTCCATTCCATTCCATTCCATTCCA;SCTG=c_10_42336001_42361001_303C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:19 DP:1219 GQ:99 PL:[0.0, 284.5, 1462.0] SR:1 DR:18 LR:303.7 LO:-5.413);ALT=]chr10:42357329]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42600177	+	chr10	42597585	+	.	8	0	6213701_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6213701_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42597585(-)-10:42600177(+)__10_42581001_42606001D;SPAN=2592;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:419 GQ:86.9 PL:[0.0, 86.9, 1192.0] SR:0 DR:8 LR:87.11 LO:9.662);ALT=]chr10:42600177]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42666935	+	chr10	42661706	+	.	14	0	6216180_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6216180_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42661706(-)-10:42666935(+)__10_42654501_42679501D;SPAN=5229;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:14 DP:202 GQ:8.2 PL:[0.0, 8.2, 505.0] SR:0 DR:14 LR:8.513 LO:24.82);ALT=]chr10:42666935]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42701593	+	chr10	42716849	+	.	21	0	6215804_1	62.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=6215804_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42701593(+)-10:42716849(-)__10_42679001_42704001D;SPAN=15256;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:27 GQ:2.6 PL:[62.0, 0.0, 2.6] SR:0 DR:21 LR:-65.13 LO:65.13);ALT=G[chr10:42716849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43272230	-	chr20	14961673	+	.	11	46	6218744_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6218744_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_43267001_43292001_393C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:72 GQ:10.4 PL:[162.2, 0.0, 10.4] SR:46 DR:11 LR:-169.6 LO:169.6);ALT=[chr20:14961673[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	54783542	+	chr10	54788830	+	T	78	64	6273873_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=6273873_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_54782001_54807001_67C;SPAN=5288;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:94 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:64 DR:78 LR:-333.4 LO:333.4);ALT=A[chr10:54788830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	55038596	+	chr20	47845568	+	.	9	32	6274225_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=6274225_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_10_55027001_55052001_268C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:38 DP:35 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:32 DR:9 LR:-112.2 LO:112.2);ALT=T[chr20:47845568[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	55038800	-	chr19	37433289	+	.	9	0	6274227_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6274227_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:55038800(-)-19:37433289(-)__10_55027001_55052001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=[chr19:37433289[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	55271528	+	chr10	107230662	+	.	4	88	6275624_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACACACACACACACACA;MAPQ=60;MATEID=6275624_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_55247501_55272501_277C;SPAN=51959134;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:86 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:88 DR:4 LR:-267.4 LO:267.4);ALT=A[chr10:107230662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	33595145	+	chr10	55894133	+	TATATATATATAA	9	46	9981844_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=TATATATATATAA;MAPQ=60;MATEID=9981844_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_33589501_33614501_140C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:85 GQ:66.2 PL:[138.8, 0.0, 66.2] SR:46 DR:9 LR:-140.0 LO:140.0);ALT=]chr18:33595145]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	56767191	-	chr10	56773197	+	.	124	106	6280440_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=6280440_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_10_56766501_56791501_184C;SPAN=6006;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:198 DP:63 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:106 DR:124 LR:-587.5 LO:587.5);ALT=[chr10:56773197[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	63034905	+	chr19	19996063	-	.	3	8	10207617_1	8.0	.	DISC_MAPQ=0;EVDNC=TSI_L;HOMSEQ=TTTCTTTCTTTCTTTCTTTCTTT;MAPQ=60;MATEID=10207617_2;MATENM=2;NM=0;NUMPARTS=3;REPSEQ=TTCTTTCTTTCTTTCTTTCT;SCTG=c_19_19992001_20017001_482C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:17 GQ:4 PL:[8.1, 0.0, 4.0] SR:8 DR:3 LR:-8.033 LO:8.033);ALT=A]chr19:19996063];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	74767593	-	chr17	32673409	+	ATACATCC	49	48	6357300_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=ATACATCC;MAPQ=60;MATEID=6357300_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_10_74749501_74774501_37C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:89 DP:116 GQ:18.2 PL:[262.4, 0.0, 18.2] SR:48 DR:49 LR:-274.8 LO:274.8);ALT=[chr17:32673409[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	74784036	+	chr10	74788477	+	.	32	0	6357513_1	74.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=6357513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:74784036(+)-10:74788477(-)__10_74774001_74799001D;SPAN=4441;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:117 GQ:74 PL:[74.0, 0.0, 209.3] SR:0 DR:32 LR:-73.93 LO:77.56);ALT=T[chr10:74788477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75848405	+	chr10	75781766	+	.	4	7	6362570_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=6362570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_75778501_75803501_75C;SPAN=66639;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:70 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:7 DR:4 LR:-10.74 LO:18.5);ALT=]chr10:75848405]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	75820294	+	chr10	75821799	-	.	5	2	6362368_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTACAGG;MAPQ=60;MATEID=6362368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_75803001_75828001_454C;SPAN=1505;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:149 GQ:20.5 PL:[0.0, 20.5, 402.6] SR:2 DR:5 LR:20.56 LO:9.19);ALT=G]chr10:75821799];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	76355531	-	chr20	4351297	+	.	47	16	6365595_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=GATCACCTGAGGTCAGGAATTCGAGACCAGCCTGGCCAACA;MAPQ=60;MATEID=6365595_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_10_76342001_76367001_393C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:62 DP:16 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:16 DR:47 LR:-181.5 LO:181.5);ALT=[chr20:4351297[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	77347393	+	chr10	77345742	+	.	91	36	6369869_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GTTG;MAPQ=60;MATEID=6369869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_77346501_77371501_279C;SPAN=1651;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:84 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:36 DR:91 LR:-316.9 LO:316.9);ALT=]chr10:77347393]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	78255578	+	chr10	78261020	+	.	120	80	6373650_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTCAGT;MAPQ=60;MATEID=6373650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_78253001_78278001_239C;SPAN=5442;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:164 DP:34 GQ:44.2 PL:[485.2, 44.2, 0.0] SR:80 DR:120 LR:-485.2 LO:485.2);ALT=T[chr10:78261020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78346604	+	chr10	78351578	+	.	58	43	6374657_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAATACTTAATTT;MAPQ=60;MATEID=6374657_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_78351001_78376001_49C;SPAN=4974;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:31 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:43 DR:58 LR:-237.7 LO:237.7);ALT=T[chr10:78351578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	79184905	+	chr22	44376043	-	.	6	30	6377270_1	69.0	.	DISC_MAPQ=5;EVDNC=ASDIS;HOMSEQ=ATGGATGGATGGATGGATGGATGGATG;MAPQ=23;MATEID=6377270_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_10_79184001_79209001_182C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:158 GQ:69.5 PL:[69.5, 0.0, 313.7] SR:30 DR:6 LR:-69.43 LO:78.28);ALT=G]chr22:44376043];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	99034873	+	chr10	99037398	+	.	195	86	6464317_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAAAGCACTG;MAPQ=60;MATEID=6464317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_99029001_99054001_296C;SPAN=2525;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:245 DP:45 GQ:66.1 PL:[726.1, 66.1, 0.0] SR:86 DR:195 LR:-726.2 LO:726.2);ALT=G[chr10:99037398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	99174549	-	chr10	99176031	+	.	8	0	6464924_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6464924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:99174549(-)-10:99176031(-)__10_99151501_99176501D;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:159 GQ:16.6 PL:[0.0, 16.6, 419.2] SR:0 DR:8 LR:16.67 LO:13.04);ALT=[chr10:99176031[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	100057897	-	chr17	68088708	+	.	4	49	9788136_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TATCTATCTATCTATCTATCTATCTATCTATCTATCTATCTAT;MAPQ=49;MATEID=9788136_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_17_68085501_68110501_90C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:38 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:49 DR:4 LR:-155.1 LO:155.1);ALT=[chr17:68088708[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	394278	+	chr11	392811	+	A	6	14	6618321_1	45.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=6618321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_392001_417001_80C;SPAN=1467;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:14 DR:6 LR:-45.01 LO:45.06);ALT=]chr11:394278]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	736910	+	chr11	3917284	+	.	9	0	6627260_1	16.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=6627260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:736910(+)-11:3917284(-)__11_3895501_3920501D;SPAN=3180374;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=T[chr11:3917284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	3917414	+	chr11	737067	+	.	41	32	6627261_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAAAGTGCTGGGATTACAGGCG;MAPQ=60;MATEID=6627261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_3895501_3920501_285C;SPAN=3180347;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:56 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:32 DR:41 LR:-178.2 LO:178.2);ALT=]chr11:3917414]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	3416273	-	chr11	3615604	+	.	3	2	6626485_1	5.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=CCAGGGGCA;MAPQ=50;MATEID=6626485_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_3601501_3626501_280C;SPAN=199331;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:4 DP:28 GQ:5.6 PL:[5.6, 0.0, 61.7] SR:2 DR:3 LR:-5.618 LO:8.419);ALT=[chr11:3615604[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	3615290	+	chr11	71310881	-	.	8	0	6626514_1	16.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6626514_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:3615290(+)-11:71310881(+)__11_3601501_3626501D;SPAN=67695591;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:0 DR:8 LR:-16.11 LO:18.33);ALT=C]chr11:71310881];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	24137201	-	chr11	87594960	+	.	47	43	6665375_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=6665375_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_24132501_24157501_11C;SPAN=63457759;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:66 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:43 DR:47 LR:-221.2 LO:221.2);ALT=[chr11:87594960[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	87594964	+	chr11	24137280	+	.	150	67	7008120_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTA;MAPQ=60;MATEID=7008120_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_87587501_87612501_793C;SPAN=63457684;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:196 DP:200 GQ:54.1 PL:[594.1, 54.1, 0.0] SR:67 DR:150 LR:-594.1 LO:594.1);ALT=]chr11:87594964]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	24137288	+	chr11	98883067	+	.	47	69	7156446_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7156446_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_98882001_98907001_64C;SPAN=74745779;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:80 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:69 DR:47 LR:-340.0 LO:340.0);ALT=G[chr11:98883067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	24137851	-	chr11	24139485	+	CTCTCTTAG	13	86	6665387_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CTCTCTTAG;MAPQ=60;MATEID=6665387_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_11_24132501_24157501_235C;SPAN=1634;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:277 GQ:99 PL:[245.2, 0.0, 426.8] SR:86 DR:13 LR:-245.2 LO:247.9);ALT=[chr11:24139485[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	24137948	+	chr11	98883577	-	.	37	51	6665389_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=6665389_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_24132501_24157501_194C;SPAN=74745629;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:68 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:51 DR:37 LR:-241.0 LO:241.0);ALT=A]chr11:98883577];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	28622230	+	chr11	24139182	+	.	190	49	6709086_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=6709086_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_28616001_28641001_391C;SPAN=4483048;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:204 DP:89 GQ:55 PL:[604.0, 55.0, 0.0] SR:49 DR:190 LR:-604.0 LO:604.0);ALT=]chr11:28622230]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	24349495	+	chr11	24355549	+	.	40	27	6667198_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAACAGAACCC;MAPQ=60;MATEID=6667198_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_24328501_24353501_145C;SPAN=6054;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:102 GQ:99 PL:[140.9, 0.0, 104.6] SR:27 DR:40 LR:-141.0 LO:141.0);ALT=C[chr11:24355549[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	25493241	+	chr11	25494361	+	.	0	51	6676200_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AATTTT;MAPQ=60;MATEID=6676200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_25480001_25505001_191C;SPAN=1120;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:219 GQ:99 PL:[109.0, 0.0, 422.6] SR:51 DR:0 LR:-109.0 LO:119.4);ALT=T[chr11:25494361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	96270545	+	chr11	25752249	+	CAT	49	23	6679352_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CAT;MAPQ=60;MATEID=6679352_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_11_25749501_25774501_104C;SPAN=70518296;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:61 DP:164 GQ:99 PL:[157.1, 0.0, 239.6] SR:23 DR:49 LR:-156.9 LO:157.9);ALT=]chr11:96270545]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	26800268	+	chr11	86700710	-	.	180	53	7002686_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=7002686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_86681001_86706001_690C;SPAN=59900442;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:214 DP:111 GQ:57.7 PL:[633.7, 57.7, 0.0] SR:53 DR:180 LR:-633.8 LO:633.8);ALT=A]chr11:86700710];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	28082157	+	chr11	26929534	+	TGCACAGCCAAACACTATG	173	77	6692844_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TGCACAGCCAAACACTATG;MAPQ=60;MATEID=6692844_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_26925501_26950501_726C;SPAN=1152623;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:212 DP:282 GQ:59.2 PL:[623.6, 0.0, 59.2] SR:77 DR:173 LR:-650.5 LO:650.5);ALT=]chr11:28082157]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	26958398	-	chr11	26959867	+	.	8	0	6692358_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6692358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:26958398(-)-11:26959867(-)__11_26950001_26975001D;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:813 GQ:99 PL:[0.0, 193.4, 2360.0] SR:0 DR:8 LR:193.9 LO:7.415);ALT=[chr11:26959867[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	97311967	+	chr11	27035783	+	.	138	52	7141563_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7141563_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_97289501_97314501_606C;SPAN=70276184;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:166 DP:165 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:52 DR:138 LR:-491.8 LO:491.8);ALT=]chr11:97311967]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	27187962	-	chr11	95942887	+	.	225	87	7125332_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7125332_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_95942001_95967001_373C;SPAN=68754925;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:281 DP:97 GQ:75.8 PL:[831.8, 75.8, 0.0] SR:87 DR:225 LR:-831.8 LO:831.8);ALT=[chr11:95942887[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	27221064	+	chr11	28082681	-	.	161	69	6703957_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=6703957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_28077001_28102001_354C;SPAN=861617;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:216 DP:241 GQ:64.9 PL:[712.9, 64.9, 0.0] SR:69 DR:161 LR:-710.4 LO:710.4);ALT=T]chr11:28082681];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	29931676	+	chr11	27273999	+	.	216	61	6715356_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=6715356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_29914501_29939501_77C;SPAN=2657677;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:235 DP:137 GQ:63.4 PL:[696.4, 63.4, 0.0] SR:61 DR:216 LR:-696.5 LO:696.5);ALT=]chr11:29931676]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	27796415	+	chr11	92124130	+	.	137	49	7083758_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7083758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_92120001_92145001_761C;SPAN=64327715;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:166 DP:347 GQ:99 PL:[454.0, 0.0, 388.0] SR:49 DR:137 LR:-454.2 LO:454.2);ALT=T[chr11:92124130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	28057512	+	chr11	28056253	+	.	22	0	6707894_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6707894_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:28056253(-)-11:28057512(+)__11_28052501_28077501D;SPAN=1259;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:22 DP:919 GQ:99 PL:[0.0, 176.1, 2584.0] SR:0 DR:22 LR:176.4 LO:28.71);ALT=]chr11:28057512]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	28116978	+	chr11	91209154	+	.	134	55	7068913_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GAC;MAPQ=60;MATEID=7068913_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_91189001_91214001_598C;SPAN=63092176;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:161 DP:242 GQ:99 PL:[466.1, 0.0, 119.5] SR:55 DR:134 LR:-477.2 LO:477.2);ALT=C[chr11:91209154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	28462216	-	chr11	96559642	+	.	115	36	7132149_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAT;MAPQ=60;MATEID=7132149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_96554501_96579501_776C;SPAN=68097426;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:137 DP:156 GQ:32.2 PL:[442.3, 32.2, 0.0] SR:36 DR:115 LR:-445.3 LO:445.3);ALT=[chr11:96559642[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	29007245	+	chr11	29012888	+	.	37	0	6711148_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6711148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:29007245(+)-11:29012888(-)__11_28983501_29008501D;SPAN=5643;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:37 DP:30 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:0 DR:37 LR:-108.9 LO:108.9);ALT=C[chr11:29012888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	29559730	+	chr11	29562002	+	ATAATAAATT	78	54	6712893_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ATAATAAATT;MAPQ=60;MATEID=6712893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_29547001_29572001_109C;SPAN=2272;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:102 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:54 DR:78 LR:-310.3 LO:310.3);ALT=G[chr11:29562002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94913814	+	chr11	29832425	+	.	254	87	7118442_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=7118442_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_94913001_94938001_133C;SPAN=65081389;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:303 DP:93 GQ:81.8 PL:[897.8, 81.8, 0.0] SR:87 DR:254 LR:-897.8 LO:897.8);ALT=]chr11:94913814]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	30537132	+	chr11	30565853	-	.	4	3	6718373_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=6718373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_30527001_30552001_426C;SPAN=28721;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:80 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:3 DR:4 LR:5.169 LO:8.632);ALT=A]chr11:30565853];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	31617372	+	chr11	31620114	+	.	0	63	6721866_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GCA;MAPQ=60;MATEID=6721866_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_31605001_31630001_302C;SPAN=2742;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:108 GQ:83 PL:[178.7, 0.0, 83.0] SR:63 DR:0 LR:-180.6 LO:180.6);ALT=A[chr11:31620114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	91209132	+	chr11	32378981	+	.	152	59	7068914_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7068914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_91189001_91214001_647C;SPAN=58830151;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:182 DP:246 GQ:62.2 PL:[534.2, 0.0, 62.2] SR:59 DR:152 LR:-555.7 LO:555.7);ALT=]chr11:91209132]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	32566061	+	chr11	95225383	+	.	145	60	6726963_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6726963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_32560501_32585501_12C;SPAN=62659322;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:189 DP:99 GQ:51.1 PL:[561.1, 51.1, 0.0] SR:60 DR:145 LR:-561.1 LO:561.1);ALT=T[chr11:95225383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	70950376	+	chr11	70951826	-	.	3	2	6901132_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGCCAGG;MAPQ=60;MATEID=6901132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_70927501_70952501_167C;SPAN=1450;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:193 GQ:35.5 PL:[0.0, 35.5, 538.0] SR:2 DR:3 LR:35.78 LO:6.696);ALT=T]chr11:70951826];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	71279868	-	chr11	71290883	+	.	23	0	6902971_1	19.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=6902971_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:71279868(-)-11:71290883(-)__11_71270501_71295501D;SPAN=11015;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:208 GQ:19.6 PL:[19.6, 0.0, 485.0] SR:0 DR:23 LR:-19.57 LO:45.66);ALT=[chr11:71290883[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	52178115	+	chr11	74064909	+	.	3	77	6925536_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGGGTGGCTGCCGGGCGGGGGCTG;MAPQ=60;MATEID=6925536_2;MATENM=7;NM=0;NUMPARTS=2;SCTG=c_11_74063501_74088501_442C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:68 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:77 DR:3 LR:-234.4 LO:234.4);ALT=]chr15:52178115]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	78024273	+	chr11	76746553	+	.	38	47	6947957_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=6947957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_76734001_76759001_456C;SPAN=1277720;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:82 DP:180 GQ:99 PL:[221.9, 0.0, 215.3] SR:47 DR:38 LR:-221.9 LO:221.9);ALT=]chr11:78024273]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	76746553	-	chr11	78024331	+	GGATCACTCTAAAGCTTTTTTTTTCCCAGCACTTTTTTTTTCAGTT	113	120	6962192_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTT;INSERTION=GGATCACTCTAAAGCTTTTTTTTTCCCAGCACTTTTTTTTTCAGTT;MAPQ=60;MATEID=6962192_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_78008001_78033001_528C;SPAN=1277778;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:214 DP:131 GQ:57.7 PL:[633.7, 57.7, 0.0] SR:120 DR:113 LR:-633.8 LO:633.8);ALT=[chr11:78024331[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	76959289	-	chrX	47119458	+	.	3	4	6951018_1	0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=TGAGCTGAGATTGCACCACTGCACTCCAGCCTGG;MAPQ=51;MATEID=6951018_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_76954501_76979501_868C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:252 GQ:48.1 PL:[0.0, 48.1, 706.3] SR:4 DR:3 LR:48.47 LO:7.816);ALT=[chrX:47119458[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	77119794	+	chr11	77167712	-	.	126	53	6955182_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6955182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77150501_77175501_723C;SPAN=47918;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:164 DP:112 GQ:44.2 PL:[485.2, 44.2, 0.0] SR:53 DR:126 LR:-485.2 LO:485.2);ALT=A]chr11:77167712];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	77886100	-	chr11	77889450	+	.	8	0	6960645_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6960645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:77886100(-)-11:77889450(-)__11_77885501_77910501D;SPAN=3350;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:286 GQ:50.9 PL:[0.0, 50.9, 795.4] SR:0 DR:8 LR:51.08 LO:10.98);ALT=[chr11:77889450[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	78772191	+	chr11	79022582	-	.	226	59	6972254_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=6972254_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_79012501_79037501_352C;SPAN=250391;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:270 DP:66 GQ:73 PL:[802.0, 73.0, 0.0] SR:59 DR:226 LR:-802.1 LO:802.1);ALT=A]chr11:79022582];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	92488775	+	chr11	79005423	+	AAAC	71	29	7092821_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AAAC;MAPQ=60;MATEID=7092821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_92487501_92512501_1101C;SPAN=13483352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:84 DP:312 GQ:99 PL:[193.0, 0.0, 562.7] SR:29 DR:71 LR:-192.8 LO:202.9);ALT=]chr11:92488775]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	84723396	-	chr15	90114725	+	.	18	71	6989613_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CCATTTCTACTAAAAATACAAAATT;MAPQ=60;MATEID=6989613_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_84721001_84746001_29C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:34 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:71 DR:18 LR:-237.7 LO:237.7);ALT=[chr15:90114725[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	85199785	+	chr11	86907737	+	AGAGCTCTCAAAAAAAT	37	16	7004101_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AGAGCTCTCAAAAAAAT;MAPQ=60;MATEID=7004101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_86901501_86926501_470C;SPAN=1707952;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:48 DP:71 GQ:30.5 PL:[139.4, 0.0, 30.5] SR:16 DR:37 LR:-142.9 LO:142.9);ALT=T[chr11:86907737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85310436	-	chr11	85312027	+	.	8	0	6992495_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6992495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85310436(-)-11:85312027(-)__11_85309001_85334001D;SPAN=1591;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:130 GQ:8.7 PL:[0.0, 8.7, 333.3] SR:0 DR:8 LR:8.812 LO:13.76);ALT=[chr11:85312027[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	86120028	-	chr11	88865273	+	.	165	58	7024244_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7024244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_88861501_88886501_146C;SPAN=2745245;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:206 DP:146 GQ:55.6 PL:[610.6, 55.6, 0.0] SR:58 DR:165 LR:-610.7 LO:610.7);ALT=[chr11:88865273[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	88642548	+	chr11	96184889	+	.	91	37	7129015_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7129015_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_96162501_96187501_877C;SPAN=7542341;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:111 DP:272 GQ:99 PL:[292.9, 0.0, 365.6] SR:37 DR:91 LR:-292.7 LO:293.2);ALT=T[chr11:96184889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	88964485	+	chr11	88967931	+	.	156	108	7025014_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TGT;MAPQ=60;MATEID=7025014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_88959501_88984501_562C;SPAN=3446;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:254 DP:176 GQ:68.5 PL:[752.5, 68.5, 0.0] SR:108 DR:156 LR:-752.6 LO:752.6);ALT=T[chr11:88967931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	90065772	+	chr11	89168420	+	.	135	36	7029067_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=7029067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_89155501_89180501_642C;SPAN=897352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:154 DP:232 GQ:99 PL:[445.7, 0.0, 115.6] SR:36 DR:135 LR:-456.1 LO:456.1);ALT=]chr11:90065772]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	89908896	+	chr11	89916290	+	.	12	7	7047782_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=7047782_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_89890501_89915501_282C;SPAN=7394;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:215 GQ:1.3 PL:[1.3, 0.0, 519.5] SR:7 DR:12 LR:-1.169 LO:33.45);ALT=A[chr11:89916290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	95417865	+	chr11	90315029	+	T	159	65	7122454_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=T;MAPQ=56;MATEID=7122454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_95403001_95428001_350C;SPAN=5102836;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:196 DP:110 GQ:52.9 PL:[580.9, 52.9, 0.0] SR:65 DR:159 LR:-580.9 LO:580.9);ALT=]chr11:95417865]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	92501163	+	chr11	98883386	+	ATGGTTTGGCT	136	37	7093106_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ATGGTTTGGCT;MAPQ=60;MATEID=7093106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_92487501_92512501_764C;SPAN=6382223;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:163 DP:206 GQ:16.9 PL:[482.3, 0.0, 16.9] SR:37 DR:136 LR:-508.4 LO:508.4);ALT=C[chr11:98883386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	92869804	+	chr11	92875914	+	ATACATAAC	38	47	7096593_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=ATACATAAC;MAPQ=60;MATEID=7096593_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_92855001_92880001_562C;SPAN=6110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:85 DP:188 GQ:99 PL:[229.7, 0.0, 226.4] SR:47 DR:38 LR:-229.7 LO:229.7);ALT=T[chr11:92875914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93021139	+	chr11	93022161	+	A	0	52	7098492_1	90.0	.	EVDNC=ASSMB;INSERTION=A;MAPQ=60;MATEID=7098492_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_93002001_93027001_589C;SPAN=1022;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:301 GQ:90.4 PL:[90.4, 0.0, 638.3] SR:52 DR:0 LR:-90.1 LO:114.2);ALT=T[chr11:93022161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93486679	+	chr11	94912201	+	TTTAACTAG	115	59	7119493_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TTTAACTAG;MAPQ=60;MATEID=7119493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_94888501_94913501_28C;SPAN=1425522;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:148 DP:160 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:59 DR:115 LR:-475.3 LO:475.3);ALT=A[chr11:94912201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93679244	+	chr11	93681424	+	.	165	106	7108059_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCCTGTTGGATTCTT;MAPQ=60;MATEID=7108059_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_11_93663501_93688501_43C;SPAN=2180;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:217 DP:112 GQ:58.6 PL:[643.6, 58.6, 0.0] SR:106 DR:165 LR:-643.7 LO:643.7);ALT=T[chr11:93681424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93695221	+	chr11	93702085	+	.	66	55	7108429_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=7108429_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_93688001_93713001_504C;SPAN=6864;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:95 DP:214 GQ:99 PL:[255.8, 0.0, 262.4] SR:55 DR:66 LR:-255.6 LO:255.6);ALT=T[chr11:93702085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94970456	-	chr11	97111810	+	.	60	61	7139217_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=7139217_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_97093501_97118501_142C;SPAN=2141354;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:107 DP:162 GQ:81.8 PL:[309.5, 0.0, 81.8] SR:61 DR:60 LR:-316.5 LO:316.5);ALT=[chr11:97111810[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	95169380	+	chr11	95175432	+	.	47	51	7120316_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=7120316_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_11_95158001_95183001_96C;SPAN=6052;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:81 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:51 DR:47 LR:-247.6 LO:247.6);ALT=A[chr11:95175432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	95220767	-	chr11	97657269	+	.	68	33	7144793_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7144793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_97657001_97682001_689C;SPAN=2436502;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:93 DP:151 GQ:98 PL:[266.3, 0.0, 98.0] SR:33 DR:68 LR:-270.2 LO:270.2);ALT=[chr11:97657269[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	95746463	+	chr11	96870992	-	T	106	34	7125098_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=7125098_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_95721501_95746501_3C;SPAN=1124529;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:133 DP:46 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:34 DR:106 LR:-392.8 LO:392.8);ALT=A]chr11:96870992];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	96265856	+	chr11	96270636	-	.	19	49	7128787_1	86.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TGT;MAPQ=60;MATEID=7128787_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_96260501_96285501_318C;SPAN=4780;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:59 DP:399 GQ:86.7 PL:[86.7, 0.0, 882.2] SR:49 DR:19 LR:-86.66 LO:125.1);ALT=A]chr11:96270636];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	98880329	+	chr11	98883386	-	GATTTT	162	64	7157820_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GATTTT;MAPQ=60;MATEID=7157820_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_98857501_98882501_52C;SPAN=3057;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:214 DP:64 GQ:57.7 PL:[633.7, 57.7, 0.0] SR:64 DR:162 LR:-633.8 LO:633.8);ALT=A]chr11:98883386];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	99762143	+	chr11	99766003	+	.	64	51	7158723_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=7158723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_99764001_99789001_170C;SPAN=3860;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:11 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:51 DR:64 LR:-254.2 LO:254.2);ALT=A[chr11:99766003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	117920353	+	chr15	57019427	-	.	14	0	7206925_1	18.0	.	DISC_MAPQ=7;EVDNC=DSCRD;IMPRECISE;MAPQ=7;MATEID=7206925_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:117920353(+)-15:57019427(+)__11_117918501_117943501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:0 DR:14 LR:-18.58 LO:29.2);ALT=C]chr15:57019427];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	118293109	-	chr11	118295524	+	.	9	0	7210673_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7210673_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118293109(-)-11:118295524(-)__11_118286001_118311001D;SPAN=2415;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:140 GQ:8.1 PL:[0.0, 8.1, 356.4] SR:0 DR:9 LR:8.221 LO:15.65);ALT=[chr11:118295524[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	118707030	-	chr11	118708219	+	.	14	0	7213090_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7213090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118707030(-)-11:118708219(-)__11_118702501_118727501D;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:14 DP:205 GQ:9.1 PL:[0.0, 9.1, 514.9] SR:0 DR:14 LR:9.326 LO:24.73);ALT=[chr11:118708219[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	119082238	+	chr11	118842623	+	.	69	25	7217161_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7217161_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_119070001_119095001_568C;SPAN=239615;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:77 DP:109 GQ:39.8 PL:[224.6, 0.0, 39.8] SR:25 DR:69 LR:-232.0 LO:232.0);ALT=]chr11:119082238]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	119440683	+	chr16	72158099	+	TTTGTAGAGGC	10	55	7219882_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=TTTGTAGAGGC;MAPQ=60;MATEID=7219882_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_119437501_119462501_199C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:41 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:55 DR:10 LR:-171.6 LO:171.6);ALT=T[chr16:72158099[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	119956131	+	chr11	119954127	+	.	64	0	7223094_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=7223094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:119954127(-)-11:119956131(+)__11_119952001_119977001D;SPAN=2004;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:194 GQ:99 PL:[158.9, 0.0, 310.7] SR:0 DR:64 LR:-158.7 LO:161.4);ALT=]chr11:119956131]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	120674468	+	chr11	120792878	+	.	221	70	7227365_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TATTT;MAPQ=53;MATEID=7227365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_120785001_120810001_120C;SPAN=118410;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:249 DP:29 GQ:67.3 PL:[739.3, 67.3, 0.0] SR:70 DR:221 LR:-739.4 LO:739.4);ALT=T[chr11:120792878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6643735	+	chrX	39647397	-	CCGAGCCACATCGCTC	5	96	11093637_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;INSERTION=CCGAGCCACATCGCTC;MAPQ=60;MATEID=11093637_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_23_39641001_39666001_92C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:122 GQ:3 PL:[300.3, 3.0, 0.0] SR:96 DR:5 LR:-315.7 LO:315.7);ALT=G]chrX:39647397];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	9016803	+	chr12	9018144	-	.	4	2	7379535_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=7379535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9016001_9041001_112C;SPAN=1341;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:201 GQ:34.3 PL:[0.0, 34.3, 554.5] SR:2 DR:4 LR:34.65 LO:8.405);ALT=T]chr12:9018144];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	9016852	+	chr12	9017868	+	.	121	129	7379537_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCTCATGCCTGT;MAPQ=60;MATEID=7379537_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_9016001_9041001_344C;SPAN=1016;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:228 DP:76 GQ:61.6 PL:[676.6, 61.6, 0.0] SR:129 DR:121 LR:-676.7 LO:676.7);ALT=T[chr12:9017868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9304760	+	chr12	9243514	+	.	49	26	7381711_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GTT;MAPQ=60;MATEID=7381711_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9285501_9310501_469C;SPAN=61246;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:67 DP:104 GQ:57.8 PL:[193.1, 0.0, 57.8] SR:26 DR:49 LR:-196.9 LO:196.9);ALT=]chr12:9304760]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	9632754	+	chr12	31353964	-	.	27	0	7522211_1	65.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=7522211_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:9632754(+)-12:31353964(+)__12_31335501_31360501D;SPAN=21721210;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:89 GQ:65 PL:[65.0, 0.0, 150.8] SR:0 DR:27 LR:-65.02 LO:66.9);ALT=T]chr12:31353964];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	11192447	+	chr12	11218062	+	.	131	78	7394220_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTC;MAPQ=60;MATEID=7394220_2;MATENM=11;NM=1;NUMPARTS=2;SCTG=c_12_11196501_11221501_190C;SPAN=25615;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:166 DP:139 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:78 DR:131 LR:-491.8 LO:491.8);ALT=C[chr12:11218062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	29844030	+	chr12	29846435	+	.	22	0	7512013_1	37.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7512013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:29844030(+)-12:29846435(-)__12_29841001_29866001D;SPAN=2405;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:132 GQ:37.1 PL:[37.1, 0.0, 281.3] SR:0 DR:22 LR:-36.86 LO:47.92);ALT=C[chr12:29846435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	29844384	+	chr12	29846436	+	.	154	158	7512017_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAC;MAPQ=60;MATEID=7512017_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_29841001_29866001_225C;SPAN=2052;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:258 DP:62 GQ:69.7 PL:[765.7, 69.7, 0.0] SR:158 DR:154 LR:-765.8 LO:765.8);ALT=C[chr12:29846436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	30237245	+	chr12	30243567	+	AACA	4	159	7514330_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AACA;MAPQ=60;MATEID=7514330_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_30233001_30258001_95C;SPAN=6322;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:161 DP:62 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:159 DR:4 LR:-475.3 LO:475.3);ALT=T[chr12:30243567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	30518417	-	chr12	30519480	+	.	2	3	7515905_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTGTTG;MAPQ=60;MATEID=7515905_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_30502501_30527501_311C;SPAN=1063;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:251 GQ:54.4 PL:[0.0, 54.4, 716.2] SR:3 DR:2 LR:54.8 LO:4.522);ALT=[chr12:30519480[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr21	25532815	+	chr12	30627432	+	.	0	11	7516629_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CCCG;MAPQ=51;MATEID=7516629_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_30625001_30650001_250C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:131 GQ:1.1 PL:[1.1, 0.0, 314.6] SR:11 DR:0 LR:-0.8199 LO:20.45);ALT=]chr21:25532815]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	31944043	+	chr12	31956007	-	CTGTA	3	5	7527085_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGTA;MAPQ=60;MATEID=7527085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_31923501_31948501_206C;SPAN=11964;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:7 DP:115 GQ:7.8 PL:[0.0, 7.8, 293.7] SR:5 DR:3 LR:8.049 LO:12.0);ALT=T]chr12:31956007];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	43461084	+	chr12	43462661	+	ATAA	0	57	7569940_1	99.0	.	EVDNC=ASSMB;INSERTION=ATAA;MAPQ=60;MATEID=7569940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_43438501_43463501_111C;SPAN=1577;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:57 DP:85 GQ:39.8 PL:[165.2, 0.0, 39.8] SR:57 DR:0 LR:-169.3 LO:169.3);ALT=A[chr12:43462661[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	43977460	+	chr12	43979550	+	.	69	42	7572099_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAGACATTCCA;MAPQ=60;MATEID=7572099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_43977501_44002501_1C;SPAN=2090;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:52 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:42 DR:69 LR:-277.3 LO:277.3);ALT=A[chr12:43979550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53258192	-	chr12	65905635	+	.	7	9	7673148_1	8.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CTA;MAPQ=60;MATEID=7673148_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_65905001_65930001_14C;SPAN=12647443;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:127 GQ:8.6 PL:[8.6, 0.0, 299.0] SR:9 DR:7 LR:-8.506 LO:25.35);ALT=[chr12:65905635[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	76361989	+	chr12	58469539	+	.	26	0	7640902_1	74.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7640902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:58469539(-)-23:76361989(+)__12_58457001_58482001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:42 GQ:25.1 PL:[74.6, 0.0, 25.1] SR:0 DR:26 LR:-75.63 LO:75.63);ALT=]chrX:76361989]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	64667225	+	chr12	77771324	-	.	64	37	7765437_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=7765437_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_77763001_77788001_38C;SPAN=13104099;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:47 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:37 DR:64 LR:-277.3 LO:277.3);ALT=T]chr12:77771324];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	64756658	-	chr12	79558633	+	.	28	0	7770371_1	81.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7770371_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:64756658(-)-12:79558633(-)__12_79551501_79576501D;SPAN=14801975;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:42 GQ:18.5 PL:[81.2, 0.0, 18.5] SR:0 DR:28 LR:-83.03 LO:83.03);ALT=[chr12:79558633[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	80171338	+	chr12	64756660	+	TAGTTCTTTCATCCCCAA	0	68	7772158_1	99.0	.	EVDNC=ASSMB;INSERTION=TAGTTCTTTCATCCCCAA;MAPQ=60;MATEID=7772158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_80164001_80189001_146C;SPAN=15414678;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:53 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:68 DR:0 LR:-201.3 LO:201.3);ALT=]chr12:80171338]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	64761891	-	chr12	80917933	+	.	71	42	7665092_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=59;MATEID=7665092_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_64753501_64778501_392C;SPAN=16156042;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:93 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:42 DR:71 LR:-290.5 LO:290.5);ALT=[chr12:80917933[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	64944857	+	chr12	64939727	+	.	10	0	7666443_1	0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=7666443_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:64939727(-)-12:64944857(+)__12_64925001_64950001D;SPAN=5130;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:194 GQ:19.3 PL:[0.0, 19.3, 508.3] SR:0 DR:10 LR:19.55 LO:16.41);ALT=]chr12:64944857]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	66527651	+	chr12	66529877	+	.	164	75	7677203_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATGGTATTAATA;MAPQ=60;MATEID=7677203_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_66517501_66542501_375C;SPAN=2226;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:209 DP:51 GQ:56.5 PL:[620.5, 56.5, 0.0] SR:75 DR:164 LR:-620.6 LO:620.6);ALT=A[chr12:66529877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	67181819	-	chr12	67318749	+	.	57	14	7682363_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAA;MAPQ=60;MATEID=7682363_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_67301501_67326501_624C;SPAN=136930;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:131 GQ:99 PL:[189.2, 0.0, 126.5] SR:14 DR:57 LR:-189.6 LO:189.6);ALT=[chr12:67318749[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	68071678	+	chr14	100602967	+	CT	36	48	7690917_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CT;MAPQ=60;MATEID=7690917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_68061001_68086001_640C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:70 DP:163 GQ:99 PL:[187.1, 0.0, 206.9] SR:48 DR:36 LR:-186.9 LO:187.0);ALT=G[chr14:100602967[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	68072096	+	chr14	100603141	-	.	28	53	7690935_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7690935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_68061001_68086001_377C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:149 GQ:99 PL:[184.1, 0.0, 177.5] SR:53 DR:28 LR:-184.1 LO:184.1);ALT=G]chr14:100603141];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	79844324	+	chr12	77776071	+	.	62	53	7770800_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGTC;MAPQ=60;MATEID=7770800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_79821001_79846001_324C;SPAN=2068253;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:48 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:53 DR:62 LR:-274.0 LO:274.0);ALT=]chr12:79844324]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	78008285	+	chr12	79558904	+	.	16	38	7770373_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATTTT;MAPQ=60;MATEID=7770373_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_79551501_79576501_431C;SPAN=1550619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:38 DR:16 LR:-128.7 LO:128.7);ALT=T[chr12:79558904[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	79558905	+	chr12	78018015	+	.	15	68	7770374_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AAT;MAPQ=60;MATEID=7770374_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_79551501_79576501_306C;SPAN=1540890;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:44 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:68 DR:15 LR:-211.3 LO:211.3);ALT=]chr12:79558905]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	79607466	+	chr12	78019303	+	.	42	47	7770030_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGA;MAPQ=60;MATEID=7770030_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_79600501_79625501_180C;SPAN=1588163;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:49 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:47 DR:42 LR:-204.7 LO:204.7);ALT=]chr12:79607466]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	78019480	+	chr12	80917429	+	GGTG	22	26	7773262_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GGTG;MAPQ=60;MATEID=7773262_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_80899001_80924001_276C;SPAN=2897949;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:55 GQ:14.9 PL:[117.2, 0.0, 14.9] SR:26 DR:22 LR:-121.5 LO:121.5);ALT=G[chr12:80917429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	78019523	+	chr12	79559014	-	.	10	0	7770377_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7770377_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:78019523(+)-12:79559014(+)__12_79551501_79576501D;SPAN=1539491;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:0 DR:10 LR:-20.82 LO:23.18);ALT=C]chr12:79559014];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	79558496	+	chr12	78385564	+	.	39	0	7770378_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=7770378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:78385564(-)-12:79558496(+)__12_79551501_79576501D;SPAN=1172932;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:31 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:39 LR:-115.5 LO:115.5);ALT=]chr12:79558496]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	78385565	-	chr12	80171137	+	TACAAATTAATGCCATTGTGTCTGGAGCATATCATATAACTAATTATGCATGGCTTCTTAGAATGTTAGAAATTGTCACTTTGGGAGGCCGAGGTGAGCGGATCAAGAGGTCAGGAGTTTGAGACCATCTTGGCCAACATGGCGAAACACTGCCTCTACTAAAAATACAAAAAGTAGCCAGATGTGGTGGCGGG	25	54	7767407_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CACT;INSERTION=TACAAATTAATGCCATTGTGTCTGGAGCATATCATATAACTAATTATGCATGGCTTCTTAGAATGTTAGAAATTGTCACTTTGGGAGGCCGAGGTGAGCGGATCAAGAGGTCAGGAGTTTGAGACCATCTTGGCCAACATGGCGAAACACTGCCTCTACTAAAAATACAAAAAGTAGCCAGATGTGGTGGCGGG;MAPQ=60;MATEID=7767407_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_12_78375501_78400501_10C;SPAN=1785572;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:43 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:54 DR:25 LR:-184.8 LO:184.8);ALT=[chr12:80171137[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	79888360	+	chr12	79558153	+	ATCTTTAGAAACAATTACTTGAAG	44	36	7771532_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ATTT;INSERTION=ATCTTTAGAAACAATTACTTGAAG;MAPQ=60;MATEID=7771532_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TTT;SCTG=c_12_79870001_79895001_271C;SPAN=330207;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:33 GQ:18 PL:[198.0, 18.0, 0.0] SR:36 DR:44 LR:-198.0 LO:198.0);ALT=]chr12:79888360]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	79558454	+	chr12	80171219	-	ATCTTTAGAAACAATTACTTGAAG	17	40	7770390_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TTT;INSERTION=ATCTTTAGAAACAATTACTTGAAG;MAPQ=60;MATEID=7770390_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=TTT;SCTG=c_12_79551501_79576501_131C;SPAN=612765;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:32 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:40 DR:17 LR:-141.9 LO:141.9);ALT=T]chr12:80171219];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	79558634	-	chr12	80171214	+	.	31	30	7772162_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GTA;MAPQ=60;MATEID=7772162_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_80164001_80189001_115C;SPAN=612580;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:54 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:30 DR:31 LR:-158.4 LO:158.4);ALT=[chr12:80171214[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	79607507	+	chr12	80917418	+	.	12	0	7773264_1	25.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7773264_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:79607507(+)-12:80917418(-)__12_80899001_80924001D;SPAN=1309911;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=C[chr12:80917418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	79626495	-	chr12	79853781	+	TT	47	41	7770983_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TT;MAPQ=60;MATEID=7770983_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_12_79845501_79870501_6C;SPAN=227286;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:34 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:41 DR:47 LR:-234.4 LO:234.4);ALT=[chr12:79853781[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	79987561	+	chr12	81095100	-	.	34	0	7773918_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=7773918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:79987561(+)-12:81095100(+)__12_81070501_81095501D;SPAN=1107539;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:34 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:34 LR:-102.3 LO:102.3);ALT=C]chr12:81095100];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	90911081	+	chr12	115251922	+	.	8	44	7840672_1	99.0	.	DISC_MAPQ=11;EVDNC=ASDIS;HOMSEQ=CTTTCTTTCTTTCTTT;MAPQ=20;MATEID=7840672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_115248001_115273001_409C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:44 DP:28 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:44 DR:8 LR:-128.7 LO:128.7);ALT=]chr14:90911081]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	115681517	-	chr12	115716233	+	.	31	21	7841971_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CCCTC;MAPQ=60;MATEID=7841971_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_115713501_115738501_169C;SPAN=34716;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:70 GQ:27.2 PL:[142.7, 0.0, 27.2] SR:21 DR:31 LR:-147.2 LO:147.2);ALT=[chr12:115716233[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	115718807	+	chr16	6025564	+	.	61	42	7842002_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7842002_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_12_115713501_115738501_437C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:71 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:42 DR:61 LR:-250.9 LO:250.9);ALT=G[chr16:6025564[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	19570321	+	chr13	19568903	+	.	15	1	7929817_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGAAGG;MAPQ=60;MATEID=7929817_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_19551001_19576001_325C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:158 GQ:6.7 PL:[6.7, 0.0, 376.4] SR:1 DR:15 LR:-6.709 LO:28.73);ALT=]chr13:19570321]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	10953666	+	chr13	20050556	+	.	0	17	7931906_1	37.0	.	EVDNC=ASSMB;HOMSEQ=TACTGAAGCCTCC;MAPQ=56;MATEID=7931906_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_13_20041001_20066001_192C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:68 GQ:37.7 PL:[37.7, 0.0, 126.8] SR:17 DR:0 LR:-37.69 LO:40.42);ALT=]chr21:10953666]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr13	20825485	+	chr13	20828793	+	.	85	70	7936819_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGAT;MAPQ=60;MATEID=7936819_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_20800501_20825501_344C;SPAN=3308;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:50 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:70 DR:85 LR:-346.6 LO:346.6);ALT=T[chr13:20828793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49533337	+	chr13	49536619	+	.	28	0	8059052_1	72.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=8059052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:49533337(+)-13:49536619(-)__13_49514501_49539501D;SPAN=3282;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:74 GQ:72.5 PL:[72.5, 0.0, 105.5] SR:0 DR:28 LR:-72.38 LO:72.75);ALT=A[chr13:49536619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49951414	+	chr13	49953863	+	.	48	38	8060307_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAACAAAAACAGT;MAPQ=60;MATEID=8060307_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_49931001_49956001_206C;SPAN=2449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:76 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:38 DR:48 LR:-223.4 LO:223.4);ALT=T[chr13:49953863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	82859130	+	chr13	94778075	-	.	56	39	8233337_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8233337_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_94766001_94791001_421C;SPAN=11918945;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:73 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:39 DR:56 LR:-214.6 LO:214.6);ALT=T]chr13:94778075];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	83378291	-	chr13	94952534	+	AAAGAT	82	51	8234295_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AAAGAT;MAPQ=60;MATEID=8234295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_94937501_94962501_361C;SPAN=11574243;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:75 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:51 DR:82 LR:-307.0 LO:307.0);ALT=[chr13:94952534[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	83921691	+	chr13	83928158	+	CAACAACATTTAAG	0	39	8189103_1	99.0	.	EVDNC=ASSMB;INSERTION=CAACAACATTTAAG;MAPQ=60;MATEID=8189103_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_83912501_83937501_316C;SPAN=6467;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:84 GQ:96.2 PL:[106.1, 0.0, 96.2] SR:39 DR:0 LR:-106.0 LO:106.0);ALT=A[chr13:83928158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	95251182	+	chr13	95252198	-	.	10	0	8236368_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=8236368_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:95251182(+)-13:95252198(+)__13_95231501_95256501D;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:140 GQ:4.8 PL:[0.0, 4.8, 349.8] SR:0 DR:10 LR:4.919 LO:17.86);ALT=C]chr13:95252198];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	95783806	-	chr13	95785459	+	.	5	1	8239470_1	0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=CCCAG;MAPQ=44;MATEID=8239470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_95770501_95795501_455C;SPAN=1653;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:275 GQ:54.4 PL:[0.0, 54.4, 775.6] SR:1 DR:5 LR:54.7 LO:7.59);ALT=[chr13:95785459[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	96470642	+	chr13	96347414	+	.	85	39	8244915_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8244915_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_96456501_96481501_32C;SPAN=123228;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:125 GQ:30.3 PL:[363.0, 30.3, 0.0] SR:39 DR:85 LR:-362.9 LO:362.9);ALT=]chr13:96470642]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	96420954	+	chr13	96427829	+	.	81	49	8244020_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=8244020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_96407501_96432501_115C;SPAN=6875;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:101 DP:228 GQ:99 PL:[271.7, 0.0, 281.6] SR:49 DR:81 LR:-271.6 LO:271.6);ALT=C[chr13:96427829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	103443612	+	chr13	103451379	-	.	70	56	8289806_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGCC;MAPQ=60;MATEID=8289806_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_103439001_103464001_402C;SPAN=7767;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:135 GQ:9.9 PL:[346.5, 9.9, 0.0] SR:56 DR:70 LR:-359.6 LO:359.6);ALT=C]chr13:103451379];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	103443675	-	chr13	105854919	+	.	74	33	8298663_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=57;MATEID=8298663_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_105840001_105865001_390C;SPAN=2411244;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:78 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:33 DR:74 LR:-277.3 LO:277.3);ALT=[chr13:105854919[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	90328232	+	chr13	105798341	+	.	48	47	9060519_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=9060519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90307001_90332001_328C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:84 GQ:6 PL:[214.5, 6.0, 0.0] SR:47 DR:48 LR:-222.4 LO:222.4);ALT=]chr15:90328232]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr13	105798356	+	chr15	90328126	+	TTTTTTTTTTTTTTTTTT	45	63	8298603_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=TTTATTAAATTTTTTTT;INSERTION=TTTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=8298603_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_105791001_105816001_180C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:51 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:63 DR:45 LR:-250.9 LO:250.9);ALT=T[chr15:90328126[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr14	45769273	-	chr14	45837612	+	ATC	56	49	8477534_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ATC;MAPQ=60;MATEID=8477534_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_45766001_45791001_8C;SPAN=68339;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:64 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:49 DR:56 LR:-270.7 LO:270.7);ALT=[chr14:45837612[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	45770427	+	chr14	61463062	+	.	74	19	8540779_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTA;MAPQ=60;MATEID=8540779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_61446001_61471001_110C;SPAN=15692635;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:65 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:19 DR:74 LR:-254.2 LO:254.2);ALT=A[chr14:61463062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45775965	+	chr14	61465413	+	.	85	50	8540780_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=8540780_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_61446001_61471001_14C;SPAN=15689448;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:114 DP:125 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:50 DR:85 LR:-369.7 LO:369.7);ALT=G[chr14:61465413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45776151	-	chr14	47703224	+	.	47	43	8481656_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=8481656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_47701501_47726501_364C;SPAN=1927073;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:63 GQ:21 PL:[231.0, 21.0, 0.0] SR:43 DR:47 LR:-231.1 LO:231.1);ALT=[chr14:47703224[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	45801498	+	chr14	47703726	-	.	47	44	8481658_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=8481658_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_47701501_47726501_158C;SPAN=1902228;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:58 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:44 DR:47 LR:-247.6 LO:247.6);ALT=T]chr14:47703726];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	45855301	+	chr14	47640078	+	.	0	44	8481319_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AAGTTAA;MAPQ=60;MATEID=8481319_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_47628001_47653001_11C;SPAN=1784777;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:44 DP:28 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:44 DR:0 LR:-128.7 LO:128.7);ALT=A[chr14:47640078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	61184792	+	chr14	46283809	+	.	45	12	8539050_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=8539050_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_61176501_61201501_222C;SPAN=14900983;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:61 GQ:3 PL:[151.8, 3.0, 0.0] SR:12 DR:45 LR:-157.9 LO:157.9);ALT=]chr14:61184792]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	46646784	+	chr14	61465762	-	.	60	23	8479735_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=8479735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_46623501_46648501_263C;SPAN=14818978;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:26 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:23 DR:60 LR:-234.4 LO:234.4);ALT=T]chr14:61465762];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	47117868	-	chr14	63226284	+	.	31	40	8551095_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;MAPQ=0;MATEID=8551095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_63210001_63235001_511C;SPAN=16108416;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:54 GQ:18 PL:[198.0, 18.0, 0.0] SR:40 DR:31 LR:-198.0 LO:198.0);ALT=[chr14:63226284[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	48323968	-	chr14	48325262	+	.	42	55	8483579_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8483579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_48314001_48339001_400C;SPAN=1294;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:81 DP:113 GQ:35.6 PL:[236.9, 0.0, 35.6] SR:55 DR:42 LR:-245.1 LO:245.1);ALT=[chr14:48325262[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	55491318	+	chr22	18934743	+	.	9	0	10838800_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10838800_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55491318(+)-22:18934743(-)__22_18914001_18939001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:0 DR:9 LR:-4.784 LO:17.36);ALT=A[chr22:18934743[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr14	55904996	-	chr14	55906449	+	.	10	0	8516884_1	2.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=8516884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55904996(-)-14:55906449(-)__14_55884501_55909501D;SPAN=1453;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:115 GQ:2 PL:[2.0, 0.0, 275.9] SR:0 DR:10 LR:-1.854 LO:18.75);ALT=[chr14:55906449[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	55931135	+	chrX	48531139	-	.	13	0	11150232_1	33.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=11150232_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55931135(+)-23:48531139(+)__23_48510001_48535001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:36 GQ:33.2 PL:[33.2, 0.0, 53.0] SR:0 DR:13 LR:-33.16 LO:33.44);ALT=T]chrX:48531139];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr20	32337222	+	chr14	57466339	+	CAGTAGCTGGGATTACAAATGCCTGCCACCATGCCCAGGTAATTTAGAGACTGGGTTTCACCACGTTAGCCAGGC	6	58	8523660_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TGGTCTTGAACTCC;INSERTION=CAGTAGCTGGGATTACAAATGCCTGCCACCATGCCCAGGTAATTTAGAGACTGGGTTTCACCACGTTAGCCAGGC;MAPQ=60;MATEID=8523660_2;MATENM=3;NM=0;NUMPARTS=4;SCTG=c_14_57452501_57477501_344C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:64 DP:43 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:58 DR:6 LR:-188.1 LO:188.1);ALT=]chr20:32337222]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr14	58259348	-	chr14	58412167	+	.	29	0	8527927_1	85.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=8527927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58259348(-)-14:58412167(-)__14_58408001_58433001D;SPAN=152819;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:19 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=[chr14:58412167[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	60341398	+	chr14	60343242	+	.	133	117	8535183_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8535183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_60319001_60344001_286C;SPAN=1844;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:196 DP:40 GQ:52.9 PL:[580.9, 52.9, 0.0] SR:117 DR:133 LR:-580.9 LO:580.9);ALT=T[chr14:60343242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	62341344	+	chr14	60702364	+	.	78	50	8546452_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=8546452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_62328001_62353001_134C;SPAN=1638980;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:102 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:50 DR:78 LR:-323.5 LO:323.5);ALT=]chr14:62341344]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	73600315	+	chr14	73515049	+	.	65	30	8597299_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=52;MATEID=8597299_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73598001_73623001_414C;SPAN=85266;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:83 DP:104 GQ:5 PL:[245.9, 0.0, 5.0] SR:30 DR:65 LR:-259.6 LO:259.6);ALT=]chr14:73600315]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	74594794	+	chr14	73710471	+	.	66	38	8605749_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=8605749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74578001_74603001_198C;SPAN=884323;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:92 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:38 DR:66 LR:-270.7 LO:270.7);ALT=]chr14:74594794]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	74239795	+	chr14	74246937	+	.	134	147	8602247_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=8602247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74235001_74260001_199C;SPAN=7142;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:218 DP:130 GQ:58.9 PL:[646.9, 58.9, 0.0] SR:147 DR:134 LR:-647.0 LO:647.0);ALT=C[chr14:74246937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74534936	+	chr14	74535985	-	.	0	4	8605140_1	0	.	EVDNC=ASSMB;HOMSEQ=AAAATACAAAAATTAG;MAPQ=60;MATEID=8605140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74529001_74554001_4C;SPAN=1049;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:186 GQ:37 PL:[0.0, 37.0, 524.8] SR:4 DR:0 LR:37.19 LO:5.035);ALT=G]chr14:74535985];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	74559374	+	chr14	74561226	+	.	87	55	8605574_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=8605574_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74553501_74578501_49C;SPAN=1852;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:115 DP:157 GQ:43.4 PL:[337.1, 0.0, 43.4] SR:55 DR:87 LR:-350.1 LO:350.1);ALT=C[chr14:74561226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74667010	-	chr19	33417587	+	.	8	0	8606229_1	6.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=8606229_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:74667010(-)-19:33417587(-)__14_74651501_74676501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:0 DR:8 LR:-6.089 LO:15.75);ALT=[chr19:33417587[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	96172397	-	chr21	36792263	+	.	7	64	10770981_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=AGATAGATAGACAGACAGACAGATAGA;MAPQ=34;MATEID=10770981_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_21_36774501_36799501_64C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:46 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:64 DR:7 LR:-191.4 LO:191.4);ALT=[chr21:36792263[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr15	20022131	+	chr15	20024080	+	.	71	0	8747859_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=8747859_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:20022131(+)-15:20024080(-)__15_20016501_20041501D;SPAN=1949;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:10 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=T[chr15:20024080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	33628756	-	chr20	23541588	+	.	13	57	8838075_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=8838075_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_15_33614001_33639001_10C;SECONDARY;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:27 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:57 DR:13 LR:-204.7 LO:204.7);ALT=[chr20:23541588[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr15	42962505	+	chr15	42759006	+	.	11	10	8876105_1	38.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=8876105_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42948501_42973501_354C;SPAN=203499;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:43 GQ:38 PL:[38.0, 0.0, 64.4] SR:10 DR:11 LR:-37.87 LO:38.3);ALT=]chr15:42962505]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	43368155	-	chr20	5268410	+	AGAGGGC	16	44	8877399_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;INSERTION=AGAGGGC;MAPQ=15;MATEID=8877399_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_15_43365001_43390001_241C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:57 DP:40 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:44 DR:16 LR:-168.3 LO:168.3);ALT=[chr20:5268410[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr15	51864402	+	chr15	51801632	+	.	11	0	8896018_1	30.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=8896018_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:51801632(-)-15:51864402(+)__15_51842001_51867001D;SPAN=62770;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:21 GQ:17.6 PL:[30.8, 0.0, 17.6] SR:0 DR:11 LR:-30.73 LO:30.73);ALT=]chr15:51864402]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	51801761	+	chr15	51864510	+	.	19	0	8896019_1	52.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=8896019_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:51801761(+)-15:51864510(-)__15_51842001_51867001D;SPAN=62749;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:37 GQ:36.2 PL:[52.7, 0.0, 36.2] SR:0 DR:19 LR:-52.84 LO:52.84);ALT=A[chr15:51864510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55655547	+	chr15	55657029	+	.	86	31	8904185_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTGGGCAACAGAGCGAGGCTCCATCTCA;MAPQ=60;MATEID=8904185_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_55639501_55664501_163C;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:22 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:31 DR:86 LR:-326.8 LO:326.8);ALT=A[chr15:55657029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	68461178	+	chr15	56251135	+	.	6	25	9789700_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=9789700_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_68453001_68478001_83C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:121 GQ:69.8 PL:[69.8, 0.0, 221.6] SR:25 DR:6 LR:-69.55 LO:74.09);ALT=]chr17:68461178]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr15	81360254	+	chr20	34272339	-	CATAACATAACAAAC	6	22	9017014_1	68.0	.	DISC_MAPQ=4;EVDNC=ASDIS;INSERTION=CATAACATAACAAAC;MAPQ=16;MATEID=9017014_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_81340001_81365001_1C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:77 GQ:68.3 PL:[68.3, 0.0, 117.8] SR:22 DR:6 LR:-68.27 LO:69.01);ALT=T]chr20:34272339];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr21	27196911	+	chr16	5285837	+	.	10	8	9127770_1	47.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTTTT;MAPQ=23;MATEID=9127770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_5267501_5292501_94C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:30 GQ:24.8 PL:[47.9, 0.0, 24.8] SR:8 DR:10 LR:-48.39 LO:48.39);ALT=]chr21:27196911]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	5949478	+	chr16	7349172	+	.	55	53	9129648_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=9129648_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_16_7325501_7350501_8C;SPAN=1399694;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:42 GQ:24 PL:[264.0, 24.0, 0.0] SR:53 DR:55 LR:-264.1 LO:264.1);ALT=G[chr16:7349172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	6075881	+	chr16	6099307	+	.	55	51	9129414_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=9129414_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_16_6051501_6076501_5C;SPAN=23426;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:8 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:51 DR:55 LR:-270.7 LO:270.7);ALT=A[chr16:6099307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	6101608	+	chr16	6138466	+	ACTTT	91	77	9129353_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=ACTTT;MAPQ=60;MATEID=9129353_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_6125001_6150001_49C;SPAN=36858;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:137 DP:17 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:77 DR:91 LR:-406.0 LO:406.0);ALT=C[chr16:6138466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	6153889	+	chr16	6509091	+	GGAAATTCC	89	52	9129422_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GGAAATTCC;MAPQ=60;MATEID=9129422_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_6492501_6517501_43C;SPAN=355202;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:12 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:52 DR:89 LR:-316.9 LO:316.9);ALT=T[chr16:6509091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	6535234	+	chr16	7155803	-	ACCCTTTCCCCTGAGTCCACAAAGTCCATTGTGTCATTCTTATGCCTTTGCTTCCTCATAGCTTAGCTCCCACTTACGAGTGAGAACATACAACGTTTGGTTTTGCATTCCTGAGTTAGTCTGCAATCTCATCCAGGTTGCTGCGAATGCCATTGACCCATTCCTTTTTATGGCTGAGTCATATTCCATCATA	5	82	9129570_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TTGTGTCATTCTTATGCCTTTGCTTCCTCATAGCTTAGCTCCCACTTACGAGTGAGAACATACAACGTTTGGTTTTGCATTCCTGAGTTAGTCTGCAATCTCATCCAGGTTGCTGCGAATGCCATTGACCCATTCCTTTTTATGGCTGAGTCATATTCCATCATATCTATCT;INSERTION=ACCCTTTCCCCTGAGTCCACAAAGTCCATTGTGTCATTCTTATGCCTTTGCTTCCTCATAGCTTAGCTCCCACTTACGAGTGAGAACATACAACGTTTGGTTTTGCATTCCTGAGTTAGTCTGCAATCTCATCCAGGTTGCTGCGAATGCCATTGACCCATTCCTTTTTATGGCTGAGTCATATTCCATCATA;MAPQ=60;MATEID=9129570_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_16_7154001_7179001_160C;SECONDARY;SPAN=620569;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:28 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:82 DR:5 LR:-250.9 LO:250.9);ALT=C]chr16:7155803];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	6535234	+	chr16	7155480	+	.	94	57	9129569_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CTTCC;MAPQ=60;MATEID=9129569_2;MATENM=0;NM=2;NUMPARTS=3;REPSEQ=CCC;SCTG=c_16_7154001_7179001_160C;SPAN=620246;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:132 DP:14 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:57 DR:94 LR:-389.5 LO:389.5);ALT=C[chr16:7155480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	7172400	+	chr16	7233555	+	.	55	43	9129610_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTG;MAPQ=60;MATEID=9129610_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_7154001_7179001_6C;SPAN=61155;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:6 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:43 DR:55 LR:-237.7 LO:237.7);ALT=G[chr16:7233555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78325356	+	chr16	78339513	+	.	47	36	9431922_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=9431922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_78326501_78351501_89C;SPAN=14157;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:11 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:36 DR:47 LR:-204.7 LO:204.7);ALT=T[chr16:78339513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78615516	+	chr16	78736814	+	.	81	49	9432355_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=9432355_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_78596001_78621001_89C;SPAN=121298;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:9 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:49 DR:81 LR:-280.6 LO:280.6);ALT=A[chr16:78736814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78745811	+	chr16	78784787	+	.	74	50	9432322_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=9432322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_78767501_78792501_86C;SPAN=38976;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:12 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:50 DR:74 LR:-303.7 LO:303.7);ALT=C[chr16:78784787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78885452	+	chr16	78899365	+	.	0	33	9432627_1	95.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=9432627_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_78890001_78915001_169C;SPAN=13913;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:33 DP:21 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:33 DR:0 LR:-95.72 LO:95.72);ALT=A[chr16:78899365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	79499072	+	chr16	78925426	+	.	45	39	9434790_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=9434790_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_79478001_79503001_95C;SPAN=573646;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:36 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:45 LR:-201.3 LO:201.3);ALT=]chr16:79499072]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	79205904	+	chr16	79197893	+	.	131	83	9433634_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=9433634_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_79184001_79209001_145C;SPAN=8011;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:163 DP:146 GQ:43.9 PL:[481.9, 43.9, 0.0] SR:83 DR:131 LR:-481.9 LO:481.9);ALT=]chr16:79205904]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	79242908	+	chr16	79218751	+	TGTCTTT	81	41	9434161_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TGTCTTT;MAPQ=60;MATEID=9434161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_79233001_79258001_161C;SPAN=24157;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:112 DP:86 GQ:30 PL:[330.0, 30.0, 0.0] SR:41 DR:81 LR:-330.1 LO:330.1);ALT=]chr16:79242908]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	25536553	+	chr17	25540382	+	.	173	89	9571269_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAATTCACATGGCA;MAPQ=60;MATEID=9571269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25529001_25554001_196C;SPAN=3829;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:220 DP:59 GQ:59.5 PL:[653.5, 59.5, 0.0] SR:89 DR:173 LR:-653.6 LO:653.6);ALT=A[chr17:25540382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26356915	-	chr17	26358570	+	.	9	0	9574952_1	1.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=9574952_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:26356915(-)-17:26358570(-)__17_26337501_26362501D;SPAN=1655;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:0 DR:9 LR:-1.262 LO:16.82);ALT=[chr17:26358570[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	27126542	-	chr17	27127913	+	.	14	0	9578538_1	10.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=9578538_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:27126542(-)-17:27127913(-)__17_27121501_27146501D;SPAN=1371;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:134 GQ:10.1 PL:[10.1, 0.0, 313.7] SR:0 DR:14 LR:-9.91 LO:27.43);ALT=[chr17:27127913[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	122597535	+	chr17	33857509	+	.	8	0	9611645_1	18.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=9611645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:33857509(-)-23:122597535(+)__17_33834501_33859501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:0 DR:8 LR:-18.55 LO:19.42);ALT=]chrX:122597535]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	68455097	+	chr17	68461177	+	.	108	57	9789703_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAGATTTTGTG;MAPQ=60;MATEID=9789703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_68453001_68478001_236C;SPAN=6080;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:139 DP:154 GQ:41.5 PL:[455.5, 41.5, 0.0] SR:57 DR:108 LR:-455.5 LO:455.5);ALT=G[chr17:68461177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39044999	+	chr17	80313286	+	GAGAATCATTTGAACCTGGGAGGTAGAGGTTGCA	26	94	10288321_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_G;HOMSEQ=GTGAGCTGAGATCGCGCCATTGCACTCCA;INSERTION=GAGAATCATTTGAACCTGGGAGGTAGAGGTTGCA;MAPQ=33;MATEID=10288321_2;MATENM=2;NM=2;NUMPARTS=3;SCTG=c_19_39028501_39053501_618C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:63 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:94 DR:26 LR:-303.7 LO:303.7);ALT=]chr19:39044999]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr18	33144440	+	chr18	32973131	+	GA	7	7	9979931_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GA;MAPQ=60;MATEID=9979931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_33124001_33149001_437C;SPAN=171309;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:7 DR:7 LR:-16.31 LO:25.12);ALT=]chr18:33144440]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr18	38064076	+	chr18	67448633	+	.	47	42	10051490_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10051490_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_67448501_67473501_95C;SPAN=29384557;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:45 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:42 DR:47 LR:-201.3 LO:201.3);ALT=A[chr18:67448633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	38259893	+	chr18	38266750	+	.	58	51	9998762_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=9998762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_38244501_38269501_59C;SPAN=6857;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:19 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:51 DR:58 LR:-260.8 LO:260.8);ALT=T[chr18:38266750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	38864779	+	chr18	38868344	+	TAAAACTCTTTTAAG	0	30	9999866_1	89.0	.	EVDNC=ASSMB;INSERTION=TAAAACTCTTTTAAG;MAPQ=60;MATEID=9999866_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_38857001_38882001_211C;SPAN=3565;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:30 DP:17 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:30 DR:0 LR:-89.12 LO:89.12);ALT=T[chr18:38868344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	39819980	+	chr18	39754276	+	CA	88	50	10001331_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CA;MAPQ=60;MATEID=10001331_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_39812501_39837501_33C;SPAN=65704;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:42 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:50 DR:88 LR:-346.6 LO:346.6);ALT=]chr18:39819980]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr18	42707914	+	chr20	43033460	-	.	55	0	10560473_1	95.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=10560473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:42707914(+)-20:43033460(+)__20_43022001_43047001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:318 GQ:95.5 PL:[95.5, 0.0, 676.4] SR:0 DR:55 LR:-95.4 LO:120.8);ALT=G]chr20:43033460];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr18	68383825	+	chr18	68405444	+	.	14	0	10056313_1	17.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=10056313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:68383825(+)-18:68405444(-)__18_68404001_68429001D;SPAN=21619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:105 GQ:17.9 PL:[17.9, 0.0, 235.7] SR:0 DR:14 LR:-17.77 LO:29.01);ALT=A[chr18:68405444[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	68405855	+	chr18	68387238	+	.	53	0	10056314_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=10056314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:68387238(-)-18:68405855(+)__18_68404001_68429001D;SPAN=18617;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:62 GQ:9.9 PL:[168.3, 9.9, 0.0] SR:0 DR:53 LR:-170.1 LO:170.1);ALT=]chr18:68405855]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr18	68405811	+	chr18	68408815	+	TATTCACGATAGCAAAGACTTGCAAC	0	56	10056325_1	99.0	.	EVDNC=ASSMB;INSERTION=TATTCACGATAGCAAAGACTTGCAAC;MAPQ=60;MATEID=10056325_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_18_68404001_68429001_207C;SPAN=3004;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:154 GQ:99 PL:[143.3, 0.0, 229.1] SR:56 DR:0 LR:-143.1 LO:144.3);ALT=T[chr18:68408815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	20095911	-	chrX	29350711	+	.	23	0	11046645_1	58.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=11046645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:20095911(-)-23:29350711(-)__23_29326501_29351501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:65 GQ:58.4 PL:[58.4, 0.0, 98.0] SR:0 DR:23 LR:-58.31 LO:58.9);ALT=[chrX:29350711[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr19	20771460	+	chr19	20924894	-	.	9	0	10212359_1	9.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=10212359_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:20771460(+)-19:20924894(+)__19_20923001_20948001D;SPAN=153434;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:0 DR:9 LR:-9.119 LO:18.15);ALT=G]chr19:20924894];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	20802049	-	chr19	20883039	+	.	86	0	10211600_1	99.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=10211600_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:20802049(-)-19:20883039(-)__19_20874001_20899001D;SPAN=80990;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:98 GQ:19.8 PL:[277.2, 19.8, 0.0] SR:0 DR:86 LR:-279.4 LO:279.4);ALT=[chr19:20883039[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	21268380	+	chr19	21328014	+	.	8	0	10213770_1	6.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=10213770_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:21268380(+)-19:21328014(-)__19_21315001_21340001D;SPAN=59634;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=A[chr19:21328014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21334763	+	chr19	21272695	+	.	33	13	10213930_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGAAATTTGTACACTTTTGCCAGCATGCCAGGCTTCTGGG;MAPQ=60;MATEID=10213930_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_21266001_21291001_456C;SPAN=62068;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:35 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:13 DR:33 LR:-115.5 LO:115.5);ALT=]chr19:21334763]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	21336431	+	chr19	21274430	+	.	10	0	10213935_1	18.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=10213935_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:21274430(-)-19:21336431(+)__19_21266001_21291001D;SPAN=62001;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:54 GQ:18.5 PL:[18.5, 0.0, 110.9] SR:0 DR:10 LR:-18.38 LO:22.29);ALT=]chr19:21336431]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	33663511	+	chr19	33567307	+	.	13	0	10257931_1	26.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=10257931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:33567307(-)-19:33663511(+)__19_33638501_33663501D;SPAN=96204;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:61 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.39 LO:29.87);ALT=]chr19:33663511]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	33663725	+	chr19	33567308	+	.	13	7	10258162_1	29.0	.	DISC_MAPQ=48;EVDNC=ASDIS;MAPQ=30;MATEID=10258162_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_33663001_33688001_360C;SPAN=96417;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:62 GQ:29.6 PL:[29.6, 0.0, 118.7] SR:7 DR:13 LR:-29.42 LO:32.57);ALT=]chr19:33663725]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	33862170	-	chr19	33863742	+	.	10	0	10258604_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10258604_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:33862170(-)-19:33863742(-)__19_33859001_33884001D;SPAN=1572;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:109 GQ:3.5 PL:[3.5, 0.0, 260.9] SR:0 DR:10 LR:-3.479 LO:19.0);ALT=[chr19:33863742[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	35661081	+	chr19	35665798	+	.	92	43	10268051_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=0;MATEID=10268051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_35647501_35672501_362C;SECONDARY;SPAN=4717;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:101 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:43 DR:92 LR:-316.9 LO:316.9);ALT=C[chr19:35665798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36488006	-	chr19	36489104	+	.	8	0	10271285_1	0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=10271285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36488006(-)-19:36489104(-)__19_36480501_36505501D;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:140 GQ:11.4 PL:[0.0, 11.4, 363.0] SR:0 DR:8 LR:11.52 LO:13.49);ALT=[chr19:36489104[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	122804408	+	chr19	39044978	+	.	13	0	10288410_1	23.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=10288410_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39044978(-)-23:122804408(+)__19_39028501_39053501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:71 GQ:23.9 PL:[23.9, 0.0, 146.0] SR:0 DR:13 LR:-23.68 LO:28.9);ALT=]chrX:122804408]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr20	2803162	+	chr20	2806410	+	.	62	37	10401841_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAGAACTTGATTT;MAPQ=60;MATEID=10401841_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2793001_2818001_80C;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:32 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:37 DR:62 LR:-244.3 LO:244.3);ALT=T[chr20:2806410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	4021215	-	chr20	10505041	+	.	66	23	10421380_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=10421380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_10486001_10511001_133C;SPAN=6483826;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:43 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:23 DR:66 LR:-237.7 LO:237.7);ALT=[chr20:10505041[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	4071034	+	chr20	5546460	-	.	79	25	10412349_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10412349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_5537001_5562001_129C;SPAN=1475426;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:32 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:25 DR:79 LR:-267.4 LO:267.4);ALT=T]chr20:5546460];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	5599463	+	chr20	5600678	-	.	9	0	10412444_1	16.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=10412444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:5599463(+)-20:5600678(+)__20_5586001_5611001D;SPAN=1215;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=C]chr20:5600678];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	5906787	+	chr21	38018084	+	GTATG	9	14	10776615_1	24.0	.	DISC_MAPQ=0;EVDNC=TSI_L;HOMSEQ=AGAGAGAGAGAGAGAGAGA;INSERTION=GTATG;MAPQ=60;MATEID=10776615_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=AGAGAGAGAGAGAGAGAG;SCTG=c_21_37999501_38024501_273C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:20 DP:18 GQ:5 PL:[24.8, 5.0, 0.0] SR:14 DR:9 LR:-24.84 LO:24.84);ALT=A[chr21:38018084[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	11281584	-	chrX	81651235	+	AGTATTAAA	27	42	10424437_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AGTATTAAA;MAPQ=60;MATEID=10424437_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_20_11270001_11295001_120C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:39 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:42 DR:27 LR:-178.2 LO:178.2);ALT=[chrX:81651235[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr20	12436601	+	chr20	12180501	+	.	72	20	10429443_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTG;MAPQ=60;MATEID=10429443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_12421501_12446501_312C;SPAN=256100;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:35 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:20 DR:72 LR:-237.7 LO:237.7);ALT=]chr20:12436601]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	22151117	+	chr20	12338511	+	.	13	0	10429350_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=10429350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:12338511(-)-20:22151117(+)__20_12323501_12348501D;SPAN=9812606;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:48 GQ:29.9 PL:[29.9, 0.0, 86.0] SR:0 DR:13 LR:-29.91 LO:31.44);ALT=]chr20:22151117]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	12452382	+	chr20	12338512	+	ATATTATTTACCATTCTTCTGTAACCTCCTATTCCCTCAGCATAAAATCTACACTTTTGAAGGTACTGCATAACACCATTTGGTTCACTCAGCACTGGGCTTACAC	19	88	10429352_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=GCTC;INSERTION=ATATTATTTACCATTCTTCTGTAACCTCCTATTCCCTCAGCATAAAATCTACACTTTTGAAGGTACTGCATAACACCATTTGGTTCACTCAGCACTGGGCTTACAC;MAPQ=60;MATEID=10429352_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_12323501_12348501_51C;SPAN=113870;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:50 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:88 DR:19 LR:-300.4 LO:300.4);ALT=]chr20:12452382]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	12338512	-	chr20	12451965	+	.	26	56	10429351_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GCTC;MAPQ=60;MATEID=10429351_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TATTAT;SCTG=c_20_12323501_12348501_51C;SPAN=113453;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:50 GQ:18.8 PL:[163.8, 18.8, 0.0] SR:56 DR:26 LR:-163.9 LO:163.9);ALT=[chr20:12451965[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	12451770	-	chr20	22143554	+	ACTGTAT	40	38	10446557_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GATT;INSERTION=ACTGTAT;MAPQ=60;MATEID=10446557_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_20_22123501_22148501_34C;SPAN=9691784;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:47 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:38 DR:40 LR:-211.3 LO:211.3);ALT=[chr20:22143554[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	12451959	+	chr20	22150844	+	.	25	19	10446868_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AATTTA;MAPQ=60;MATEID=10446868_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_20_22148001_22173001_425C;SPAN=9698885;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:42 DP:61 GQ:23.3 PL:[122.3, 0.0, 23.3] SR:19 DR:25 LR:-125.6 LO:125.6);ALT=A[chr20:22150844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	22151064	+	chr20	12452247	+	ATACAGT	20	43	10428942_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AATTTA;INSERTION=ATACAGT;MAPQ=60;MATEID=10428942_2;MATENM=1;NM=0;NUMPARTS=4;SCTG=c_20_12446001_12471001_261C;SPAN=9698817;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:45 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:43 DR:20 LR:-155.1 LO:155.1);ALT=]chr20:22151064]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	14559862	+	chr20	14596956	-	.	56	0	10433442_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=10433442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:14559862(+)-20:14596956(+)__20_14577501_14602501D;SPAN=37094;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:56 DP:0 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:56 LR:-165.0 LO:165.0);ALT=A]chr20:14596956];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	14559994	-	chr20	14677065	+	CACC	60	39	10433192_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=CACC;MAPQ=0;MATEID=10433192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_14553001_14578001_66C;SECONDARY;SPAN=117071;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:24 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:39 DR:60 LR:-274.0 LO:274.0);ALT=[chr20:14677065[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	14732422	+	chr20	14869025	+	.	83	70	10433124_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGTC;MAPQ=60;MATEID=10433124_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_14847001_14872001_0C;SPAN=136603;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:119 DP:13 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:70 DR:83 LR:-353.2 LO:353.2);ALT=C[chr20:14869025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	15016452	+	chr20	15126125	+	.	59	51	10433566_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAT;MAPQ=60;MATEID=10433566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_15116501_15141501_159C;SPAN=109673;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:9 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:51 DR:59 LR:-257.5 LO:257.5);ALT=T[chr20:15126125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16079002	+	chr20	16085370	+	CATGCATATAATTGACTA	0	59	10435030_1	99.0	.	EVDNC=ASSMB;INSERTION=CATGCATATAATTGACTA;MAPQ=60;MATEID=10435030_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_16072001_16097001_138C;SPAN=6368;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:21 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:59 DR:0 LR:-174.9 LO:174.9);ALT=G[chr20:16085370[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16239637	+	chr20	16238391	+	.	9	0	10435504_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=10435504_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:16238391(-)-20:16239637(+)__20_16219001_16244001D;SPAN=1246;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:122 GQ:3 PL:[0.0, 3.0, 300.3] SR:0 DR:9 LR:3.344 LO:16.21);ALT=]chr20:16239637]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	21286134	+	chr20	21288751	+	.	60	0	10445197_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=10445197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:21286134(+)-20:21288751(-)__20_21266001_21291001D;SPAN=2617;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:8 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=C[chr20:21288751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	22143553	-	chr20	22150835	+	.	16	0	10446871_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10446871_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:22143553(-)-20:22150835(-)__20_22148001_22173001D;SPAN=7282;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:53 GQ:38.6 PL:[38.6, 0.0, 88.1] SR:0 DR:16 LR:-38.46 LO:39.6);ALT=[chr20:22150835[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	23963022	+	chr22	24642332	+	.	9	0	10455526_1	18.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=10455526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:23963022(+)-22:24642332(-)__20_23961001_23986001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:43 GQ:18.2 PL:[18.2, 0.0, 84.2] SR:0 DR:9 LR:-18.06 LO:20.6);ALT=A[chr22:24642332[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	32815938	+	chr20	32819226	+	.	111	67	10490839_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAGAACTTTC;MAPQ=60;MATEID=10490839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32805501_32830501_355C;SPAN=3288;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:162 DP:697 GQ:99 PL:[346.1, 0.0, 1346.0] SR:67 DR:111 LR:-345.9 LO:379.2);ALT=C[chr20:32819226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42024612	+	chr20	42025793	+	.	61	38	10553253_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGGTAAAACCCCATTTCT;MAPQ=60;MATEID=10553253_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_42017501_42042501_116C;SPAN=1181;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:79 DP:122 GQ:66.2 PL:[227.9, 0.0, 66.2] SR:38 DR:61 LR:-232.5 LO:232.5);ALT=T[chr20:42025793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42271923	+	chr20	42274577	+	.	84	0	10555285_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=10555285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:42271923(+)-20:42274577(-)__20_42262501_42287501D;SPAN=2654;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:103 GQ:1.2 PL:[250.8, 1.2, 0.0] SR:0 DR:84 LR:-264.7 LO:264.7);ALT=T[chr20:42274577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43033706	+	chr20	43030775	+	.	8	0	10560526_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10560526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:43030775(-)-20:43033706(+)__20_43022001_43047001D;SPAN=2931;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:625 GQ:99 PL:[0.0, 142.6, 1802.0] SR:0 DR:8 LR:142.9 LO:8.299);ALT=]chr20:43033706]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	43305847	+	chr20	43312215	-	.	111	109	10562662_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=10562662_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_43291501_43316501_589C;SPAN=6368;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:192 DP:175 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:109 DR:111 LR:-567.7 LO:567.7);ALT=T]chr20:43312215];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	55224961	-	chr20	55228175	+	.	8	0	10641244_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=10641244_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:55224961(-)-20:55228175(-)__20_55223001_55248001D;SPAN=3214;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:163 GQ:17.5 PL:[0.0, 17.5, 429.1] SR:0 DR:8 LR:17.75 LO:12.95);ALT=[chr20:55228175[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	23852644	+	chr20	55239234	+	.	15	79	10853097_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10853097_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_22_23838501_23863501_260C;SECONDARY;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:33 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:79 DR:15 LR:-237.7 LO:237.7);ALT=]chr22:23852644]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr21	37511992	-	chr21	37513242	+	.	11	0	10774303_1	4.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=10774303_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:37511992(-)-21:37513242(-)__21_37509501_37534501D;SPAN=1250;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:117 GQ:4.7 PL:[4.7, 0.0, 278.6] SR:0 DR:11 LR:-4.613 LO:21.02);ALT=[chr21:37513242[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	18057770	+	chr22	18060458	+	.	107	74	10834459_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=ATTCTCCTGCCTCAGCCTCC;MAPQ=60;MATEID=10834459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18056501_18081501_87C;SPAN=2688;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:165 DP:47 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:74 DR:107 LR:-488.5 LO:488.5);ALT=C[chr22:18060458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24195941	+	chr22	24198506	+	.	50	47	10854072_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=GAAAAAAA;MAPQ=60;MATEID=10854072_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_22_24181501_24206501_209C;SPAN=2565;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:30 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:47 DR:50 LR:-234.4 LO:234.4);ALT=A[chr22:24198506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24276436	+	chr22	24279226	+	.	59	47	10854199_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CG;MAPQ=60;MATEID=10854199_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_22_24279501_24304501_18C;SPAN=2790;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:0 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:47 DR:59 LR:-267.4 LO:267.4);ALT=G[chr22:24279226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	4724929	+	chrX	4726799	+	.	13	11	10942620_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=10942620_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_4704001_4729001_326C;SPAN=1870;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:136 GQ:22.7 PL:[22.7, 0.0, 306.5] SR:11 DR:13 LR:-22.57 LO:37.24);ALT=T[chrX:4726799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	5055347	+	chrX	5057500	+	.	115	112	10943938_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTTA;MAPQ=60;MATEID=10943938_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_5047001_5072001_334C;SPAN=2153;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:183 DP:38 GQ:49.3 PL:[541.3, 49.3, 0.0] SR:112 DR:115 LR:-541.3 LO:541.3);ALT=A[chrX:5057500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	5729125	-	chrX	5730607	+	.	80	93	10946926_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCCAC;MAPQ=60;MATEID=10946926_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_5708501_5733501_88C;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:160 DP:125 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:93 DR:80 LR:-475.3 LO:475.3);ALT=[chrX:5730607[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	5729126	+	chrX	5730792	-	.	60	93	10946927_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10946927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_5708501_5733501_138C;SPAN=1666;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:147 DP:130 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:93 DR:60 LR:-435.7 LO:435.7);ALT=T]chrX:5730792];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	6010547	+	chrX	6004436	+	.	68	63	10947869_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10947869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_6002501_6027501_135C;SPAN=6111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:191 GQ:99 PL:[268.7, 0.0, 192.8] SR:63 DR:68 LR:-269.1 LO:269.1);ALT=]chrX:6010547]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	6933200	+	chrX	6942585	+	.	59	33	10952136_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10952136_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_6909001_6934001_202C;SPAN=9385;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:44 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:33 DR:59 LR:-227.8 LO:227.8);ALT=A[chrX:6942585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	7001689	+	chrX	7135424	+	CC	14	4	10952376_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CC;MAPQ=60;MATEID=10952376_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_6982501_7007501_249C;SPAN=133735;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:100 GQ:29 PL:[29.0, 0.0, 213.8] SR:4 DR:14 LR:-29.02 LO:37.19);ALT=C[chrX:7135424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	7029390	+	chrX	7069941	+	.	65	19	10952397_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GCT;MAPQ=60;MATEID=10952397_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_7056001_7081001_17C;SPAN=40551;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:28 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:19 DR:65 LR:-211.3 LO:211.3);ALT=T[chrX:7069941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	7623882	+	chrX	7673883	+	.	124	115	10954579_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=10954579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_7668501_7693501_186C;SPAN=50001;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:192 DP:17 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:115 DR:124 LR:-567.7 LO:567.7);ALT=C[chrX:7673883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	10738668	+	chrX	10788674	+	.	134	0	10968469_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=10968469_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:10738668(+)-23:10788674(-)__23_10780001_10805001D;SPAN=50006;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:6 GQ:36 PL:[396.0, 36.0, 0.0] SR:0 DR:134 LR:-396.1 LO:396.1);ALT=A[chrX:10788674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	84823534	+	chrX	11042090	+	TTGGTGACCTTTGA	7	42	11285111_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;INSERTION=TTGGTGACCTTTGA;MAPQ=38;MATEID=11285111_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_23_84819001_84844001_126C;SPAN=73781444;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:71 GQ:27.2 PL:[142.7, 0.0, 27.2] SR:42 DR:7 LR:-146.7 LO:146.7);ALT=]chrX:84823534]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	11953199	+	chrX	11959436	+	.	69	33	10973040_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGGTGATTTTTTTT;MAPQ=60;MATEID=10973040_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_11931501_11956501_197C;SPAN=6237;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:65 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:33 DR:69 LR:-260.8 LO:260.8);ALT=T[chrX:11959436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	13675608	-	chrX	13678652	+	.	10	0	10980287_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10980287_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:13675608(-)-23:13678652(-)__23_13671001_13696001D;SPAN=3044;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:129 GQ:1.8 PL:[0.0, 1.8, 316.8] SR:0 DR:10 LR:1.939 LO:18.23);ALT=[chrX:13678652[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	48134220	+	chrX	48037226	+	.	8	0	11145948_1	10.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=11145948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48037226(-)-23:48134220(+)__23_48118001_48143001D;SPAN=96994;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=]chrX:48134220]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	48091714	+	chrX	48093011	+	.	31	0	11145762_1	82.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=11145762_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48091714(+)-23:48093011(-)__23_48069001_48094001D;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:75 GQ:82.1 PL:[82.1, 0.0, 98.6] SR:0 DR:31 LR:-82.01 LO:82.11);ALT=T[chrX:48093011[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48104369	+	chrX	48306103	-	.	25	0	11145582_1	72.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=11145582_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48104369(+)-23:48306103(+)__23_48093501_48118501D;SPAN=201734;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:25 DP:20 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:0 DR:25 LR:-72.62 LO:72.62);ALT=T]chrX:48306103];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	48104636	-	chrX	48305935	+	.	17	0	11145584_1	42.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=11145584_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48104636(-)-23:48305935(-)__23_48093501_48118501D;SPAN=201299;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:0 DR:17 LR:-42.84 LO:43.35);ALT=[chrX:48305935[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	48140635	+	chrX	52641884	+	.	25	0	11146065_1	65.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=11146065_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48140635(+)-23:52641884(-)__23_48118001_48143001D;SPAN=4501249;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:65 GQ:65 PL:[65.0, 0.0, 91.4] SR:0 DR:25 LR:-64.92 LO:65.19);ALT=T[chrX:52641884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	52642058	+	chrX	48140737	+	.	16	0	11146066_1	42.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=11146066_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48140737(-)-23:52642058(+)__23_48118001_48143001D;SPAN=4501321;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:38 GQ:42.5 PL:[42.5, 0.0, 49.1] SR:0 DR:16 LR:-42.52 LO:42.55);ALT=]chrX:52642058]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	54002189	+	chrX	53742007	+	.	58	13	11174110_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=11174110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_53998001_54023001_199C;SPAN=260182;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:81 GQ:11.3 PL:[182.9, 0.0, 11.3] SR:13 DR:58 LR:-191.3 LO:191.3);ALT=]chrX:54002189]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	54938971	-	chrX	54940218	+	.	9	0	11178673_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=11178673_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:54938971(-)-23:54940218(-)__23_54929001_54954001D;SPAN=1247;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:142 GQ:8.4 PL:[0.0, 8.4, 359.7] SR:0 DR:9 LR:8.762 LO:15.59);ALT=[chrX:54940218[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	55702405	+	chrX	55709883	+	.	53	0	11182734_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=11182734_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:55702405(+)-23:55709883(-)__23_55688501_55713501D;SPAN=7478;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:50 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:0 DR:53 LR:-155.1 LO:155.1);ALT=G[chrX:55709883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	75417348	+	chrX	75298131	+	.	72	36	11250413_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=11250413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_75411001_75436001_80C;SPAN=119217;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:69 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:36 DR:72 LR:-280.6 LO:280.6);ALT=]chrX:75417348]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	76508484	-	chrX	76510025	+	.	10	0	11254711_1	2.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=11254711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:76508484(-)-23:76510025(-)__23_76489001_76514001D;SPAN=1541;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:115 GQ:2 PL:[2.0, 0.0, 275.9] SR:0 DR:10 LR:-1.854 LO:18.75);ALT=[chrX:76510025[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	77121417	+	chrX	77123867	+	.	88	43	11256835_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTCACGCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=60;MATEID=11256835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_77101501_77126501_416C;SPAN=2450;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:107 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:43 DR:88 LR:-346.6 LO:346.6);ALT=C[chrX:77123867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	81096653	+	chrX	81102693	+	.	62	39	11271553_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGGCAATTTGG;MAPQ=60;MATEID=11271553_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_81095001_81120001_237C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:81 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:39 DR:62 LR:-247.6 LO:247.6);ALT=G[chrX:81102693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	81982373	+	chrX	81988116	+	.	45	0	11274717_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=11274717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:81982373(+)-23:81988116(-)__23_81977001_82002001D;SPAN=5743;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:99 GQ:99 PL:[121.7, 0.0, 118.4] SR:0 DR:45 LR:-121.7 LO:121.7);ALT=G[chrX:81988116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	84096004	+	chrX	84145023	-	.	20	43	11282007_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAA;MAPQ=60;MATEID=11282007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_84133001_84158001_74C;SPAN=49019;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:61 DP:71 GQ:12.3 PL:[194.7, 12.3, 0.0] SR:43 DR:20 LR:-196.2 LO:196.2);ALT=A]chrX:84145023];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	84098028	-	chrX	84144890	+	.	8	0	11282008_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=11282008_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:84098028(-)-23:84144890(-)__23_84133001_84158001D;SPAN=46862;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=[chrX:84144890[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	85605183	+	chrX	85609864	+	.	114	75	11287981_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=AAAACAAAACAA;MAPQ=60;MATEID=11287981_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_85603001_85628001_68C;SPAN=4681;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:169 DP:36 GQ:45.7 PL:[501.7, 45.7, 0.0] SR:75 DR:114 LR:-501.7 LO:501.7);ALT=A[chrX:85609864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	86279051	+	chrX	86280137	+	TG	0	60	11290173_1	99.0	.	EVDNC=ASSMB;INSERTION=TG;MAPQ=60;MATEID=11290173_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_86264501_86289501_372C;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:66 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:60 DR:0 LR:-194.7 LO:194.7);ALT=A[chrX:86280137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	123127643	+	chrX	123122701	+	.	60	49	11370567_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=11370567_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_123112501_123137501_246C;SPAN=4942;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:87 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:49 DR:60 LR:-274.0 LO:274.0);ALT=]chrX:123127643]G;VARTYPE=BND:DUP-th;JOINTYPE=th
