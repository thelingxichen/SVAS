chr5	23065367	-	chr5	23067021	+	.	9	0	3287426_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3287426_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:23065367(-)-5:23067021(-)__5_23054501_23079501D;SPAN=1654;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:199 GQ:24.1 PL:[0.0, 24.1, 531.4] SR:0 DR:9 LR:24.21 LO:14.25);ALT=[chr5:23067021[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
