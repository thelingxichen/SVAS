chr2	53992724	+	chr2	54013958	+	.	13	3	797190_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=797190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_53998001_54023001_75C;SPAN=21234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:44 GQ:37.7 PL:[37.7, 0.0, 67.4] SR:3 DR:13 LR:-37.59 LO:38.11);ALT=T[chr2:54013958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	54111588	+	chr14	40317397	-	.	12	47	5714070_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GGATCACAAGGTCAAGAGATTGAGACCATCCTGGCCAACATG;MAPQ=49;MATEID=5714070_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_14_40302501_40327501_111C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:25 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:47 DR:12 LR:-174.9 LO:174.9);ALT=C]chr14:40317397];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	54342895	+	chr2	54365775	+	GTTTGCTTCAGAAT	11	6	798064_1	22.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=GTTTGCTTCAGAAT;MAPQ=60;MATEID=798064_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_2_54365501_54390501_264C;SPAN=22880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:6 DR:11 LR:-22.49 LO:25.34);ALT=T[chr2:54365775[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	54565493	+	chr2	54567474	+	TA	62	24	798570_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TA;MAPQ=0;MATEID=798570_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_54561501_54586501_287C;SPAN=1981;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:55 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:24 DR:62 LR:-217.9 LO:217.9);ALT=G[chr2:54567474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55200334	+	chr2	55201831	+	TTAGCCATAGCATCTTTAACATTCTTATTTGCAAGTCCTAGATAATGATCTATCTGTGCCTGATGCCGTTCATAAATAACAGGAACACTGAAGAGTGAAATGAGAG	3	18	800178_1	33.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTAGCCATAGCATCTTTAACATTCTTATTTGCAAGTCCTAGATAATGATCTATCTGTGCCTGATGCCGTTCATAAATAACAGGAACACTGAAGAGTGAAATGAGAG;MAPQ=60;MATEID=800178_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_55198501_55223501_256C;SPAN=1497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:96 GQ:33.5 PL:[33.5, 0.0, 198.5] SR:18 DR:3 LR:-33.41 LO:40.23);ALT=T[chr2:55201831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55201902	+	chr2	55209651	+	.	2	9	800183_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=800183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_55198501_55223501_162C;SPAN=7749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:9 DR:2 LR:-13.82 LO:22.76);ALT=T[chr2:55209651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55209791	+	chr2	55214626	+	.	8	3	800211_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=800211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_55198501_55223501_146C;SPAN=4835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:3 DR:8 LR:-10.79 LO:20.31);ALT=T[chr2:55214626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55214835	+	chr2	55237223	+	.	3	4	800224_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=800224_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_55198501_55223501_44C;SPAN=22388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:41 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:4 DR:3 LR:-5.397 LO:10.15);ALT=C[chr2:55237223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55746950	+	chr2	55749235	+	.	11	0	801847_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=801847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:55746950(+)-2:55749235(-)__2_55737501_55762501D;SPAN=2285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:0 DR:11 LR:-11.39 LO:22.24);ALT=G[chr2:55749235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55747052	+	chr2	55750857	+	TTTTTGATGATGAAGAAGAAAGCAAATTGACCTATACAGAGATTCATCAGGAATACAAAGAACTA	7	28	801849_1	78.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=TTTTTGATGATGAAGAAGAAAGCAAATTGACCTATACAGAGATTCATCAGGAATACAAAGAACTA;MAPQ=60;MATEID=801849_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_55737501_55762501_69C;SPAN=3805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:88 GQ:78.5 PL:[78.5, 0.0, 134.6] SR:28 DR:7 LR:-78.49 LO:79.31);ALT=G[chr2:55750857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	55750959	+	chr2	55761008	+	CCATTTTGCAACCTGTGTTGGCAGCAGAAGATTTTACTATCTTTAAAGCAATGATGGTCCAGAAAAACATTGAAATGCAGCTGCAAGCCATTCGAATAATTCAAGAGAGAAAT	0	15	801875_1	31.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=CCATTTTGCAACCTGTGTTGGCAGCAGAAGATTTTACTATCTTTAAAGCAATGATGGTCCAGAAAAACATTGAAATGCAGCTGCAAGCCATTCGAATAATTCAAGAGAGAAAT;MAPQ=60;MATEID=801875_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_55737501_55762501_52C;SPAN=10049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:66 GQ:31.7 PL:[31.7, 0.0, 127.4] SR:15 DR:0 LR:-31.63 LO:34.94);ALT=G[chr2:55761008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	56652302	+	chr2	56655883	+	AA	19	16	804356_1	85.0	.	DISC_MAPQ=15;EVDNC=ASDIS;INSERTION=AA;MAPQ=0;MATEID=804356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_56644001_56669001_119C;SPAN=3581;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:64 GQ:68.6 PL:[85.1, 0.0, 68.6] SR:16 DR:19 LR:-85.06 LO:85.06);ALT=G[chr2:56655883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39644642	+	chr14	39645749	+	.	16	0	5711875_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5711875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:39644642(+)-14:39645749(-)__14_39641001_39666001D;SPAN=1107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:122 GQ:20 PL:[20.0, 0.0, 274.1] SR:0 DR:16 LR:-19.76 LO:33.03);ALT=C[chr14:39645749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39645354	+	chr14	39646614	+	CGTGGATTCTCAGATAGTGGAGGAGGACCCCCAGCCAAACAGAGAGACCTTGAAGGGGCAGTCAGT	0	98	5711878_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CGTGGATTCTCAGATAGTGGAGGAGGACCCCCAGCCAAACAGAGAGACCTTGAAGGGGCAGTCAGT;MAPQ=60;MATEID=5711878_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_39641001_39666001_271C;SPAN=1260;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:98 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:98 DR:0 LR:-290.5 LO:290.5);ALT=G[chr14:39646614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39646892	+	chr14	39648294	+	AACCGGCGAATATTTGGCTTGTTGATGGGTACCCTTCAAAAATTTAAACAAGAATCCACTGTTGCTACTGAAAG	0	25	5711884_1	58.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AACCGGCGAATATTTGGCTTGTTGATGGGTACCCTTCAAAAATTTAAACAAGAATCCACTGTTGCTACTGAAAG;MAPQ=60;MATEID=5711884_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_39641001_39666001_47C;SPAN=1402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:88 GQ:58.7 PL:[58.7, 0.0, 154.4] SR:25 DR:0 LR:-58.68 LO:61.08);ALT=G[chr14:39648294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39647120	+	chr14	39648294	+	.	6	12	5711885_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5711885_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_14_39641001_39666001_47C;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:81 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:12 DR:6 LR:-27.57 LO:33.43);ALT=G[chr14:39648294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39648666	+	chr14	39649706	+	.	21	23	5711891_1	93.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5711891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_39641001_39666001_226C;SPAN=1040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:94 GQ:93.5 PL:[93.5, 0.0, 133.1] SR:23 DR:21 LR:-93.37 LO:93.78);ALT=G[chr14:39649706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39736728	+	chr14	39746137	+	.	5	4	5712301_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5712301_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_39739001_39764001_135C;SPAN=9409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:36 GQ:13.4 PL:[13.4, 0.0, 72.8] SR:4 DR:5 LR:-13.35 LO:15.77);ALT=T[chr14:39746137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	40098409	+	chr14	40100214	+	.	69	36	5713221_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAGTCCTGAAATAACTT;MAPQ=60;MATEID=5713221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_40082001_40107001_239C;SPAN=1805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:22 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:36 DR:69 LR:-247.6 LO:247.6);ALT=T[chr14:40100214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	40609815	+	chr14	40617673	+	CAGGCTCCTTTGTAAATAA	0	59	5713997_1	99.0	.	EVDNC=ASSMB;INSERTION=CAGGCTCCTTTGTAAATAA;MAPQ=60;MATEID=5713997_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_40596501_40621501_82C;SPAN=7858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:25 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:59 DR:0 LR:-174.9 LO:174.9);ALT=A[chr14:40617673[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
