chr9	77131030	-	chr9	77132356	+	.	8	0	4277475_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4277475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:77131030(-)-9:77132356(-)__9_77126001_77151001D;SPAN=1326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=[chr9:77132356[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	77703643	+	chr9	77745493	+	GCAAGTTAAAGTCTTCAGAGCCCTGTATACGTTTGAACCCAGAACTCCAGATGAATTATACTTTGAGGAAGGTGATATTATCTACATTACTGACAT	0	96	4279400_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GCAAGTTAAAGTCTTCAGAGCCCTGTATACGTTTGAACCCAGAACTCCAGATGAATTATACTTTGAGGAAGGTGATATTATCTACATTACTGACAT;MAPQ=60;MATEID=4279400_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_9_77738501_77763501_2C;SPAN=41850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:47 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:96 DR:0 LR:-283.9 LO:283.9);ALT=G[chr9:77745493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	77755848	+	chr9	77761596	+	.	2	6	4279460_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4279460_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_77738501_77763501_306C;SPAN=5748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:93 GQ:1.8 PL:[0.0, 1.8, 227.7] SR:6 DR:2 LR:2.089 LO:12.67);ALT=G[chr9:77761596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
