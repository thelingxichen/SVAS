chrX	72652681	+	chrX	72916723	+	.	0	10	11239442_1	17.0	.	EVDNC=ASSMB;HOMSEQ=ATCTCTCAGCA;MAPQ=60;MATEID=11239442_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_72642501_72667501_220C;SPAN=264042;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=A[chrX:72916723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
