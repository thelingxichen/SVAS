chr3	80925314	+	chr3	80926605	+	.	29	18	1506983_1	97.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=1506983_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_80923501_80948501_64C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:273 GQ:97.9 PL:[97.9, 0.0, 563.3] SR:18 DR:29 LR:-97.69 LO:116.6);ALT=T[chr3:80926605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
