chr20	7096793	+	chr20	7102847	+	.	37	32	10415730_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GACAAAATTTTT;MAPQ=60;MATEID=10415730_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_7080501_7105501_186C;SPAN=6054;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:57 DP:29 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:32 DR:37 LR:-168.3 LO:168.3);ALT=T[chr20:7102847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
