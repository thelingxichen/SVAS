chr20	42024612	+	chr20	42025793	+	.	95	20	7019739_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGGTAAAACCCCATTTCT;MAPQ=0;MATEID=7019739_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_42017501_42042501_270C;SECONDARY;SPAN=1181;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:30 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:20 DR:95 LR:-310.3 LO:310.3);ALT=T[chr20:42025793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42219700	+	chr20	42223330	+	.	14	0	7020730_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7020730_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:42219700(+)-20:42223330(-)__20_42213501_42238501D;SPAN=3630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:117 GQ:14.6 PL:[14.6, 0.0, 268.7] SR:0 DR:14 LR:-14.52 LO:28.31);ALT=G[chr20:42223330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42223457	+	chr20	42225073	+	.	0	14	7020740_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7020740_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_42213501_42238501_54C;SPAN=1616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:14 DR:0 LR:-21.29 LO:29.89);ALT=G[chr20:42225073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42271920	+	chr20	42274577	+	.	89	0	7020847_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7020847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:42271920(+)-20:42274577(-)__20_42262501_42287501D;SPAN=2657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:13 GQ:24 PL:[264.0, 24.0, 0.0] SR:0 DR:89 LR:-264.1 LO:264.1);ALT=G[chr20:42274577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42481277	+	chr20	42483783	+	.	51	32	7021824_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GCCCAGCTA;MAPQ=60;MATEID=7021824_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_42483001_42508001_128C;SPAN=2506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:30 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:32 DR:51 LR:-224.5 LO:224.5);ALT=A[chr20:42483783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	42826380	+	chr20	42831599	+	.	2	2	7023112_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=7023112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_42826001_42851001_346C;SPAN=5219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:2 DR:2 LR:13.62 LO:6.133);ALT=C[chr20:42831599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43142727	+	chr20	43150612	+	.	21	0	7024531_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7024531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:43142727(+)-20:43150612(-)__20_43120001_43145001D;SPAN=7885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:56 GQ:54.2 PL:[54.2, 0.0, 80.6] SR:0 DR:21 LR:-54.15 LO:54.46);ALT=T[chr20:43150612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43160671	+	chr20	43243171	+	.	19	0	7024747_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7024747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:43160671(+)-20:43243171(-)__20_43242501_43267501D;SPAN=82500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:74 GQ:42.8 PL:[42.8, 0.0, 135.2] SR:0 DR:19 LR:-42.67 LO:45.43);ALT=T[chr20:43243171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43218508	+	chr20	43243172	+	.	0	14	7024749_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=7024749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43242501_43267501_46C;SPAN=24664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:14 DR:0 LR:-26.17 LO:31.35);ALT=G[chr20:43243172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43255240	+	chr20	43257687	+	.	2	24	7024789_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7024789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43242501_43267501_317C;SPAN=2447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:120 GQ:53.3 PL:[53.3, 0.0, 238.1] SR:24 DR:2 LR:-53.32 LO:59.95);ALT=C[chr20:43257687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43255286	+	chr20	43280270	+	.	13	0	7025016_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=7025016_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:43255286(+)-20:43280270(-)__20_43267001_43292001D;SPAN=24984;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:51 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:0 DR:13 LR:-29.1 LO:31.04);ALT=T[chr20:43280270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43257813	+	chr20	43280214	+	CCATAGTATAAGATGGTTTCAGGCTTGATGGATCCGTCTAGGTGGACATGCAGTTCT	79	91	7025018_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=CCATAGTATAAGATGGTTTCAGGCTTGATGGATCCGTCTAGGTGGACATGCAGTTCT;MAPQ=60;MATEID=7025018_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_43267001_43292001_375C;SPAN=22401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:47 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:91 DR:79 LR:-392.8 LO:392.8);ALT=G[chr20:43280214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43264926	+	chr20	43280214	+	T	45	41	7025019_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CCTG;INSERTION=T;MAPQ=60;MATEID=7025019_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_43267001_43292001_375C;SPAN=15288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:47 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:41 DR:45 LR:-158.4 LO:158.4);ALT=C[chr20:43280214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43514528	+	chr20	43530171	+	.	93	74	7025943_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7025943_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43512001_43537001_89C;SPAN=15643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:166 GQ:28.3 PL:[458.8, 28.3, 0.0] SR:74 DR:93 LR:-465.2 LO:465.2);ALT=G[chr20:43530171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43514528	+	chr20	43516288	+	.	0	11	7025942_1	1.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=7025942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43512001_43537001_379C;SPAN=1760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:131 GQ:1.1 PL:[1.1, 0.0, 314.6] SR:11 DR:0 LR:-0.8199 LO:20.45);ALT=G[chr20:43516288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43516384	+	chr20	43530170	+	.	0	11	7025948_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7025948_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43512001_43537001_283C;SPAN=13786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:132 GQ:0.8 PL:[0.8, 0.0, 317.6] SR:11 DR:0 LR:-0.549 LO:20.42);ALT=G[chr20:43530170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43530475	+	chr20	43532633	+	.	8	9	7026000_1	12.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7026000_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43512001_43537001_209C;SPAN=2158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:99 GQ:12.8 PL:[12.8, 0.0, 227.3] SR:9 DR:8 LR:-12.79 LO:24.33);ALT=G[chr20:43532633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43532757	+	chr20	43534641	+	CCACTGTGTCGAACTCCCAGCAGGCTTACCAGGAAGCATTTGAAATTAGTAAGAAAGAAATGCAGCCTACACACCCAATTCGTCTTGGTCTGGCACTAAATTTCTCAGTCTTTTACTATGAGATTCTAAACTCTCCTGAAAAGGCCTGTAGCCTGGCAAAAAC	0	51	7026009_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=CCACTGTGTCGAACTCCCAGCAGGCTTACCAGGAAGCATTTGAAATTAGTAAGAAAGAAATGCAGCCTACACACCCAATTCGTCTTGGTCTGGCACTAAATTTCTCAGTCTTTTACTATGAGATTCTAAACTCTCCTGAAAAGGCCTGTAGCCTGGCAAAAAC;MAPQ=60;MATEID=7026009_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_43512001_43537001_27C;SPAN=1884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:115 GQ:99 PL:[137.3, 0.0, 140.6] SR:51 DR:0 LR:-137.2 LO:137.2);ALT=A[chr20:43534641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43547919	+	chr20	43550233	+	.	2	2	7025759_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7025759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43536501_43561501_105C;SPAN=2314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:121 GQ:19.2 PL:[0.0, 19.2, 330.0] SR:2 DR:2 LR:19.58 LO:5.781);ALT=G[chr20:43550233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43585128	+	chr20	43588846	+	.	0	16	7026129_1	41.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=7026129_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43561001_43586001_37C;SPAN=3718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:42 GQ:41.6 PL:[41.6, 0.0, 58.1] SR:16 DR:0 LR:-41.44 LO:41.63);ALT=T[chr20:43588846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43595245	+	chr20	43600718	+	.	87	10	7026193_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7026193_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43585501_43610501_190C;SPAN=5473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:135 GQ:69.2 PL:[257.3, 0.0, 69.2] SR:10 DR:87 LR:-263.1 LO:263.1);ALT=G[chr20:43600718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43595277	+	chr20	43607081	+	.	26	0	7026196_1	51.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7026196_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:43595277(+)-20:43607081(-)__20_43585501_43610501D;SPAN=11804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:126 GQ:51.8 PL:[51.8, 0.0, 253.1] SR:0 DR:26 LR:-51.69 LO:59.32);ALT=G[chr20:43607081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43600801	+	chr20	43607083	+	.	0	21	7026222_1	31.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7026222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43585501_43610501_155C;SPAN=6282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:142 GQ:31.1 PL:[31.1, 0.0, 311.6] SR:21 DR:0 LR:-30.85 LO:44.54);ALT=T[chr20:43607083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43607212	+	chr20	43610468	+	.	0	16	7026245_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7026245_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43585501_43610501_304C;SPAN=3256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:116 GQ:21.5 PL:[21.5, 0.0, 259.1] SR:16 DR:0 LR:-21.39 LO:33.41);ALT=G[chr20:43610468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43630000	+	chr20	43653618	+	.	2	2	7026454_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7026454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43610001_43635001_299C;SPAN=23618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:42 GQ:2 PL:[2.0, 0.0, 97.7] SR:2 DR:2 LR:-1.825 LO:7.667);ALT=G[chr20:43653618[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	43994326	+	chr20	43995514	+	.	0	5	7027575_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7027575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_43977501_44002501_37C;SPAN=1188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:113 GQ:13.8 PL:[0.0, 13.8, 300.3] SR:5 DR:0 LR:14.11 LO:7.866);ALT=G[chr20:43995514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44050225	+	chr20	44052856	+	.	2	3	7028103_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=7028103_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_44051001_44076001_330C;SPAN=2631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:67 GQ:4.8 PL:[0.0, 4.8, 171.6] SR:3 DR:2 LR:4.948 LO:6.824);ALT=T[chr20:44052856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44326234	-	chr20	44327395	+	.	8	0	7028731_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7028731_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:44326234(-)-20:44327395(-)__20_44320501_44345501D;SPAN=1161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:0 DR:8 LR:5.561 LO:14.1);ALT=[chr20:44327395[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	44420722	+	chr20	44422557	+	.	13	0	7029402_1	13.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7029402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:44420722(+)-20:44422557(-)__20_44418501_44443501D;SPAN=1835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:111 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:0 DR:13 LR:-12.84 LO:26.15);ALT=G[chr20:44422557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44421386	+	chr20	44422558	+	.	0	21	7029407_1	37.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7029407_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_44418501_44443501_403C;SPAN=1172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:117 GQ:37.7 PL:[37.7, 0.0, 245.6] SR:21 DR:0 LR:-37.62 LO:46.49);ALT=G[chr20:44422558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44441395	+	chr20	44443021	+	.	11	0	7029483_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7029483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:44441395(+)-20:44443021(-)__20_44418501_44443501D;SPAN=1626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:103 GQ:8.6 PL:[8.6, 0.0, 239.6] SR:0 DR:11 LR:-8.406 LO:21.66);ALT=G[chr20:44443021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44441436	+	chr20	44444179	+	CTACAGCAGGAGCTGATGACCCTCAT	6	7	7029485_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTACAGCAGGAGCTGATGACCCTCAT;MAPQ=60;MATEID=7029485_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_44418501_44443501_270C;SPAN=2743;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:52 GQ:22.4 PL:[22.4, 0.0, 101.6] SR:7 DR:6 LR:-22.22 LO:25.23);ALT=G[chr20:44444179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44483934	+	chr20	44485827	+	.	0	14	7029561_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7029561_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_44467501_44492501_420C;SPAN=1893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:126 GQ:12.2 PL:[12.2, 0.0, 292.7] SR:14 DR:0 LR:-12.08 LO:27.83);ALT=G[chr20:44485827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44523805	+	chr20	44526353	+	.	8	0	7029683_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7029683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:44523805(+)-20:44526353(-)__20_44516501_44541501D;SPAN=2548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=G[chr20:44526353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44563443	+	chr20	44566054	+	.	52	4	7030003_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7030003_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_44565501_44590501_403C;SPAN=2611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:52 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:4 DR:52 LR:-155.1 LO:155.1);ALT=G[chr20:44566054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44566226	+	chr20	44567619	+	.	0	4	7030006_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7030006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_44565501_44590501_182C;SPAN=1393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:137 GQ:23.7 PL:[0.0, 23.7, 379.5] SR:4 DR:0 LR:23.91 LO:5.565);ALT=T[chr20:44567619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	44987424	+	chr20	44993009	+	.	11	0	7031463_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7031463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:44987424(+)-20:44993009(-)__20_44982001_45007001D;SPAN=5585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:0 DR:11 LR:-12.74 LO:22.52);ALT=T[chr20:44993009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
