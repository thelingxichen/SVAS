chr1	209929596	+	chr1	209932375	+	.	17	0	523170_1	23.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=523170_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:209929596(+)-1:209932375(-)__1_209916001_209941001D;SPAN=2779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:123 GQ:23 PL:[23.0, 0.0, 273.8] SR:0 DR:17 LR:-22.79 LO:35.52);ALT=A[chr1:209932375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	209929654	+	chr1	209933324	+	CAGCCTTATTGAGGTACAATTCATGTGCTTGTGGGTTTGGATGGCACAATCTGTGTCTGGGCTAAGGAAAGCAGACTTGGCACCAACATTAACCCTGA	0	34	523172_1	81.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=CAGCCTTATTGAGGTACAATTCATGTGCTTGTGGGTTTGGATGGCACAATCTGTGTCTGGGCTAAGGAAAGCAGACTTGGCACCAACATTAACCCTGA;MAPQ=60;MATEID=523172_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_209916001_209941001_63C;SPAN=3670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:113 GQ:81.8 PL:[81.8, 0.0, 190.7] SR:34 DR:0 LR:-81.62 LO:84.1);ALT=G[chr1:209933324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	209946364	+	chr1	209948691	+	.	0	7	523336_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=523336_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_209940501_209965501_115C;SPAN=2327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=G[chr1:209948691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	210078055	+	chr1	210085978	+	GAATTA	85	72	523603_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GAATTA;MAPQ=60;MATEID=523603_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_210063001_210088001_187C;SPAN=7923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:36 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:72 DR:85 LR:-369.7 LO:369.7);ALT=A[chr1:210085978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
