chr5	98345117	+	chr5	98347483	+	AC	65	41	2537572_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=AC;MAPQ=60;MATEID=2537572_2;MATENM=1;NM=5;NUMPARTS=2;SCTG=c_5_98343001_98368001_118C;SPAN=2366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:19 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:41 DR:65 LR:-247.6 LO:247.6);ALT=C[chr5:98347483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	98610746	+	chr17	60434032	+	.	19	36	6459211_1	99.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=0;MATEID=6459211_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TATA;SCTG=c_17_60417001_60442001_337C;SECONDARY;SPAN=-1;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:45 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:36 DR:19 LR:-145.2 LO:145.2);ALT=G[chr17:60434032[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	98839889	+	chr5	98842907	+	TG	30	43	2538510_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;INSERTION=TG;MAPQ=11;MATEID=2538510_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_98833001_98858001_38C;SPAN=3018;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:19 GQ:15 PL:[165.0, 15.0, 0.0] SR:43 DR:30 LR:-165.0 LO:165.0);ALT=C[chr5:98842907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
