chr10	61450941	+	chr10	61452114	+	.	0	55	6298306_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6298306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_61446001_61471001_112C;SPAN=1173;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:87 GQ:52.4 PL:[158.0, 0.0, 52.4] SR:55 DR:0 LR:-160.8 LO:160.8);ALT=T[chr10:61452114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
