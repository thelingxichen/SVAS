chr7	22434803	+	chr7	22436761	+	.	171	107	4610043_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=4610043_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_22417501_22442501_259C;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:241 DP:118 GQ:64.9 PL:[712.9, 64.9, 0.0] SR:107 DR:171 LR:-713.0 LO:713.0);ALT=C[chr7:22436761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23320762	+	chr7	23321782	-	.	8	0	4616191_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4616191_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:23320762(+)-7:23321782(+)__7_23299501_23324501D;SPAN=1020;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:201 GQ:27.7 PL:[0.0, 27.7, 541.3] SR:0 DR:8 LR:28.05 LO:12.21);ALT=A]chr7:23321782];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	23815666	-	chr7	23838143	+	.	19	17	4620105_1	60.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGAAAAAGCCTTTGATAAAATT;MAPQ=60;MATEID=4620105_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_23814001_23839001_61C;SPAN=22477;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:181 GQ:60.1 PL:[60.1, 0.0, 377.0] SR:17 DR:19 LR:-59.9 LO:73.3);ALT=[chr7:23838143[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	23815979	+	chr7	23837984	-	.	16	0	4620112_1	0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4620112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:23815979(+)-7:23837984(+)__7_23814001_23839001D;SPAN=22005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:16 DP:201 GQ:1.3 PL:[0.0, 1.3, 488.5] SR:0 DR:16 LR:1.64 LO:29.36);ALT=G]chr7:23837984];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	24038165	+	chr7	24040071	+	.	172	148	4621632_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATAT;MAPQ=60;MATEID=4621632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_24034501_24059501_49C;SPAN=1906;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:252 DP:52 GQ:67.9 PL:[745.9, 67.9, 0.0] SR:148 DR:172 LR:-746.0 LO:746.0);ALT=T[chr7:24040071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
