chr8	130883742	+	chr8	130891635	+	.	2	20	4076250_1	44.0	.	DISC_MAPQ=36;EVDNC=ASDIS;MAPQ=60;MATEID=4076250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_130879001_130904001_216C;SPAN=7893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:94 GQ:44 PL:[44.0, 0.0, 182.6] SR:20 DR:2 LR:-43.85 LO:48.74);ALT=T[chr8:130891635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	130891764	+	chr8	131028614	+	.	12	0	4076858_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4076858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:130891764(+)-8:131028614(-)__8_131026001_131051001D;SPAN=136850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:10 GQ:3 PL:[33.0, 3.0, 0.0] SR:0 DR:12 LR:-33.01 LO:33.01);ALT=A[chr8:131028614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	130983244	+	chr8	131028615	+	.	17	12	4076863_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=4076863_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_131026001_131051001_431C;SPAN=45371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:11 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:12 DR:17 LR:-62.72 LO:62.72);ALT=G[chr8:131028615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	131274647	+	chr8	131248115	+	.	19	10	4077723_1	70.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=4077723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_131271001_131296001_34C;SPAN=26532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:45 GQ:37.4 PL:[70.4, 0.0, 37.4] SR:10 DR:19 LR:-70.82 LO:70.82);ALT=]chr8:131274647]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	131850749	+	chr8	131852739	+	A	43	31	4079267_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4079267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_131834501_131859501_262C;SPAN=1990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:48 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:31 DR:43 LR:-181.5 LO:181.5);ALT=A[chr8:131852739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
