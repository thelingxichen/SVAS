chr2	128839980	+	chr3	185150146	+	.	14	28	1331375_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTTTTGTGTTTTTAGTAGAGACAGGGTTTCAC;MAPQ=60;MATEID=1331375_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_128821001_128846001_640C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:38 DP:57 GQ:27.5 PL:[110.0, 0.0, 27.5] SR:28 DR:14 LR:-112.7 LO:112.7);ALT=C[chr3:185150146[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	129438422	+	chr13	53034838	+	.	13	0	8075149_1	28.0	.	DISC_MAPQ=8;EVDNC=DSCRD;IMPRECISE;MAPQ=8;MATEID=8075149_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:129438422(+)-13:53034838(-)__13_53018001_53043001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:0 DR:13 LR:-28.55 LO:30.78);ALT=C[chr13:53034838[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	129560395	+	chr2	129561909	+	.	58	35	1333057_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=1333057_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_129556001_129581001_155C;SPAN=1514;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:61 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:35 DR:58 LR:-208.0 LO:208.0);ALT=T[chr2:129561909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	129638421	+	chr2	129646204	+	.	72	63	1333148_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=1333148_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_129629501_129654501_359C;SPAN=7783;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:120 GQ:19.2 PL:[330.0, 19.2, 0.0] SR:63 DR:72 LR:-335.9 LO:335.9);ALT=C[chr2:129646204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	129703738	+	chr2	129722264	-	.	58	0	1334207_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=1334207_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:129703738(+)-2:129722264(+)__2_129703001_129728001D;SPAN=18526;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:113 GQ:99 PL:[161.0, 0.0, 111.5] SR:0 DR:58 LR:-161.3 LO:161.3);ALT=T]chr2:129722264];VARTYPE=BND:INV-hh;JOINTYPE=hh
