chr7	16171773	+	chr7	16174073	+	.	72	53	3183590_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3183590_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_16170001_16195001_353C;SPAN=2300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:76 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:53 DR:72 LR:-293.8 LO:293.8);ALT=C[chr7:16174073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16291092	-	chr7	16293041	+	.	14	0	3184069_1	31.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=3184069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:16291092(-)-7:16293041(-)__7_16292501_16317501D;SPAN=1949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:55 GQ:31.4 PL:[31.4, 0.0, 100.7] SR:0 DR:14 LR:-31.31 LO:33.42);ALT=[chr7:16293041[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	16685913	+	chr7	16705059	+	.	27	11	3185280_1	65.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=3185280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_16684501_16709501_270C;SPAN=19146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:114 GQ:65 PL:[65.0, 0.0, 210.2] SR:11 DR:27 LR:-64.84 LO:69.21);ALT=G[chr7:16705059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16685964	+	chr7	16714034	+	.	71	0	3185366_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3185366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:16685964(+)-7:16714034(-)__7_16709001_16734001D;SPAN=28070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:53 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=A[chr7:16714034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16705126	+	chr7	16720925	+	ATGAAAAAGAGAAATTCGAACCCACAGTCTTCAGGGATACACTTGTCCAGGGGCTTAATGAGGCTGGTGATGACCTTGAAGCTGTAGCCAAATTTCTGGACTCTACAGGCTCAAGATTAGATTATCGTCGCTATGCAGACACACTCTTCGATATCCTGGTGGCTGGCAGTATGCTT	0	67	3185351_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGAAAAAGAGAAATTCGAACCCACAGTCTTCAGGGATACACTTGTCCAGGGGCTTAATGAGGCTGGTGATGACCTTGAAGCTGTAGCCAAATTTCTGGACTCTACAGGCTCAAGATTAGATTATCGTCGCTATGCAGACACACTCTTCGATATCCTGGTGGCTGGCAGTATGCTT;MAPQ=60;MATEID=3185351_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_16684501_16709501_51C;SPAN=15799;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:65 GQ:18 PL:[198.0, 18.0, 0.0] SR:67 DR:0 LR:-198.0 LO:198.0);ALT=G[chr7:16720925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16714213	+	chr7	16720925	+	.	4	14	3185382_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3185382_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_7_16709001_16734001_103C;SPAN=6712;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:103 GQ:25.1 PL:[25.1, 0.0, 223.1] SR:14 DR:4 LR:-24.91 LO:34.31);ALT=G[chr7:16720925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16737811	+	chr7	16744170	+	.	4	9	3185553_1	13.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3185553_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_16733501_16758501_172C;SPAN=6359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:96 GQ:13.7 PL:[13.7, 0.0, 218.3] SR:9 DR:4 LR:-13.6 LO:24.51);ALT=G[chr7:16744170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16737811	+	chr7	16745683	+	CTGATGTTCTGAGCGAAGAAGCAATACTGAAATGGTATAAGGAAGCACATGTTGCTAAAGGCAAAAGTGTTTTTCTTGACCAGATGAAGAAATTTGTTGAGTGGTTACAAAATGCAGAAGA	4	25	3185554_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTGATGTTCTGAGCGAAGAAGCAATACTGAAATGGTATAAGGAAGCACATGTTGCTAAAGGCAAAAGTGTTTTTCTTGACCAGATGAAGAAATTTGTTGAGTGGTTACAAAATGCAGAAGA;MAPQ=60;MATEID=3185554_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_16733501_16758501_172C;SPAN=7872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:112 GQ:52.4 PL:[52.4, 0.0, 217.4] SR:25 DR:4 LR:-52.18 LO:58.02);ALT=G[chr7:16745683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16744294	+	chr7	16745683	+	.	2	12	3185570_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3185570_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_7_16733501_16758501_172C;SPAN=1389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:118 GQ:4.6 PL:[4.6, 0.0, 207.4] SR:12 DR:2 LR:-4.459 LO:18.53);ALT=G[chr7:16745683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16793655	+	chr7	16815836	+	.	0	8	3185928_1	8.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3185928_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_16782501_16807501_82C;SPAN=22181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:8 DR:0 LR:-8.798 LO:16.28);ALT=C[chr7:16815836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	16841462	+	chr7	16844558	+	.	41	0	3185666_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3185666_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:16841462(+)-7:16844558(-)__7_16831501_16856501D;SPAN=3096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:115 GQ:99 PL:[104.3, 0.0, 173.6] SR:0 DR:41 LR:-104.2 LO:105.2);ALT=A[chr7:16844558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	17349747	+	chr7	17362124	+	.	2	6	3187374_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3187374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_17346001_17371001_90C;SPAN=12377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:111 GQ:6.6 PL:[0.0, 6.6, 280.5] SR:6 DR:2 LR:6.966 LO:12.11);ALT=G[chr7:17362124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	17370511	+	chr7	17373535	+	.	9	17	3187502_1	46.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3187502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_17370501_17395501_284C;SPAN=3024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:108 GQ:46.7 PL:[46.7, 0.0, 215.0] SR:17 DR:9 LR:-46.66 LO:52.84);ALT=G[chr7:17373535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	18330138	+	chr7	18365134	+	.	10	10	3190282_1	33.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3190282_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_18326001_18351001_68C;SPAN=34996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:59 GQ:33.5 PL:[33.5, 0.0, 109.4] SR:10 DR:10 LR:-33.53 LO:35.79);ALT=G[chr7:18365134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	18330182	+	chr7	18367067	+	.	30	0	3190283_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3190283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:18330182(+)-7:18367067(-)__7_18326001_18351001D;SPAN=36885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:49 GQ:32.9 PL:[85.7, 0.0, 32.9] SR:0 DR:30 LR:-87.03 LO:87.03);ALT=A[chr7:18367067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	18365215	+	chr7	18367068	+	.	0	14	3190242_1	17.0	.	EVDNC=ASSMB;HOMSEQ=ACAG;MAPQ=60;MATEID=3190242_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_18350501_18375501_88C;SPAN=1853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:108 GQ:17 PL:[17.0, 0.0, 244.7] SR:14 DR:0 LR:-16.95 LO:28.83);ALT=G[chr7:18367068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
