chr18	18571289	+	chr18	18572791	+	.	2	3	6553802_1	6.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6553802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_18546501_18571501_24C;SPAN=1502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:38 GQ:6.2 PL:[6.2, 0.0, 85.4] SR:3 DR:2 LR:-6.21 LO:10.33);ALT=T[chr18:18572791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	19192404	+	chr18	19202684	+	.	7	14	6555591_1	33.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6555591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_19183501_19208501_348C;SPAN=10280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:14 DR:7 LR:-33.63 LO:38.73);ALT=G[chr18:19202684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	19192421	+	chr18	19203705	+	.	47	0	6555592_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6555592_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:19192421(+)-18:19203705(-)__18_19183501_19208501D;SPAN=11284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:87 GQ:78.8 PL:[131.6, 0.0, 78.8] SR:0 DR:47 LR:-132.3 LO:132.3);ALT=G[chr18:19203705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
