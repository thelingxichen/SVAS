chr17	75073118	-	chr17	75074901	+	.	17	0	9821917_1	23.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=9821917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:75073118(-)-17:75074901(-)__17_75068001_75093001D;SPAN=1783;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:122 GQ:23.3 PL:[23.3, 0.0, 270.8] SR:0 DR:17 LR:-23.06 LO:35.58);ALT=[chr17:75074901[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
