chr10	18850429	+	chr10	18858152	-	.	8	0	4532920_1	3.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=4532920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:18850429(+)-10:18858152(+)__10_18840501_18865501D;SPAN=7723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=G]chr10:18858152];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	18858636	+	chr10	18857446	+	.	17	0	4532967_1	31.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4532967_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:18857446(-)-10:18858636(+)__10_18840501_18865501D;SPAN=1190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:91 GQ:31.7 PL:[31.7, 0.0, 186.8] SR:0 DR:17 LR:-31.46 LO:37.96);ALT=]chr10:18858636]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	18861400	+	chr10	18860398	+	.	14	0	4532977_1	21.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4532977_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:18860398(-)-10:18861400(+)__10_18840501_18865501D;SPAN=1002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:90 GQ:21.8 PL:[21.8, 0.0, 196.7] SR:0 DR:14 LR:-21.83 LO:30.03);ALT=]chr10:18861400]A;VARTYPE=BND:DUP-th;JOINTYPE=th
