chr12	96010456	+	chr12	96012415	+	.	73	52	7800667_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCC;MAPQ=43;MATEID=7800667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95991001_96016001_272C;SPAN=1959;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:22 GQ:27 PL:[297.0, 27.0, 0.0] SR:52 DR:73 LR:-297.1 LO:297.1);ALT=C[chr12:96012415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96340355	+	chr12	96342955	+	.	86	60	7801392_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAGACTGC;MAPQ=60;MATEID=7801392_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96334001_96359001_33C;SPAN=2600;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:126 DP:47 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:60 DR:86 LR:-373.0 LO:373.0);ALT=C[chr12:96342955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
