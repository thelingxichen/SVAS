chr7	157275641	+	chr7	157273983	+	.	109	0	3704548_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=3704548_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:157273983(-)-7:157275641(+)__7_157265501_157290501D;SPAN=1658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:60 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:0 DR:109 LR:-323.5 LO:323.5);ALT=]chr7:157275641]C;VARTYPE=BND:DUP-th;JOINTYPE=th
