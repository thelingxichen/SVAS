chr5	148891437	+	chr5	148892633	+	.	2	5	2610003_1	3.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2610003_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_148886501_148911501_186C;SPAN=1196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:59 GQ:3.8 PL:[3.8, 0.0, 139.1] SR:5 DR:2 LR:-3.821 LO:11.68);ALT=T[chr5:148892633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	148922271	+	chr13	33229519	+	.	2	18	5447274_1	59.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTT;MAPQ=60;MATEID=5447274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_33222001_33247001_298C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:16 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:18 DR:2 LR:-59.41 LO:59.41);ALT=T[chr13:33229519[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	149460576	+	chr5	149466022	+	.	8	0	2611474_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2611474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149460576(+)-5:149466022(-)__5_149450001_149475001D;SPAN=5446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:0 DR:8 LR:-11.51 LO:16.91);ALT=G[chr5:149466022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149778059	+	chr5	149779370	+	.	8	0	2612128_1	10.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=2612128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149778059(+)-5:149779370(-)__5_149768501_149793501D;SPAN=1311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=C[chr5:149779370[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149781858	+	chr5	149784644	+	.	18	0	2612149_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612149_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149781858(+)-5:149784644(-)__5_149768501_149793501D;SPAN=2786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:112 GQ:29.3 PL:[29.3, 0.0, 240.5] SR:0 DR:18 LR:-29.07 LO:38.89);ALT=T[chr5:149784644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149781865	+	chr5	149784242	+	.	37	0	2612150_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612150_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149781865(+)-5:149784242(-)__5_149768501_149793501D;SPAN=2377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:123 GQ:89 PL:[89.0, 0.0, 207.8] SR:0 DR:37 LR:-88.81 LO:91.51);ALT=G[chr5:149784242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149782190	+	chr5	149784243	+	.	11	89	2612153_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2612153_2;MATENM=0;NM=0;NUMPARTS=6;REPSEQ=TCTC;SCTG=c_5_149768501_149793501_67C;SPAN=2053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:98 DP:201 GQ:99 PL:[269.3, 0.0, 216.5] SR:89 DR:11 LR:-269.3 LO:269.3);ALT=T[chr5:149784243[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149782234	+	chr5	149784644	+	.	25	0	2612154_1	54.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2612154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149782234(+)-5:149784644(-)__5_149768501_149793501D;SPAN=2410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:104 GQ:54.5 PL:[54.5, 0.0, 196.4] SR:0 DR:25 LR:-54.35 LO:58.94);ALT=C[chr5:149784644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149782238	+	chr5	149785821	+	.	19	0	2612155_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149782238(+)-5:149785821(-)__5_149768501_149793501D;SPAN=3583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:164 GQ:18.4 PL:[18.4, 0.0, 378.2] SR:0 DR:19 LR:-18.29 LO:38.13);ALT=A[chr5:149785821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149782916	+	chr5	149784644	+	.	9	0	2612159_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612159_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149782916(+)-5:149784644(-)__5_149768501_149793501D;SPAN=1728;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:106 GQ:1.1 PL:[1.1, 0.0, 255.2] SR:0 DR:9 LR:-0.991 LO:16.78);ALT=G[chr5:149784644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149784370	+	chr5	149786443	+	.	10	0	2612164_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612164_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149784370(+)-5:149786443(-)__5_149768501_149793501D;SPAN=2073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:157 GQ:9.4 PL:[0.0, 9.4, 399.3] SR:0 DR:10 LR:9.525 LO:17.35);ALT=C[chr5:149786443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149784372	+	chr5	149785821	+	.	27	0	2612165_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612165_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149784372(+)-5:149785821(-)__5_149768501_149793501D;SPAN=1449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:164 GQ:44.9 PL:[44.9, 0.0, 351.8] SR:0 DR:27 LR:-44.7 LO:58.65);ALT=C[chr5:149785821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149784745	+	chr5	149785822	+	.	11	73	2612166_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2612166_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_5_149768501_149793501_67C;SPAN=1077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:252 GQ:99 PL:[205.9, 0.0, 404.0] SR:73 DR:11 LR:-205.7 LO:209.3);ALT=T[chr5:149785822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149784792	+	chr5	149786753	+	.	22	0	2612168_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612168_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149784792(+)-5:149786753(-)__5_149768501_149793501D;SPAN=1961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:22 DP:1130 GQ:99 PL:[0.0, 233.3, 3212.0] SR:0 DR:22 LR:233.5 LO:26.75);ALT=A[chr5:149786753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149785937	+	chr5	149792248	+	.	25	0	2612176_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2612176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:149785937(+)-5:149792248(-)__5_149768501_149793501D;SPAN=6311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:25 DP:733 GQ:99 PL:[0.0, 115.7, 2010.0] SR:0 DR:25 LR:116.1 LO:36.47);ALT=T[chr5:149792248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149786889	+	chr5	149792188	+	.	295	45	2612182_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2612182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_149768501_149793501_50C;SPAN=5299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:303 DP:847 GQ:99 PL:[770.9, 0.0, 1286.0] SR:45 DR:295 LR:-770.7 LO:777.8);ALT=T[chr5:149792188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	149827299	+	chr5	149829049	+	.	0	8	2611945_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2611945_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_149817501_149842501_159C;SPAN=1750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:8 DR:0 LR:0.6845 LO:14.7);ALT=C[chr5:149829049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150073804	+	chr5	150075068	+	.	0	10	2612308_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2612308_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150062501_150087501_151C;SPAN=1264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:10 DR:0 LR:-20.01 LO:22.86);ALT=T[chr5:150075068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150078243	+	chr5	150080493	+	.	19	0	2612319_1	46.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2612319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150078243(+)-5:150080493(-)__5_150062501_150087501D;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:61 GQ:46.4 PL:[46.4, 0.0, 99.2] SR:0 DR:19 LR:-46.19 LO:47.34);ALT=A[chr5:150080493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150133221	+	chr5	150135979	+	.	0	12	2612605_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2612605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150111501_150136501_135C;SPAN=2758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:72 GQ:20.3 PL:[20.3, 0.0, 152.3] SR:12 DR:0 LR:-20.11 LO:26.14);ALT=T[chr5:150135979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150136051	+	chr5	150138419	+	.	16	11	2612612_1	56.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=2612612_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150111501_150136501_10C;SPAN=2368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:36 GQ:29.9 PL:[56.3, 0.0, 29.9] SR:11 DR:16 LR:-56.66 LO:56.66);ALT=T[chr5:150138419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150158534	+	chr5	150174991	+	.	109	93	2612487_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2612487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150160501_150185501_283C;SPAN=16457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:55 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:93 DR:109 LR:-435.7 LO:435.7);ALT=G[chr5:150174991[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150415309	+	chr5	150418656	+	.	8	0	2612841_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612841_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150415309(+)-5:150418656(-)__5_150405501_150430501D;SPAN=3347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=C[chr5:150418656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150416484	+	chr5	150422101	+	TGTTGAGCCGCTGGATCTCCTTTTCCTGGTACTCACGCTGTCGGGTGAGTGGGCTCAGCTGATCCTGCAGGTACTTGACCTTTTGGCGCAGCTCCTTGGCCTCTGCTGTCAGCTGCTCCTTGTCGGT	0	12	2612844_1	21.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGTTGAGCCGCTGGATCTCCTTTTCCTGGTACTCACGCTGTCGGGTGAGTGGGCTCAGCTGATCCTGCAGGTACTTGACCTTTTGGCGCAGCTCCTTGGCCTCTGCTGTCAGCTGCTCCTTGTCGGT;MAPQ=60;MATEID=2612844_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_150405501_150430501_53C;SPAN=5617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:12 DR:0 LR:-21.19 LO:26.47);ALT=T[chr5:150422101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150444740	+	chr5	150460497	+	.	35	0	2612869_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612869_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150444740(+)-5:150460497(-)__5_150454501_150479501D;SPAN=15757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:18 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:35 LR:-102.3 LO:102.3);ALT=G[chr5:150460497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150481070	+	chr5	150483130	+	.	3	4	2612912_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2612912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150479001_150504001_296C;SPAN=2060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:58 GQ:7.4 PL:[7.4, 0.0, 132.8] SR:4 DR:3 LR:-7.393 LO:14.18);ALT=T[chr5:150483130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150497399	+	chr5	150501707	+	CTCCTTATAGGCCTCATTGATGGCCCGGATTTCAGCATTGGTCCGAGTGGCCAGGATTTCAATAAGAGCCTTTTCATCTGTGCCGGCTC	3	14	2612940_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTCCTTATAGGCCTCATTGATGGCCCGGATTTCAGCATTGGTCCGAGTGGCCAGGATTTCAATAAGAGCCTTTTCATCTGTGCCGGCTC;MAPQ=60;MATEID=2612940_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_150479001_150504001_115C;SPAN=4308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:66 GQ:35 PL:[35.0, 0.0, 124.1] SR:14 DR:3 LR:-34.94 LO:37.79);ALT=C[chr5:150501707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150515921	+	chr5	150518237	+	.	8	0	2612991_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2612991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150515921(+)-5:150518237(-)__5_150503501_150528501D;SPAN=2316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=G[chr5:150518237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150516883	+	chr5	150518238	+	.	0	6	2612994_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2612994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_150503501_150528501_134C;SPAN=1355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:57 GQ:4.4 PL:[4.4, 0.0, 133.1] SR:6 DR:0 LR:-4.363 LO:11.78);ALT=C[chr5:150518238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150518402	+	chr5	150537239	+	.	9	0	2613202_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2613202_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150518402(+)-5:150537239(-)__5_150528001_150553001D;SPAN=18837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=T[chr5:150537239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150519064	+	chr5	150537239	+	.	29	0	2613203_1	95.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2613203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150519064(+)-5:150537239(-)__5_150528001_150553001D;SPAN=18175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:33 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:0 DR:29 LR:-94.28 LO:94.28);ALT=C[chr5:150537239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150519863	+	chr5	150537236	+	.	54	0	2613206_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2613206_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:150519863(+)-5:150537236(-)__5_150528001_150553001D;SPAN=17373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:32 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=C[chr5:150537236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	150632858	+	chr5	150639314	+	.	6	2	2613064_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2613064_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_150626001_150651001_259C;SPAN=6456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:2 DR:6 LR:-10.37 LO:14.87);ALT=G[chr5:150639314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151122522	+	chr5	151125839	+	.	13	99	2613974_1	99.0	.	DISC_MAPQ=37;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2613974_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CCCCC;SCTG=c_5_151116001_151141001_228C;SPAN=3317;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:130 GQ:14.1 PL:[308.9, 14.1, 0.0] SR:99 DR:13 LR:-318.4 LO:318.4);ALT=T[chr5:151125839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151122522	+	chr5	151138107	+	GCCCCCTTTGGTCCATCCTGTGGGCTGTGGGGACCAGGCCCCTGCTACTCAAGGCCAAGGTAGGAAACAGTCTTTCCTGTTTTCTTCAGGGTTGCAAGCAGAGTGTCCATGCTGTGCTCAGATTCAATGCAGACCTTCTTGTTGGGCAGGTCAATGTCATACTTAACTCCTCCAAGCTTATTGAGGACCCGAGAGACAGCTTCAGCACAGCCTCCACAGGTCATGTCCACAGAGAACTCGTGCTT	11	127	2613975_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GCCCCCTTTGGTCCATCCTGTGGGCTGTGGGGACCAGGCCCCTGCTACTCAAGGCCAAGGTAGGAAACAGTCTTTCCTGTTTTCTTCAGGGTTGCAAGCAGAGTGTCCATGCTGTGCTCAGATTCAATGCAGACCTTCTTGTTGGGCAGGTCAATGTCATACTTAACTCCTCCAAGCTTATTGAGGACCCGAGAGACAGCTTCAGCACAGCCTCCACAGGTCATGTCCACAGAGAACTCGTGCTT;MAPQ=60;MATEID=2613975_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_151116001_151141001_228C;SPAN=15585;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:111 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:127 DR:11 LR:-382.9 LO:382.9);ALT=T[chr5:151138107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151126012	+	chr5	151131264	+	.	5	40	2613985_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2613985_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_151116001_151141001_228C;SPAN=5252;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:94 GQ:99 PL:[123.2, 0.0, 103.4] SR:40 DR:5 LR:-123.2 LO:123.2);ALT=T[chr5:151131264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151126059	+	chr5	151138106	+	.	76	0	2613986_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2613986_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:151126059(+)-5:151138106(-)__5_151116001_151141001D;SPAN=12047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:86 GQ:19.8 PL:[247.5, 19.8, 0.0] SR:0 DR:76 LR:-247.8 LO:247.8);ALT=C[chr5:151138106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151131341	+	chr5	151138107	+	.	14	12	2614009_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2614009_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_151116001_151141001_228C;SPAN=6766;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:89 GQ:48.5 PL:[48.5, 0.0, 167.3] SR:12 DR:14 LR:-48.51 LO:52.18);ALT=C[chr5:151138107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151151600	+	chr5	151166144	+	.	12	0	2614113_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2614113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:151151600(+)-5:151166144(-)__5_151165001_151190001D;SPAN=14544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:25 GQ:26.3 PL:[32.9, 0.0, 26.3] SR:0 DR:12 LR:-32.86 LO:32.86);ALT=A[chr5:151166144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	151456430	+	chr5	151462448	+	.	35	24	2614687_1	88.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAAAATTACATGGTGGA;MAPQ=60;MATEID=2614687_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_5_151459001_151484001_126C;SPAN=6018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:234 GQ:88.6 PL:[88.6, 0.0, 478.1] SR:24 DR:35 LR:-88.45 LO:103.9);ALT=A[chr5:151462448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	33000094	+	chr13	33002040	+	.	0	16	5446680_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5446680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_32977001_33002001_47C;SPAN=1946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:63 GQ:35.9 PL:[35.9, 0.0, 115.1] SR:16 DR:0 LR:-35.75 LO:38.17);ALT=T[chr13:33002040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	33092140	+	chr13	33095509	+	.	2	6	5446829_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5446829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_33075001_33100001_334C;SPAN=3369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:81 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:6 DR:2 LR:-1.162 LO:13.11);ALT=C[chr13:33095509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	33101671	+	chr13	33112778	+	.	13	0	5446945_1	15.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5446945_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:33101671(+)-13:33112778(-)__13_33099501_33124501D;SPAN=11107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:0 DR:13 LR:-15.01 LO:26.61);ALT=T[chr13:33112778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	33111166	+	chr13	33112755	+	.	98	20	5446976_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5446976_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_33099501_33124501_236C;SPAN=1589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:106 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:20 DR:98 LR:-313.6 LO:313.6);ALT=T[chr13:33112755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	33223017	+	chr13	33225939	+	.	3	3	5447288_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5447288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_33222001_33247001_216C;SPAN=2922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:3 DR:3 LR:6.574 LO:6.671);ALT=G[chr13:33225939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
