chr6	64282624	+	chr6	64286341	+	.	54	56	2878902_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=2878902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_64263501_64288501_311C;SPAN=3717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:128 GQ:64.4 PL:[245.9, 0.0, 64.4] SR:56 DR:54 LR:-251.8 LO:251.8);ALT=T[chr6:64286341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	64346055	+	chr6	64389900	+	.	3	3	2879270_1	3.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2879270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_64386001_64411001_337C;SPAN=43845;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:3 DR:3 LR:-3.23 LO:9.742);ALT=G[chr6:64389900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	64667011	+	chr6	64668347	+	.	42	40	2879964_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGAA;MAPQ=60;MATEID=2879964_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_64655501_64680501_276C;SPAN=1336;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:76 GQ:7.2 PL:[198.0, 7.2, 0.0] SR:40 DR:42 LR:-204.2 LO:204.2);ALT=A[chr6:64668347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
