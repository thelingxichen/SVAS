chr7	97769422	+	chr7	31183924	+	.	14	8	5068681_1	62.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTTTCTTTCTTTCTTTCTTTCTTTCTTTC;MAPQ=34;MATEID=5068681_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_7_97755001_97780001_124C;SPAN=66585498;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:36 GQ:23.3 PL:[62.9, 0.0, 23.3] SR:8 DR:14 LR:-63.79 LO:63.79);ALT=]chr7:97769422]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	96475901	+	chr7	96481995	+	.	125	45	5062924_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCAACTGGAACTTTC;MAPQ=60;MATEID=5062924_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_96456501_96481501_314C;SPAN=6094;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:146 DP:18 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:45 DR:125 LR:-432.4 LO:432.4);ALT=C[chr7:96481995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	97420483	+	chr7	97402640	+	.	29	57	5066663_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCCT;MAPQ=60;MATEID=5066663_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_97387501_97412501_320C;SPAN=17843;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:41 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:57 DR:29 LR:-221.2 LO:221.2);ALT=]chr7:97420483]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	98381952	-	chr7	98383249	+	.	3	2	5071682_1	0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CCTCGGCCTCCCA;MAPQ=56;MATEID=5071682_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98367501_98392501_391C;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:183 GQ:36.1 PL:[0.0, 36.1, 514.9] SR:2 DR:3 LR:36.38 LO:5.063);ALT=[chr7:98383249[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
