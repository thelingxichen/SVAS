chr1	81404772	+	chr1	81410949	+	.	61	20	218433_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AAAGTCTCACTTCTT;MAPQ=60;MATEID=218433_2;MATENM=1;NM=22;NUMPARTS=2;SCTG=c_1_81389001_81414001_235C;SPAN=6177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:522 GQ:99 PL:[162.5, 0.0, 1103.0] SR:20 DR:61 LR:-162.3 LO:202.9);ALT=T[chr1:81410949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	81660351	+	chr1	81661558	-	.	40	58	218365_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=218365_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_81658501_81683501_166C;SPAN=1207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:58 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:58 DR:40 LR:-254.2 LO:254.2);ALT=T]chr1:81661558];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	81660357	-	chr1	81661371	+	ATTTTAAATTATTAAAAAA	26	42	218366_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTTTAAATTATTAAAAAA;MAPQ=60;MATEID=218366_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_81658501_81683501_91C;SPAN=1014;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:56 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:42 DR:26 LR:-168.3 LO:168.3);ALT=[chr1:81661371[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
