chr4	167677048	+	chr4	167683072	+	.	94	37	3053022_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAGAGATTTGGG;MAPQ=60;MATEID=3053022_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_167678001_167703001_38C;SPAN=6024;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:122 DP:28 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:37 DR:94 LR:-359.8 LO:359.8);ALT=G[chr4:167683072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	168371943	+	chr4	168373137	+	.	45	34	3054945_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAT;MAPQ=60;MATEID=3054945_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_168364001_168389001_43C;SPAN=1194;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:60 GQ:18 PL:[198.0, 18.0, 0.0] SR:34 DR:45 LR:-198.0 LO:198.0);ALT=T[chr4:168373137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	169116816	+	chr4	169118418	+	.	76	59	3057982_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCA;MAPQ=60;MATEID=3057982_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_169099001_169124001_322C;SPAN=1602;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:84 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:59 DR:76 LR:-333.4 LO:333.4);ALT=A[chr4:169118418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	169979191	+	chr4	169980310	-	.	8	0	3061879_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3061879_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:169979191(+)-4:169980310(+)__4_169956501_169981501D;SPAN=1119;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:146 GQ:12.9 PL:[0.0, 12.9, 379.5] SR:0 DR:8 LR:13.15 LO:13.34);ALT=G]chr4:169980310];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	170445446	-	chr4	170446453	+	.	7	2	3063685_1	0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TCTCTACTAAAAATA;MAPQ=15;MATEID=3063685_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_170422001_170447001_43C;SPAN=1007;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:132 GQ:9 PL:[0.0, 9.0, 336.6] SR:2 DR:7 LR:9.354 LO:13.7);ALT=[chr4:170446453[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	171240407	-	chr4	171282328	+	.	10	0	3067148_1	13.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=3067148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:171240407(-)-4:171282328(-)__4_171279501_171304501D;SPAN=41921;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:73 GQ:13.4 PL:[13.4, 0.0, 161.9] SR:0 DR:10 LR:-13.23 LO:20.85);ALT=[chr4:171282328[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	171866752	+	chr4	171855225	+	.	64	74	3068917_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3068917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_171843001_171868001_160C;SPAN=11527;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:109 DP:150 GQ:45.2 PL:[319.1, 0.0, 45.2] SR:74 DR:64 LR:-331.1 LO:331.1);ALT=]chr4:171866752]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	172374412	+	chr4	172379426	+	.	108	85	3070662_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3070662_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_4_172357501_172382501_56C;SPAN=5014;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:165 DP:35 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:85 DR:108 LR:-488.5 LO:488.5);ALT=G[chr4:172379426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	172988639	+	chr4	172992932	+	C	56	42	3072695_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=3072695_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_172970001_172995001_232C;SPAN=4293;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:82 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:42 DR:56 LR:-241.0 LO:241.0);ALT=A[chr4:172992932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	173425032	+	chr4	173433521	+	A	141	103	3074291_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=3074291_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_173411001_173436001_50C;SPAN=8489;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:186 DP:38 GQ:50.2 PL:[551.2, 50.2, 0.0] SR:103 DR:141 LR:-551.2 LO:551.2);ALT=A[chr4:173433521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
