chr16	86379235	-	chr16	86385544	+	.	8	0	9449259_1	0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=9449259_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:86379235(-)-16:86385544(-)__16_86362501_86387501D;SPAN=6309;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:0 DR:8 LR:3.123 LO:14.39);ALT=[chr16:86385544[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
