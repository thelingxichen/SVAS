chr4	48712716	+	chr4	48782095	+	.	6	7	1959443_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1959443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_48706001_48731001_36C;SPAN=69379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:30 GQ:31.4 PL:[31.4, 0.0, 41.3] SR:7 DR:6 LR:-31.48 LO:31.56);ALT=C[chr4:48782095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48833416	+	chr4	48834636	+	.	28	3	1959383_1	80.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1959383_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_48828501_48853501_64C;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:70 GQ:80 PL:[80.0, 0.0, 89.9] SR:3 DR:28 LR:-80.07 LO:80.1);ALT=G[chr4:48834636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48833442	+	chr4	48835415	+	.	30	0	1959384_1	82.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1959384_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:48833442(+)-4:48835415(-)__4_48828501_48853501D;SPAN=1973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:62 GQ:65.9 PL:[82.4, 0.0, 65.9] SR:0 DR:30 LR:-82.3 LO:82.3);ALT=T[chr4:48835415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48834699	+	chr4	48851964	+	ACATAGGGCCTGATTACATTCCAACAGAGGAAGAAAGGAGAGTCTTCGCAGAATGCAATGATGAAAGCTTCTGGTTCAGATCTGTGCCTTTGGCTGCAACAAGTATGTTGATTACTCAAGGATTAATTAGTAAAGGAATACTTTCAAGTCATCCCAAATATGGTTCCATCCCTAAACTTATAC	0	47	1959388_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ACATAGGGCCTGATTACATTCCAACAGAGGAAGAAAGGAGAGTCTTCGCAGAATGCAATGATGAAAGCTTCTGGTTCAGATCTGTGCCTTTGGCTGCAACAAGTATGTTGATTACTCAAGGATTAATTAGTAAAGGAATACTTTCAAGTCATCCCAAATATGGTTCCATCCCTAAACTTATAC;MAPQ=60;MATEID=1959388_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_4_48828501_48853501_43C;SPAN=17265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:55 GQ:8.1 PL:[148.5, 8.1, 0.0] SR:47 DR:0 LR:-150.8 LO:150.8);ALT=C[chr4:48851964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48853993	+	chr4	48859228	+	.	9	8	1959503_1	28.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1959503_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_48853001_48878001_93C;SPAN=5235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:8 DR:9 LR:-28.55 LO:30.78);ALT=G[chr4:48859228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48859382	+	chr4	48862740	+	.	5	3	1959506_1	10.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1959506_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_48853001_48878001_203C;SPAN=3358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:46 GQ:10.7 PL:[10.7, 0.0, 99.8] SR:3 DR:5 LR:-10.64 LO:14.94);ALT=G[chr4:48862740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48901945	+	chr4	48908675	+	CTTGCTTGGTGGTGGAAAATGGGCATCTTTATCTTGGTTTCCACGAGCAGACGCTGAAGCCATGATGACTTTGTGCTTGCTCTCCTTCCAGTTGTTTATCCTCTGCTTACTCCTTGACCCAGTGT	15	45	1959585_1	99.0	.	DISC_MAPQ=37;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTTGCTTGGTGGTGGAAAATGGGCATCTTTATCTTGGTTTCCACGAGCAGACGCTGAAGCCATGATGACTTTGTGCTTGCTCTCCTTCCAGTTGTTTATCCTCTGCTTACTCCTTGACCCAGTGT;MAPQ=60;MATEID=1959585_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_48877501_48902501_42C;SPAN=6730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:28 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:45 DR:15 LR:-148.5 LO:148.5);ALT=G[chr4:48908675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	48906630	+	chr4	48908675	+	.	49	12	1959741_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1959741_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_4_48902001_48927001_219C;SPAN=2045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:57 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:12 DR:49 LR:-168.3 LO:168.3);ALT=T[chr4:48908675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	49150380	+	chr4	49149163	+	.	9	0	1962699_1	0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=1962699_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:49149163(-)-4:49150380(+)__4_49147001_49172001D;SPAN=1217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:115 GQ:1.2 PL:[0.0, 1.2, 280.5] SR:0 DR:9 LR:1.447 LO:16.45);ALT=]chr4:49150380]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	49637128	+	chr4	49635891	+	.	14	0	1964122_1	24.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=1964122_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:49635891(-)-4:49637128(+)__4_49612501_49637501D;SPAN=1237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:82 GQ:24.2 PL:[24.2, 0.0, 172.7] SR:0 DR:14 LR:-24.0 LO:30.65);ALT=]chr4:49637128]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	49659869	+	chr4	49658836	+	.	16	0	1967152_1	13.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=1967152_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:49658836(-)-4:49659869(+)__4_49637001_49662001D;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:147 GQ:13.1 PL:[13.1, 0.0, 343.1] SR:0 DR:16 LR:-12.99 LO:31.65);ALT=]chr4:49659869]T;VARTYPE=BND:DUP-th;JOINTYPE=th
