chr21	33032155	+	chr21	33039569	+	AAAGTAATGGACCAGTGAAGGTGTGGGGAAGCATTAAAGGACTGACTGAAGGCCTGCATGGATTCCATGTTCATGAGTTTGGAGATAATACAGCAGGCTGTACCAGTGCAGGTCCTCACTTTAATCCTCTATCCAGAAAACACGGTGGGCCAAAGGATGAAGAG	0	159	7157607_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAAGTAATGGACCAGTGAAGGTGTGGGGAAGCATTAAAGGACTGACTGAAGGCCTGCATGGATTCCATGTTCATGAGTTTGGAGATAATACAGCAGGCTGTACCAGTGCAGGTCCTCACTTTAATCCTCTATCCAGAAAACACGGTGGGCCAAAGGATGAAGAG;MAPQ=60;MATEID=7157607_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_21_33026001_33051001_61C;SPAN=7414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:159 DP:116 GQ:43 PL:[472.0, 43.0, 0.0] SR:159 DR:0 LR:-472.0 LO:472.0);ALT=G[chr21:33039569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33032155	+	chr21	33036100	+	.	75	85	7157606_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AAGG;MAPQ=60;MATEID=7157606_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_21_33026001_33051001_61C;SPAN=3945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:121 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:85 DR:75 LR:-382.9 LO:382.9);ALT=G[chr21:33036100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33032165	+	chr21	33038758	+	.	31	0	7157608_1	75.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7157608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:33032165(+)-21:33038758(-)__21_33026001_33051001D;SPAN=6593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:101 GQ:75.2 PL:[75.2, 0.0, 167.6] SR:0 DR:31 LR:-74.97 LO:77.0);ALT=G[chr21:33038758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33039690	+	chr21	33040783	+	.	7	93	7157627_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=7157627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_33026001_33051001_87C;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:118 GQ:5.4 PL:[297.0, 5.4, 0.0] SR:93 DR:7 LR:-310.9 LO:310.9);ALT=T[chr21:33040783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33253902	+	chr21	33250497	+	.	37	0	7158278_1	91.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7158278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:33250497(-)-21:33253902(+)__21_33246501_33271501D;SPAN=3405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:114 GQ:91.4 PL:[91.4, 0.0, 183.8] SR:0 DR:37 LR:-91.25 LO:93.01);ALT=]chr21:33253902]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	33976595	+	chr21	33979959	+	.	3	3	7160410_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=7160410_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_33957001_33982001_228C;SPAN=3364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:70 GQ:0.8 PL:[0.8, 0.0, 169.1] SR:3 DR:3 LR:-0.8413 LO:11.21);ALT=T[chr21:33979959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33980028	+	chr21	33982148	+	.	0	7	7160418_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7160418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_33957001_33982001_4C;SPAN=2120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:35 GQ:13.7 PL:[13.7, 0.0, 69.8] SR:7 DR:0 LR:-13.62 LO:15.86);ALT=T[chr21:33982148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	33982317	+	chr21	33984415	+	.	0	11	7160499_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7160499_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_33981501_34006501_74C;SPAN=2098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:11 DR:0 LR:-8.677 LO:21.71);ALT=T[chr21:33984415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34633032	+	chr21	34634865	+	.	0	18	7162152_1	35.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7162152_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34618501_34643501_260C;SPAN=1833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:18 DR:0 LR:-35.58 LO:40.99);ALT=G[chr21:34634865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34638819	+	chr21	34640697	+	.	16	2	7162176_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7162176_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34618501_34643501_108C;SPAN=1878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:84 GQ:33.5 PL:[33.5, 0.0, 168.8] SR:2 DR:16 LR:-33.36 LO:38.63);ALT=G[chr21:34640697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34697368	+	chr21	34707827	+	.	10	0	7162483_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7162483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:34697368(+)-21:34707827(-)__21_34692001_34717001D;SPAN=10459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:0 DR:10 LR:-8.085 LO:19.77);ALT=T[chr21:34707827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34775922	+	chr21	34787193	+	.	0	36	7162677_1	94.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7162677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34765501_34790501_74C;SPAN=11271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:92 GQ:94.1 PL:[94.1, 0.0, 127.1] SR:36 DR:0 LR:-93.91 LO:94.22);ALT=G[chr21:34787193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34787327	+	chr21	34793787	+	.	0	11	7162709_1	25.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7162709_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34765501_34790501_65C;SPAN=6460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:42 GQ:25.1 PL:[25.1, 0.0, 74.6] SR:11 DR:0 LR:-24.93 LO:26.41);ALT=A[chr21:34793787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34839430	+	chr21	34841094	+	.	0	16	7163086_1	26.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7163086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34839001_34864001_106C;SPAN=1664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:98 GQ:26.3 PL:[26.3, 0.0, 211.1] SR:16 DR:0 LR:-26.27 LO:34.69);ALT=C[chr21:34841094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34841231	+	chr21	34852143	+	.	19	0	7163096_1	43.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7163096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:34841231(+)-21:34852143(-)__21_34839001_34864001D;SPAN=10912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:71 GQ:43.7 PL:[43.7, 0.0, 126.2] SR:0 DR:19 LR:-43.48 LO:45.84);ALT=A[chr21:34852143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34907672	+	chr21	34914367	+	.	8	0	7163050_1	16.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7163050_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:34907672(+)-21:34914367(-)__21_34888001_34913001D;SPAN=6695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=C[chr21:34914367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34915475	+	chr21	34918517	+	.	66	21	7162925_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7162925_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34912501_34937501_10C;SPAN=3042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:98 GQ:6.5 PL:[230.9, 0.0, 6.5] SR:21 DR:66 LR:-243.7 LO:243.7);ALT=G[chr21:34918517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34918685	+	chr21	34921780	+	.	0	44	7162934_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7162934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34912501_34937501_203C;SPAN=3095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:104 GQ:99 PL:[117.2, 0.0, 133.7] SR:44 DR:0 LR:-117.1 LO:117.1);ALT=G[chr21:34921780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34994376	+	chr21	34996989	+	.	0	25	7163704_1	61.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7163704_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_34986001_35011001_309C;SPAN=2613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:78 GQ:61.4 PL:[61.4, 0.0, 127.4] SR:25 DR:0 LR:-61.39 LO:62.68);ALT=T[chr21:34996989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34994421	+	chr21	35013982	+	.	15	0	7163705_1	41.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7163705_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:34994421(+)-21:35013982(-)__21_34986001_35011001D;SPAN=19561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:29 GQ:28.4 PL:[41.6, 0.0, 28.4] SR:0 DR:15 LR:-41.78 LO:41.78);ALT=C[chr21:35013982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	34997110	+	chr21	35013986	+	.	10	0	7163715_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7163715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:34997110(+)-21:35013986(-)__21_34986001_35011001D;SPAN=16876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:34 GQ:23.9 PL:[23.9, 0.0, 56.9] SR:0 DR:10 LR:-23.8 LO:24.62);ALT=C[chr21:35013986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35276325	+	chr21	35279645	+	.	0	46	7164391_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7164391_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_35255501_35280501_188C;SPAN=3320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:92 GQ:94.1 PL:[127.1, 0.0, 94.1] SR:46 DR:0 LR:-127.1 LO:127.1);ALT=G[chr21:35279645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35279757	+	chr21	35281394	+	TGATCAGG	0	46	7164570_1	99.0	.	EVDNC=ASSMB;INSERTION=TGATCAGG;MAPQ=60;MATEID=7164570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_35280001_35305001_180C;SPAN=1637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:53 GQ:10.8 PL:[148.5, 10.8, 0.0] SR:46 DR:0 LR:-148.7 LO:148.7);ALT=T[chr21:35281394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35279809	+	chr21	35288028	+	.	12	0	7164572_1	15.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7164572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:35279809(+)-21:35288028(-)__21_35280001_35305001D;SPAN=8219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:88 GQ:15.8 PL:[15.8, 0.0, 197.3] SR:0 DR:12 LR:-15.77 LO:24.99);ALT=T[chr21:35288028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35281515	+	chr21	35288029	+	TGCTACTCTCAACAACTCCTTTTCTACTTGCTCCAGCTTATTCTGTTTTGATGCAGCAGAATAAAGAGCTGTGGCATAGCGACCTTCAATACCGTATACCTGAACAGGAGGCCTCACAAGCTTGGCAAATGGTCTGACCACAGAGGTACTGAAGCATCG	96	108	7164584_1	99.0	.	DISC_MAPQ=47;EVDNC=TSI_G;HOMSEQ=CACCT;INSERTION=TGCTACTCTCAACAACTCCTTTTCTACTTGCTCCAGCTTATTCTGTTTTGATGCAGCAGAATAAAGAGCTGTGGCATAGCGACCTTCAATACCGTATACCTGAACAGGAGGCCTCACAAGCTTGGCAAATGGTCTGACCACAGAGGTACTGAAGCATCG;MAPQ=60;MATEID=7164584_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_21_35280001_35305001_91C;SPAN=6514;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:164 DP:148 GQ:44.2 PL:[485.2, 44.2, 0.0] SR:108 DR:96 LR:-485.2 LO:485.2);ALT=G[chr21:35288029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35281515	+	chr21	35284593	+	.	4	94	7164583_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=7164583_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_21_35280001_35305001_91C;SPAN=3078;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:113 GQ:20.4 PL:[313.5, 20.4, 0.0] SR:94 DR:4 LR:-316.6 LO:316.6);ALT=G[chr21:35284593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35284748	+	chr21	35288025	+	.	125	0	7164592_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7164592_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:35284748(+)-21:35288025(-)__21_35280001_35305001D;SPAN=3277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:103 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:0 DR:125 LR:-369.7 LO:369.7);ALT=C[chr21:35288025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35286806	+	chr21	35288029	+	.	14	12	7164600_1	19.0	.	DISC_MAPQ=18;EVDNC=TSI_L;HOMSEQ=CACCT;MAPQ=60;MATEID=7164600_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_21_35280001_35305001_91C;SPAN=1223;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:137 GQ:19.1 PL:[19.1, 0.0, 312.8] SR:12 DR:14 LR:-19.0 LO:34.66);ALT=T[chr21:35288029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35446022	+	chr21	35514706	+	.	10	0	7165007_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7165007_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:35446022(+)-21:35514706(-)__21_35500501_35525501D;SPAN=68684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:0 DR:10 LR:-20.28 LO:22.97);ALT=T[chr21:35514706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35446045	+	chr21	35497640	+	.	0	39	7164781_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7164781_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_35476001_35501001_134C;SPAN=51595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:39 DR:0 LR:-115.5 LO:115.5);ALT=G[chr21:35497640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35747911	+	chr21	35757770	+	.	19	0	7165672_1	42.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7165672_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:35747911(+)-21:35757770(-)__21_35745501_35770501D;SPAN=9859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:75 GQ:42.5 PL:[42.5, 0.0, 138.2] SR:0 DR:19 LR:-42.4 LO:45.3);ALT=A[chr21:35757770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	35751817	+	chr21	35757772	+	.	4	15	7165680_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTTC;MAPQ=60;MATEID=7165680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_35745501_35770501_330C;SPAN=5955;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:70 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:15 DR:4 LR:-37.15 LO:40.17);ALT=T[chr21:35757772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
