chr4	156588571	+	chr4	156617908	+	.	0	8	2287707_1	10.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2287707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_156604001_156629001_275C;SPAN=29337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:8 DR:0 LR:-9.882 LO:16.52);ALT=A[chr4:156617908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	156588933	+	chr4	156617905	+	.	13	0	2287708_1	26.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2287708_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:156588933(+)-4:156617905(-)__4_156604001_156629001D;SPAN=28972;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.66 LO:29.98);ALT=A[chr4:156617905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	156629447	+	chr4	156631691	+	.	0	7	2287647_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=2287647_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_156628501_156653501_231C;SPAN=2244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:7 DR:0 LR:0.4634 LO:12.88);ALT=G[chr4:156631691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
