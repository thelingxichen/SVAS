chr11	80785602	+	chr11	81093780	+	.	38	27	4935514_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGTT;MAPQ=60;MATEID=4935514_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_81070501_81095501_113C;SPAN=308178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:28 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:27 DR:38 LR:-161.7 LO:161.7);ALT=T[chr11:81093780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
