chr5	10250528	+	chr5	10254784	+	.	17	0	2413918_1	38.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2413918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:10250528(+)-5:10254784(-)__5_10241001_10266001D;SPAN=4256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:66 GQ:38.3 PL:[38.3, 0.0, 120.8] SR:0 DR:17 LR:-38.24 LO:40.68);ALT=T[chr5:10254784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10250557	+	chr5	10254255	+	.	5	16	2413919_1	36.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2413919_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_10241001_10266001_153C;SPAN=3698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:16 DR:5 LR:-36.83 LO:38.71);ALT=G[chr5:10254255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10250557	+	chr5	10256066	+	TCTCATATAATGGCAGCAAAGGCTGTAGCAAATACAATGAGAACATCACTTGGACCAAATGGGCTTGATAAGATGATGGTGGATAAGGATGGGGATGTGACTGTAACTAATGATGGGGCCACCATCTTAAGCATGATGGATGTTGATCATCAGATTGCCAAGCTGATGGTGGAACTGTCCAAGTCTCAGGATGATGAAATTGGAGATGGAACCACAGGAGTGGTT	0	26	2413920_1	71.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TCTCATATAATGGCAGCAAAGGCTGTAGCAAATACAATGAGAACATCACTTGGACCAAATGGGCTTGATAAGATGATGGTGGATAAGGATGGGGATGTGACTGTAACTAATGATGGGGCCACCATCTTAAGCATGATGGATGTTGATCATCAGATTGCCAAGCTGATGGTGGAACTGTCCAAGTCTCAGGATGATGAAATTGGAGATGGAACCACAGGAGTGGTT;MAPQ=60;MATEID=2413920_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_10241001_10266001_153C;SPAN=5509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:52 GQ:52.1 PL:[71.9, 0.0, 52.1] SR:26 DR:0 LR:-71.86 LO:71.86);ALT=G[chr5:10256066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10254950	+	chr5	10256066	+	.	4	11	2413932_1	33.0	.	DISC_MAPQ=48;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2413932_2;MATENM=0;NM=1;NUMPARTS=4;REPSEQ=CC;SCTG=c_5_10241001_10266001_153C;SPAN=1116;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:11 DR:4 LR:-33.8 LO:35.92);ALT=G[chr5:10256066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10263426	+	chr5	10264767	+	.	0	10	2413954_1	17.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=2413954_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_10241001_10266001_66C;SPAN=1341;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=G[chr5:10264767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10290895	+	chr5	10307737	+	.	6	8	2413732_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2413732_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_10290001_10315001_102C;SPAN=16842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:8 DR:6 LR:-15.72 LO:23.22);ALT=T[chr5:10307737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10354029	+	chr5	10377908	+	.	0	11	2414008_1	30.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2414008_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_10363501_10388501_238C;SPAN=23879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:20 GQ:17.6 PL:[30.8, 0.0, 17.6] SR:11 DR:0 LR:-31.09 LO:31.09);ALT=G[chr5:10377908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10415781	+	chr5	10417381	+	.	4	3	2414095_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2414095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_10412501_10437501_124C;SPAN=1600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:66 GQ:2 PL:[2.0, 0.0, 157.1] SR:3 DR:4 LR:-1.925 LO:11.37);ALT=G[chr5:10417381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10681282	+	chr5	10748287	+	CGGGCGATGACCCCAGAGATGAACACAGTGGGTTTAGGTGGA	2	9	2414530_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTGG;INSERTION=CGGGCGATGACCCCAGAGATGAACACAGTGGGTTTAGGTGGA;MAPQ=60;MATEID=2414530_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_10657501_10682501_142C;SPAN=67005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:9 DR:2 LR:-21.31 LO:22.09);ALT=C[chr5:10748287[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	10748384	+	chr5	10761126	+	.	0	20	2414693_1	57.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2414693_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_10731001_10756001_55C;SPAN=12742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:30 GQ:14.9 PL:[57.8, 0.0, 14.9] SR:20 DR:0 LR:-59.31 LO:59.31);ALT=C[chr5:10761126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
