chr5	28787996	+	chr5	28963096	+	.	36	23	2441210_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=2441210_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_28787501_28812501_165C;SPAN=175100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:19 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:23 DR:36 LR:-145.2 LO:145.2);ALT=T[chr5:28963096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
