chr3	49221838	-	chr3	49224050	+	.	8	0	2004959_1	0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2004959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:49221838(-)-3:49224050(-)__3_49220501_49245501D;SPAN=2212;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:172 GQ:19.9 PL:[0.0, 19.9, 455.5] SR:0 DR:8 LR:20.19 LO:12.76);ALT=[chr3:49224050[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	49587558	-	chr3	49589605	+	.	8	0	2007336_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2007336_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:49587558(-)-3:49589605(-)__3_49563501_49588501D;SPAN=2047;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=[chr3:49589605[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
