chr3	42838373	+	chr3	42840811	+	.	135	107	1973921_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGAATCTTATAACTTCC;MAPQ=60;MATEID=1973921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_42826001_42851001_42C;SPAN=2438;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:220 DP:41 GQ:59.5 PL:[653.5, 59.5, 0.0] SR:107 DR:135 LR:-653.6 LO:653.6);ALT=C[chr3:42840811[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
