chr8	87526780	+	chr8	87540762	+	.	35	0	3956463_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3956463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:87526780(+)-8:87540762(-)__8_87514001_87539001D;SPAN=13982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:37 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:0 DR:35 LR:-108.9 LO:108.9);ALT=G[chr8:87540762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	87544809	+	chr8	87556966	+	ATCTATTTGGAAAGTCAGACCCATACCTGGAATTCCACAAGCAGACATCTGATGGAAACTGGCTAATGGTTCATCGGACAGAGGTTGTTAAAAACAACTTGAATCCTGTTTGGAGGCCTTTCAAGATCTCTCTTAACTCACTGTGTTACGGAGATATGGACAAAACCATTA	0	16	3956364_1	31.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=ATCTATTTGGAAAGTCAGACCCATACCTGGAATTCCACAAGCAGACATCTGATGGAAACTGGCTAATGGTTCATCGGACAGAGGTTGTTAAAAACAACTTGAATCCTGTTTGGAGGCCTTTCAAGATCTCTCTTAACTCACTGTGTTACGGAGATATGGACAAAACCATTA;MAPQ=60;MATEID=3956364_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_87538501_87563501_82C;SPAN=12157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:80 GQ:31.1 PL:[31.1, 0.0, 163.1] SR:16 DR:0 LR:-31.14 LO:36.26);ALT=G[chr8:87556966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
