chr5	66481847	+	chr5	66492380	+	.	3	4	2491127_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2491127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_66468501_66493501_91C;SPAN=10533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:55 GQ:1.7 PL:[1.7, 0.0, 130.4] SR:4 DR:3 LR:-1.604 LO:9.478);ALT=T[chr5:66492380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
