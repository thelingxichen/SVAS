chrX	128914130	+	chrX	128921949	+	.	0	14	7523998_1	35.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7523998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_128919001_128944001_57C;SPAN=7819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:40 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:14 DR:0 LR:-35.38 LO:35.77);ALT=G[chrX:128921949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	129290579	+	chrX	129299524	+	.	0	10	7524675_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7524675_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_129286501_129311501_279C;SPAN=8945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:10 DR:0 LR:-15.67 LO:21.47);ALT=T[chrX:129299524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	129479250	+	chrX	129480517	+	.	2	2	7524899_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7524899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_129458001_129483001_27C;SPAN=1267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:51 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:2 DR:2 LR:0.6132 LO:7.314);ALT=G[chrX:129480517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
