chr17	10601037	+	chr17	10608235	+	.	8	0	6313001_1	1.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6313001_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:10601037(+)-17:10608235(-)__17_10584001_10609001D;SPAN=7198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:0 DR:8 LR:-0.9411 LO:14.92);ALT=G[chr17:10608235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
