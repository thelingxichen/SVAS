chr8	27456153	+	chr8	27457294	+	.	7	6	3793549_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=3793549_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_27440001_27465001_115C;SPAN=1141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:98 GQ:13.1 PL:[13.1, 0.0, 224.3] SR:6 DR:7 LR:-13.06 LO:24.39);ALT=C[chr8:27457294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27457527	+	chr8	27462441	+	CACAGACAAGATCTCCCGGCACTTGTCACACTGGTCCTTCATCCGCAGGCAGCCCGTGGAGTTGTGGCGGATCTCCCGGCACACAGTCCGGTCATCGTCGCCTT	5	10	3793555_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CACAGACAAGATCTCCCGGCACTTGTCACACTGGTCCTTCATCCGCAGGCAGCCCGTGGAGTTGTGGCGGATCTCCCGGCACACAGTCCGGTCATCGTCGCCTT;MAPQ=60;MATEID=3793555_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_8_27440001_27465001_224C;SPAN=4914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:90 GQ:25.1 PL:[25.1, 0.0, 193.4] SR:10 DR:5 LR:-25.13 LO:32.67);ALT=C[chr8:27462441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27457527	+	chr8	27461808	+	.	5	4	3793554_1	3.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3793554_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_27440001_27465001_224C;SPAN=4281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:4 DR:5 LR:-3.158 LO:17.1);ALT=C[chr8:27461808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27462856	+	chr8	27467992	+	CGGCCAACCAGGCCTGAGCCACTTCTGCAGACGCGTGCGTAGAACTTCATGCAGGTCTGTTTCAGGCAGGGCTTACACTCTTCCCAGAGGGCCATCATGGTCTCATTGCACACTCCTGGGAGCTCCTTCAGCTTTGTCTCTGATTCCCTGGTCTCATTTAGGGCATCCTCTTTCTTCTTCTTGGCTTCTTCTAGGTTGCTGAGCAGTGTCTTGCGCTCTTCGTTTGTTTTTTCTATGAGAGTCTTTATCTGTTTCACCCCGTTGACAGCATTTTGAATTTCCTTATTGACGTACTTACTTCCCTGATTGGACATTT	0	58	3793720_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CGGCCAACCAGGCCTGAGCCACTTCTGCAGACGCGTGCGTAGAACTTCATGCAGGTCTGTTTCAGGCAGGGCTTACACTCTTCCCAGAGGGCCATCATGGTCTCATTGCACACTCCTGGGAGCTCCTTCAGCTTTGTCTCTGATTCCCTGGTCTCATTTAGGGCATCCTCTTTCTTCTTCTTGGCTTCTTCTAGGTTGCTGAGCAGTGTCTTGCGCTCTTCGTTTGTTTTTTCTATGAGAGTCTTTATCTGTTTCACCCCGTTGACAGCATTTTGAATTTCCTTATTGACGTACTTACTTCCCTGATTGGACATTT;MAPQ=60;MATEID=3793720_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_27464501_27489501_34C;SPAN=5136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:69 GQ:5.4 PL:[178.2, 5.4, 0.0] SR:58 DR:0 LR:-184.9 LO:184.9);ALT=G[chr8:27467992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27462856	+	chr8	27463871	+	.	7	8	3793572_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTGG;MAPQ=60;MATEID=3793572_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_8_27440001_27465001_336C;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:127 GQ:8.6 PL:[8.6, 0.0, 299.0] SR:8 DR:7 LR:-8.506 LO:25.35);ALT=G[chr8:27463871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27464043	+	chr8	27466454	+	.	8	10	3793722_1	44.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=3793722_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TTT;SCTG=c_8_27464501_27489501_34C;SPAN=2411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:43 GQ:44.6 PL:[44.6, 0.0, 57.8] SR:10 DR:8 LR:-44.47 LO:44.59);ALT=T[chr8:27466454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27466604	+	chr8	27467992	+	.	0	43	3793729_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3793729_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_27464501_27489501_34C;SPAN=1388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:134 GQ:99 PL:[105.8, 0.0, 218.0] SR:43 DR:0 LR:-105.6 LO:107.8);ALT=C[chr8:27467992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27466645	+	chr8	27472171	+	.	43	0	3793730_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3793730_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:27466645(+)-8:27472171(-)__8_27464501_27489501D;SPAN=5526;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:123 GQ:99 PL:[108.8, 0.0, 188.0] SR:0 DR:43 LR:-108.6 LO:109.8);ALT=A[chr8:27472171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27468133	+	chr8	27472171	+	.	22	0	3793734_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3793734_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:27468133(+)-8:27472171(-)__8_27464501_27489501D;SPAN=4038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:127 GQ:38.3 PL:[38.3, 0.0, 269.3] SR:0 DR:22 LR:-38.21 LO:48.32);ALT=G[chr8:27472171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	27610149	+	chr8	27630062	+	.	10	0	3794105_1	18.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=3794105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:27610149(+)-8:27630062(-)__8_27611501_27636501D;SPAN=19913;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:54 GQ:18.5 PL:[18.5, 0.0, 110.9] SR:0 DR:10 LR:-18.38 LO:22.29);ALT=A[chr8:27630062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
