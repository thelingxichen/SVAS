chr2	162017034	+	chr2	162036122	+	.	8	0	1067012_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1067012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:162017034(+)-2:162036122(-)__2_161994001_162019001D;SPAN=19088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=C[chr2:162036122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	162165116	+	chr2	162172946	+	.	21	12	1067737_1	73.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1067737_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_162141001_162166001_93C;SPAN=7830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:45 GQ:34.1 PL:[73.7, 0.0, 34.1] SR:12 DR:21 LR:-74.35 LO:74.35);ALT=G[chr2:162172946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	162173080	+	chr2	162224295	+	AAATATGGACAGACTTCTTAGACTTGGAGGAGGTATGCCTGGACTGGGCCAGGGGCCACCTACAGATGCTCCTGCAGTGGACACAGCAGAACAAGTCTATATCTCTTCCCTGGCACTGTTAAAA	0	18	1067504_1	51.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAATATGGACAGACTTCTTAGACTTGGAGGAGGTATGCCTGGACTGGGCCAGGGGCCACCTACAGATGCTCCTGCAGTGGACACAGCAGAACAAGTCTATATCTCTTCCCTGGCACTGTTAAAA;MAPQ=60;MATEID=1067504_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_162165501_162190501_357C;SPAN=51215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:29 GQ:18.5 PL:[51.5, 0.0, 18.5] SR:18 DR:0 LR:-52.4 LO:52.4);ALT=G[chr2:162224295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	162332271	+	chr2	162334042	+	.	105	80	1067856_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GCCA;MAPQ=60;MATEID=1067856_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_162312501_162337501_27C;SPAN=1771;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:36 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:80 DR:105 LR:-429.1 LO:429.1);ALT=A[chr2:162334042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	163200785	+	chr2	163204087	+	.	28	16	1069766_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1069766_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_163194501_163219501_150C;SPAN=3302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:16 DR:28 LR:-91.97 LO:92.16);ALT=G[chr2:163204087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
