chr4	128904202	+	chr4	128905492	+	.	0	8	2200072_1	1.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2200072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_128894501_128919501_24C;SPAN=1290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:8 DR:0 LR:-0.9411 LO:14.92);ALT=G[chr4:128905492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	128982556	+	chr4	128995613	+	.	2	5	2200914_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2200914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_128992501_129017501_109C;SPAN=13057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:43 GQ:5 PL:[5.0, 0.0, 97.4] SR:5 DR:2 LR:-4.855 LO:10.04);ALT=G[chr4:128995613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
