chr18	11509708	+	chr18	11511475	+	.	77	47	9898992_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGT;MAPQ=60;MATEID=9898992_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_11490501_11515501_212C;SPAN=1767;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:95 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:47 DR:77 LR:-323.5 LO:323.5);ALT=T[chr18:11511475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12134799	+	chr18	12146288	+	.	39	72	9902565_1	99.0	.	DISC_MAPQ=29;EVDNC=ASDIS;HOMSEQ=G;MAPQ=34;MATEID=9902565_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_12127501_12152501_148C;SPAN=11489;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:101 GQ:27 PL:[297.0, 27.0, 0.0] SR:72 DR:39 LR:-294.9 LO:294.9);ALT=G[chr18:12146288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
