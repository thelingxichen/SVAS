chr8	42190455	+	chr8	42194367	+	.	64	0	5455450_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5455450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:42190455(+)-8:42194367(-)__8_42189001_42214001D;SPAN=3912;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:64 DP:14 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=G[chr8:42194367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	43097523	+	chr8	43096054	+	.	23	0	5457363_1	55.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5457363_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:43096054(-)-8:43097523(+)__8_43095501_43120501D;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:76 GQ:55.4 PL:[55.4, 0.0, 128.0] SR:0 DR:23 LR:-55.33 LO:56.96);ALT=]chr8:43097523]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	43226576	-	chr14	36674745	+	.	14	12	8442542_1	71.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=8442542_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_36652001_36677001_169C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:42 GQ:28.4 PL:[71.3, 0.0, 28.4] SR:12 DR:14 LR:-72.01 LO:72.01);ALT=[chr14:36674745[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	43472430	+	chr8	43470750	+	.	11	0	5458126_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5458126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:43470750(-)-8:43472430(+)__8_43463001_43488001D;SPAN=1680;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:0 DR:11 LR:-15.99 LO:23.29);ALT=]chr8:43472430]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	43514714	+	chr8	43510735	+	.	61	21	5458212_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTCTTTTGATTCAGCAGATTG;MAPQ=60;MATEID=5458212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_43512001_43537001_216C;SPAN=3979;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:42 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:21 DR:61 LR:-221.2 LO:221.2);ALT=]chr8:43514714]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	35507715	+	chr14	35509508	+	.	0	73	8436509_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AAGACTTACGAATAG;MAPQ=60;MATEID=8436509_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_35500501_35525501_71C;SPAN=1793;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:55 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:73 DR:0 LR:-214.6 LO:214.6);ALT=G[chr14:35509508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35605641	+	chr14	35615069	+	.	110	60	8437121_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TTGTTGCCCAGGCTAGAGTGCAATGGC;MAPQ=60;MATEID=8437121_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_35598501_35623501_133C;SPAN=9428;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:154 DP:40 GQ:41.5 PL:[455.5, 41.5, 0.0] SR:60 DR:110 LR:-455.5 LO:455.5);ALT=C[chr14:35615069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	36418745	+	chr14	36417604	+	.	56	0	8440874_1	99.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=8440874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:36417604(-)-14:36418745(+)__14_36407001_36432001D;SPAN=1141;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:98 GQ:79.1 PL:[158.3, 0.0, 79.1] SR:0 DR:56 LR:-159.7 LO:159.7);ALT=]chr14:36418745]G;VARTYPE=BND:DUP-th;JOINTYPE=th
