chr18	14280465	+	chr18	14283681	+	.	68	27	9912486_1	99.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=TCAACACCAG;MAPQ=60;MATEID=9912486_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_14259001_14284001_26C;SPAN=3216;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:76 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:27 DR:68 LR:-260.8 LO:260.8);ALT=G[chr18:14283681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	14552177	+	chr18	14568726	+	.	44	28	9914726_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=TGGAACAT;MAPQ=0;MATEID=9914726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_14528501_14553501_431C;SPAN=16549;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:57 DP:33 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:28 DR:44 LR:-168.3 LO:168.3);ALT=T[chr18:14568726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
