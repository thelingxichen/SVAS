chr1	56831124	+	chr1	56834962	+	.	75	65	163717_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAAGAACCACTGCCTC;MAPQ=60;MATEID=163717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_56815501_56840501_43C;SPAN=3838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:50 GQ:30 PL:[330.0, 30.0, 0.0] SR:65 DR:75 LR:-330.1 LO:330.1);ALT=C[chr1:56834962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
