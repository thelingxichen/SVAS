chr4	49151360	+	chr4	49150189	+	.	22	0	2714026_1	0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2714026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:49150189(-)-4:49151360(+)__4_49147001_49172001D;SPAN=1171;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:22 DP:321 GQ:14 PL:[0.0, 14.0, 805.3] SR:0 DR:22 LR:14.34 LO:38.89);ALT=]chr4:49151360]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	49158225	+	chr4	49156678	+	.	8	0	2714079_1	0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=2714079_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:49156678(-)-4:49158225(+)__4_49147001_49172001D;SPAN=1547;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:317 GQ:59.3 PL:[0.0, 59.3, 887.9] SR:0 DR:8 LR:59.48 LO:10.62);ALT=]chr4:49158225]C;VARTYPE=BND:DUP-th;JOINTYPE=th
