chr1	892652	+	chr1	894592	+	.	9	0	2348_1	8.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:892652(+)-1:894592(-)__1_882001_907001D;SPAN=1940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:77 GQ:8.9 PL:[8.9, 0.0, 177.2] SR:0 DR:9 LR:-8.848 LO:18.1);ALT=G[chr1:894592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1159348	+	chr1	1163847	+	.	3	5	3263_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3263_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1151501_1176501_117C;SPAN=4499;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:81 GQ:1.8 PL:[0.0, 1.8, 198.0] SR:5 DR:3 LR:2.139 LO:10.82);ALT=C[chr1:1163847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1164327	+	chr1	1167272	+	.	130	11	3276_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1151501_1176501_123C;SPAN=2945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:66 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:11 DR:130 LR:-389.5 LO:389.5);ALT=C[chr1:1167272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1203374	+	chr1	1209046	+	.	0	10	3558_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1200501_1225501_230C;SPAN=5672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:10 DR:0 LR:-14.59 LO:21.18);ALT=T[chr1:1209046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1254907	+	chr1	1256376	+	ATGATCACACAGTCCAGGAAGTCTGTTAGGCGGCCGTTCTGGGTGATGTAGGAGAAGTCAGGGAAGCGTCG	0	38	4154_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTA;INSERTION=ATGATCACACAGTCCAGGAAGTCTGTTAGGCGGCCGTTCTGGGTGATGTAGGAGAAGTCAGGGAAGCGTCG;MAPQ=60;MATEID=4154_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_1_1249501_1274501_303C;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:90 GQ:99 PL:[101.0, 0.0, 117.5] SR:38 DR:0 LR:-101.1 LO:101.1);ALT=A[chr1:1256376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1254942	+	chr1	1259957	+	.	11	0	4155_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:1254942(+)-1:1259957(-)__1_1249501_1274501D;SPAN=5015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:0 DR:11 LR:-13.55 LO:22.7);ALT=T[chr1:1259957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1255958	+	chr1	1259957	+	.	18	0	4158_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:1255958(+)-1:1259957(-)__1_1249501_1274501D;SPAN=3999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:0 DR:18 LR:-35.58 LO:40.99);ALT=A[chr1:1259957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1256495	+	chr1	1259957	+	.	19	0	4159_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4159_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:1256495(+)-1:1259957(-)__1_1249501_1274501D;SPAN=3462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:84 GQ:40.1 PL:[40.1, 0.0, 162.2] SR:0 DR:19 LR:-39.96 LO:44.22);ALT=A[chr1:1259957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1337638	+	chr1	1341189	+	.	2	22	3734_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1323001_1348001_63C;SPAN=3551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:84 GQ:56.6 PL:[56.6, 0.0, 145.7] SR:22 DR:2 LR:-56.47 LO:58.71);ALT=T[chr1:1341189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1341266	+	chr1	1342289	+	.	0	48	3749_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1323001_1348001_291C;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:100 GQ:99 PL:[131.3, 0.0, 111.5] SR:48 DR:0 LR:-131.4 LO:131.4);ALT=G[chr1:1342289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1480382	+	chr1	1500153	+	.	7	12	4394_1	45.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=4394_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1494501_1519501_152C;SPAN=19771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:12 DR:7 LR:-45.01 LO:45.06);ALT=G[chr1:1500153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1480426	+	chr1	1509857	+	.	8	0	4395_1	18.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4395_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:1480426(+)-1:1509857(-)__1_1494501_1519501D;SPAN=29431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:30 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.28 LO:19.28);ALT=T[chr1:1509857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1500300	+	chr1	1509858	+	.	39	27	4411_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTGA;MAPQ=60;MATEID=4411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1494501_1519501_218C;SPAN=9558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:92 GQ:80.9 PL:[140.3, 0.0, 80.9] SR:27 DR:39 LR:-140.9 LO:140.9);ALT=A[chr1:1509858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	1718879	+	chr1	1720490	+	.	4	3	5344_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=5344_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_1715001_1740001_233C;SPAN=1611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:74 GQ:0 PL:[0.0, 0.0, 178.2] SR:3 DR:4 LR:0.2424 LO:11.06);ALT=G[chr1:1720490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2323397	+	chr1	2327221	+	.	30	9	7225_1	90.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7225_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_2303001_2328001_259C;SPAN=3824;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:67 GQ:71 PL:[90.8, 0.0, 71.0] SR:9 DR:30 LR:-90.9 LO:90.9);ALT=G[chr1:2327221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2323413	+	chr1	2328551	+	.	20	0	7293_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:2323413(+)-1:2328551(-)__1_2327501_2352501D;SPAN=5138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:39 GQ:38.9 PL:[55.4, 0.0, 38.9] SR:0 DR:20 LR:-55.6 LO:55.6);ALT=G[chr1:2328551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2327310	+	chr1	2328553	+	.	0	36	7294_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_2327501_2352501_18C;SPAN=1243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:36 DR:0 LR:-118.8 LO:118.8);ALT=G[chr1:2328553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2328660	+	chr1	2330851	+	.	0	11	7297_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=7297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_2327501_2352501_300C;SPAN=2191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:11 DR:0 LR:-16.53 LO:23.43);ALT=G[chr1:2330851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2332375	+	chr1	2334472	+	CATGCGGCTACCAAGGGCATCCTTGTGGCTATGGTCTGTACTTTCTTCGACGCTTTCAACGTCCCGGTGTTCTGGCCGATTCTGGTGATGTACTTCATCATGCTCTTCTGTATCACGATGAAGAGGCAAATCA	0	28	7306_1	69.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CATGCGGCTACCAAGGGCATCCTTGTGGCTATGGTCTGTACTTTCTTCGACGCTTTCAACGTCCCGGTGTTCTGGCCGATTCTGGTGATGTACTTCATCATGCTCTTCTGTATCACGATGAAGAGGCAAATCA;MAPQ=60;MATEID=7306_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_2327501_2352501_174C;SPAN=2097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:84 GQ:69.8 PL:[69.8, 0.0, 132.5] SR:28 DR:0 LR:-69.67 LO:70.79);ALT=G[chr1:2334472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2332375	+	chr1	2333645	+	.	2	5	7305_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=7305_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_2327501_2352501_174C;SPAN=1270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:75 GQ:0.3 PL:[0.0, 0.3, 181.5] SR:5 DR:2 LR:0.5133 LO:11.02);ALT=G[chr1:2333645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	2341891	+	chr1	2343827	+	.	0	10	7335_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=7335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_2327501_2352501_33C;SPAN=1936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=C[chr1:2343827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	3326686	+	chr1	3324958	+	.	15	0	9931_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:3324958(-)-1:3326686(+)__1_3307501_3332501D;SPAN=1728;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:98 GQ:23 PL:[23.0, 0.0, 214.4] SR:0 DR:15 LR:-22.96 LO:32.06);ALT=]chr1:3326686]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	3564125	+	chr1	3566494	+	.	7	2	10399_1	5.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=10399_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_3552501_3577501_194C;SPAN=2369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:66 GQ:5.3 PL:[5.3, 0.0, 153.8] SR:2 DR:7 LR:-5.226 LO:13.76);ALT=C[chr1:3566494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	3807656	+	chr1	3816735	+	.	8	0	11853_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=11853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:3807656(+)-1:3816735(-)__1_3797501_3822501D;SPAN=9079;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:0 DR:8 LR:-8.798 LO:16.28);ALT=T[chr1:3816735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	3809595	+	chr1	3816586	+	.	12	0	11857_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=11857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:3809595(+)-1:3816586(-)__1_3797501_3822501D;SPAN=6991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:0 DR:12 LR:-17.67 LO:25.46);ALT=C[chr1:3816586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
