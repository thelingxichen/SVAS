chr8	115516632	+	chr8	115598206	-	.	11	0	4032997_1	19.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4032997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:115516632(+)-8:115598206(+)__8_115591001_115616001D;SPAN=81574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:0 DR:11 LR:-19.51 LO:24.29);ALT=T]chr8:115598206];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	115887041	-	chr8	115888057	+	.	11	0	4033314_1	12.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4033314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:115887041(-)-8:115888057(-)__8_115885001_115910001D;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:89 GQ:12.2 PL:[12.2, 0.0, 203.6] SR:0 DR:11 LR:-12.2 LO:22.41);ALT=[chr8:115888057[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
