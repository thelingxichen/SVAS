chr18	52551749	+	chr18	52425822	+	TGAAATCATGAA	72	62	10025045_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=TGAAATCATGAA;MAPQ=60;MATEID=10025045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_52528001_52553001_208C;SPAN=125927;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:52 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:62 DR:72 LR:-300.4 LO:300.4);ALT=]chr18:52551749]A;VARTYPE=BND:DUP-th;JOINTYPE=th
