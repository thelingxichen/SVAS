chr8	80029360	+	chr8	80137002	+	.	17	0	5515795_1	50.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=5515795_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:80029360(+)-8:80137002(-)__8_80115001_80140001D;SPAN=107642;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:23 GQ:3.8 PL:[50.0, 0.0, 3.8] SR:0 DR:17 LR:-51.89 LO:51.89);ALT=C[chr8:80137002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
