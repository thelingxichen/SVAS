chr10	97208025	+	chr10	97206786	+	.	0	42	6456218_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TGCTC;MAPQ=60;MATEID=6456218_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_97191501_97216501_178C;SPAN=1239;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:42 DP:123 GQ:99 PL:[105.5, 0.0, 191.3] SR:42 DR:0 LR:-105.3 LO:106.7);ALT=]chr10:97208025]T;VARTYPE=BND:DUP-th;JOINTYPE=th
