chr1	76900621	+	chr1	76903367	+	.	42	22	359595_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=ATTCTCCTGCCTCAGCCTCTTGAGTAGCTGGGACTACAGGCA;MAPQ=60;MATEID=359595_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_1_76881001_76906001_13C;SPAN=2746;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:60 DP:76 GQ:5.9 PL:[177.5, 0.0, 5.9] SR:22 DR:42 LR:-187.0 LO:187.0);ALT=A[chr1:76903367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
