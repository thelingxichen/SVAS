chr2	10155443	+	chr2	10154282	+	.	9	0	910712_1	8.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=910712_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:10154282(-)-2:10155443(+)__2_10143001_10168001D;SPAN=1161;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-8.035 LO:17.94);ALT=]chr2:10155443]C;VARTYPE=BND:DUP-th;JOINTYPE=th
