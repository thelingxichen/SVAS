chr3	162525742	+	chr3	162547643	-	.	46	34	1759754_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=1759754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_162533001_162558001_293C;SPAN=21901;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:27 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:34 DR:46 LR:-217.9 LO:217.9);ALT=T]chr3:162547643];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	162545363	-	chr3	162547659	+	C	49	39	1759771_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=1759771_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_162533001_162558001_26C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:70 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:39 DR:49 LR:-221.2 LO:221.2);ALT=[chr3:162547659[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	162764901	+	chr3	162769085	+	GT	42	35	1760292_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GT;MAPQ=60;MATEID=1760292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_162753501_162778501_26C;SPAN=4184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:58 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:35 DR:42 LR:-184.8 LO:184.8);ALT=T[chr3:162769085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
