chr15	54199918	+	chr15	54203166	+	TT	0	42	5954419_1	99.0	.	EVDNC=ASSMB;INSERTION=TT;MAPQ=60;MATEID=5954419_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_54194001_54219001_99C;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:21 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:42 DR:0 LR:-122.1 LO:122.1);ALT=A[chr15:54203166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
