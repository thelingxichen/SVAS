chr2	18478317	+	chr18	70839198	+	.	0	7	6671584_1	19.0	.	EVDNC=ASSMB;HOMSEQ=ACTATATATAGTGTATATATACAC;MAPQ=54;MATEID=6671584_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_70829501_70854501_313C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:7 DP:6 GQ:1.8 PL:[19.8, 1.8, 0.0] SR:7 DR:0 LR:-19.8 LO:19.8);ALT=C[chr18:70839198[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	18906149	+	chr2	18907349	+	.	30	32	705881_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTT;MAPQ=60;MATEID=705881_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_18889501_18914501_206C;SPAN=1200;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:81 GQ:47.6 PL:[146.6, 0.0, 47.6] SR:32 DR:30 LR:-149.0 LO:149.0);ALT=T[chr2:18907349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	18907656	+	chr2	18906161	+	.	0	34	705882_1	87.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=705882_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_18889501_18914501_254C;SPAN=1495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:93 GQ:87.2 PL:[87.2, 0.0, 136.7] SR:34 DR:0 LR:-87.04 LO:87.69);ALT=]chr2:18907656]T;VARTYPE=BND:DUP-th;JOINTYPE=th
