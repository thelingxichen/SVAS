chr5	6374539	+	chr5	6377279	+	.	0	9	2408013_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2408013_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_6370001_6395001_1C;SPAN=2740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:9 DR:0 LR:-12.1 LO:18.81);ALT=T[chr5:6377279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	6377362	+	chr5	6378474	+	.	0	15	2408015_1	33.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2408015_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_6370001_6395001_219C;SPAN=1112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:61 GQ:33.2 PL:[33.2, 0.0, 112.4] SR:15 DR:0 LR:-32.99 LO:35.54);ALT=C[chr5:6378474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
