chr3	81957140	-	chr3	81958385	+	.	4	2	1509514_1	0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTG;MAPQ=60;MATEID=1509514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_81952501_81977501_149C;SPAN=1245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:131 GQ:21.9 PL:[0.0, 21.9, 359.7] SR:2 DR:4 LR:22.29 LO:5.643);ALT=[chr3:81958385[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
