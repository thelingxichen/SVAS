chr12	80191178	+	chr12	80199946	+	TGTTGATCTTCTAGATTGTCTTGCTTGTCTAGATCTTGCTTTTCTTTGGGATTCAGACTCTTCATCCCTAACAGGAGTGAGGTATGAT	0	12	5260915_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGTTGATCTTCTAGATTGTCTTGCTTGTCTAGATCTTGCTTTTCTTTGGGATTCAGACTCTTCATCCCTAACAGGAGTGAGGTATGAT;MAPQ=60;MATEID=5260915_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_80188501_80213501_142C;SPAN=8768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:83 GQ:17.3 PL:[17.3, 0.0, 182.3] SR:12 DR:0 LR:-17.13 LO:25.33);ALT=G[chr12:80199946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	80266720	+	chr12	80328474	+	.	0	7	5261102_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5261102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_80262001_80287001_26C;SPAN=61754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:43 GQ:11.6 PL:[11.6, 0.0, 90.8] SR:7 DR:0 LR:-11.46 LO:15.17);ALT=T[chr12:80328474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
