chr5	17144637	+	chr5	17145828	-	.	9	0	3246409_1	0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=3246409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:17144637(+)-5:17145828(+)__5_17125501_17150501D;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:181 GQ:19 PL:[0.0, 19.0, 475.3] SR:0 DR:9 LR:19.33 LO:14.62);ALT=T]chr5:17145828];VARTYPE=BND:INV-hh;JOINTYPE=hh
