chr4	155078005	+	chr4	155133914	+	.	9	0	3007808_1	13.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=3007808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:155078005(+)-4:155133914(-)__4_155060501_155085501D;SPAN=55909;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:61 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.18 LO:19.08);ALT=G[chr4:155133914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
