chr2	50925555	-	chr15	60831403	+	.	61	59	8916568_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=8916568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_60809001_60834001_17C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:51 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:59 DR:61 LR:-277.3 LO:277.3);ALT=[chr15:60831403[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
