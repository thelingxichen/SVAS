chr5	60001709	+	chr5	60003666	+	.	55	29	2482242_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACTAA;MAPQ=60;MATEID=2482242_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_60000501_60025501_102C;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:14 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:29 DR:55 LR:-208.0 LO:208.0);ALT=A[chr5:60003666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	60224834	+	chr5	60240822	+	.	10	0	2482501_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2482501_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:60224834(+)-5:60240822(-)__5_60221001_60246001D;SPAN=15988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:0 DR:10 LR:-20.28 LO:22.97);ALT=T[chr5:60240822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
