chr11	80766886	+	chr11	81440358	+	.	50	29	6975159_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TATTT;MAPQ=60;MATEID=6975159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_81438001_81463001_58C;SPAN=673472;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:6 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:29 DR:50 LR:-208.0 LO:208.0);ALT=T[chr11:81440358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
