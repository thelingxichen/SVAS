chr4	6651593	+	chr4	6652911	+	.	59	62	2620639_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CAGA;MAPQ=60;MATEID=2620639_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_6639501_6664501_103C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:21 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:62 DR:59 LR:-313.6 LO:313.6);ALT=A[chr4:6652911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
