chr14	85297116	+	chr14	85302156	+	.	53	29	8650270_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTTTCTAA;MAPQ=60;MATEID=8650270_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_85284501_85309501_315C;SPAN=5040;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:67 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:29 DR:53 LR:-208.0 LO:208.0);ALT=A[chr14:85302156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
