chr4	177241370	+	chr4	177245332	+	AAAAAATGTAGAAGATTTCACTGGACCTAGAGAAAGAAGTGATCTGGGATTTATCACATTTGATATAACTGCTG	3	23	2351718_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AT;INSERTION=AAAAAATGTAGAAGATTTCACTGGACCTAGAGAAAGAAGTGATCTGGGATTTATCACATTTGATATAACTGCTG;MAPQ=60;MATEID=2351718_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_177233001_177258001_240C;SPAN=3962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:97 GQ:56.3 PL:[56.3, 0.0, 178.4] SR:23 DR:3 LR:-56.25 LO:59.83);ALT=T[chr4:177245332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	177241370	+	chr4	177243321	+	.	11	17	2351717_1	23.0	.	DISC_MAPQ=58;EVDNC=TSI_L;MAPQ=60;MATEID=2351717_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAAA;SCTG=c_4_177233001_177258001_240C;SPAN=1951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:124 GQ:23.6 PL:[23.6, 0.0, 242.5] SR:17 DR:11 LR:-23.41 LO:34.92);ALT=T[chr4:177243321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	177245409	+	chr4	177249349	+	CTCTGAACCAAGTTGTCCTATGGGACAAGATTGTTTTGAGAGGTGATAATCCGAAGCTGCTGCTGAAAGATATGAAAACAAAATATTTTTTCTTTGACGATGGAAATGGTCTCAA	0	22	2351732_1	44.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTCTGAACCAAGTTGTCCTATGGGACAAGATTGTTTTGAGAGGTGATAATCCGAAGCTGCTGCTGAAAGATATGAAAACAAAATATTTTTTCTTTGACGATGGAAATGGTCTCAA;MAPQ=60;MATEID=2351732_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_177233001_177258001_229C;SPAN=3940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:103 GQ:44.9 PL:[44.9, 0.0, 203.3] SR:22 DR:0 LR:-44.72 LO:50.57);ALT=G[chr4:177249349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
