chr22	25663781	+	chr22	25921028	+	.	9	0	10858250_1	20.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=10858250_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:25663781(+)-22:25921028(-)__22_25921001_25946001D;SPAN=257247;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=G[chr22:25921028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	25980983	+	chr22	25684716	+	.	11	0	10858315_1	24.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=10858315_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:25684716(-)-22:25980983(+)__22_25970001_25995001D;SPAN=296267;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:43 GQ:24.8 PL:[24.8, 0.0, 77.6] SR:0 DR:11 LR:-24.66 LO:26.28);ALT=]chr22:25980983]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	25981267	+	chr22	25684761	+	.	12	0	10858316_1	25.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=10858316_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:25684761(-)-22:25981267(+)__22_25970001_25995001D;SPAN=296506;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=]chr22:25981267]T;VARTYPE=BND:DUP-th;JOINTYPE=th
