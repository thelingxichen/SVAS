chr8	128190458	-	chr8	128300943	+	.	70	31	5687742_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CACT;MAPQ=60;MATEID=5687742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_128282001_128307001_264C;SPAN=110485;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:96 DP:130 GQ:34.1 PL:[281.6, 0.0, 34.1] SR:31 DR:70 LR:-293.0 LO:293.0);ALT=[chr8:128300943[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
