chr3	107037949	+	chr3	107040333	+	AAAAT	66	24	2224601_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AAAAT;MAPQ=60;MATEID=2224601_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107040501_107065501_242C;SPAN=2384;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:0 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:24 DR:66 LR:-224.5 LO:224.5);ALT=G[chr3:107040333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107976819	-	chr4	160636493	+	.	12	0	3027994_1	21.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=3027994_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:107976819(-)-4:160636493(-)__4_160622001_160647001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:0 DR:12 LR:-21.73 LO:26.64);ALT=[chr4:160636493[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	155277476	+	chr4	160103543	+	ATTCC	4	16	4458204_1	52.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=ATTCC;MAPQ=60;MATEID=4458204_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_155256501_155281501_269C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:26 GQ:9.5 PL:[52.4, 0.0, 9.5] SR:16 DR:4 LR:-53.93 LO:53.93);ALT=]chr6:155277476]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	161013814	+	chr4	161019650	+	.	65	68	3028646_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3028646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_160989501_161014501_276C;SPAN=5836;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:42 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:68 DR:65 LR:-307.0 LO:307.0);ALT=G[chr4:161019650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	161579970	+	chr4	161739627	+	TG	0	50	3030667_1	99.0	.	EVDNC=ASSMB;INSERTION=TG;MAPQ=60;MATEID=3030667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_161724501_161749501_316C;SPAN=159657;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:46 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:50 DR:0 LR:-148.5 LO:148.5);ALT=C[chr4:161739627[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	161973471	-	chr4	179040992	+	.	7	2	3031471_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TATATATATATATATAT;MAPQ=60;MATEID=3031471_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TATATATATATATATA;SCTG=c_4_161969501_161994501_263C;SPAN=17067521;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:26 GQ:5.9 PL:[5.9, 0.0, 12.8] SR:2 DR:7 LR:-5.537 LO:5.903);ALT=[chr4:179040992[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	162449277	+	chr4	162451667	+	.	32	37	3033194_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=40;MATEID=3033194_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_162435001_162460001_276C;SPAN=2390;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:58 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:37 DR:32 LR:-174.9 LO:174.9);ALT=T[chr4:162451667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	163278361	+	chr4	163281513	+	CTTTTTTTTTTTTTTTCAAAAAAAA	71	49	3035978_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTTTTTTTTTTTTTTTCAAAAAAAA;MAPQ=60;MATEID=3035978_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_163268001_163293001_123C;SPAN=3152;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:87 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:49 DR:71 LR:-287.2 LO:287.2);ALT=G[chr4:163281513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	163394005	+	chr4	163396421	+	.	70	61	3036484_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=3036484_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_163390501_163415501_363C;SPAN=2416;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:88 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:61 DR:70 LR:-300.4 LO:300.4);ALT=A[chr4:163396421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	163579619	+	chr4	163578515	+	A	22	63	3037075_1	99.0	.	DISC_MAPQ=1;EVDNC=TSI_L;INSERTION=A;MAPQ=29;MATEID=3037075_2;MATENM=1;NM=1;NUMPARTS=3;SCTG=c_4_163562001_163587001_249C;SPAN=1104;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:68 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:63 DR:22 LR:-201.3 LO:201.3);ALT=]chr4:163579619]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	179614293	-	chr4	179758025	+	.	48	26	3097105_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3097105_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_179756501_179781501_171C;SPAN=143732;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:35 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:26 DR:48 LR:-208.0 LO:208.0);ALT=[chr4:179758025[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	179756231	-	chr4	179757248	+	.	10	0	3097106_1	24.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3097106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:179756231(-)-4:179757248(-)__4_179756501_179781501D;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:33 GQ:24.2 PL:[24.2, 0.0, 53.9] SR:0 DR:10 LR:-24.07 LO:24.77);ALT=[chr4:179757248[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	180088964	-	chr4	183738455	+	.	12	0	3108620_1	29.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=3108620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:180088964(-)-4:183738455(-)__4_183725501_183750501D;SPAN=3649491;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=[chr4:183738455[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	181108559	+	chr4	182770465	+	.	89	71	3104375_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=3104375_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_182770001_182795001_171C;SPAN=1661906;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:39 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:71 DR:89 LR:-340.0 LO:340.0);ALT=A[chr4:182770465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	181876802	+	chr4	181878289	+	.	62	32	3103035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTCTACAGCACTTTCT;MAPQ=60;MATEID=3103035_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_181863501_181888501_241C;SPAN=1487;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:26 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:32 DR:62 LR:-234.4 LO:234.4);ALT=T[chr4:181878289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	184655833	+	chr4	184658970	+	.	52	24	3112338_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGCCAGACCTATTATT;MAPQ=60;MATEID=3112338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_184632001_184657001_314C;SPAN=3137;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:26 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:24 DR:52 LR:-184.8 LO:184.8);ALT=T[chr4:184658970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	184674269	+	chr4	184675715	+	.	47	0	3112835_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3112835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:184674269(+)-4:184675715(-)__4_184656501_184681501D;SPAN=1446;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:103 GQ:99 PL:[127.4, 0.0, 120.8] SR:0 DR:47 LR:-127.2 LO:127.2);ALT=C[chr4:184675715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	155291071	+	chr7	90331761	+	.	26	0	5036930_1	70.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5036930_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:155291071(+)-7:90331761(-)__7_90331501_90356501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:57 GQ:67.1 PL:[70.4, 0.0, 67.1] SR:0 DR:26 LR:-70.39 LO:70.39);ALT=T[chr7:90331761[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	91862935	+	chr7	91272565	+	.	67	49	5043420_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=5043420_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_91850501_91875501_384C;SPAN=590370;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:86 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:49 DR:67 LR:-274.0 LO:274.0);ALT=]chr7:91862935]T;VARTYPE=BND:DUP-th;JOINTYPE=th
