chr2	83066855	+	chr2	83068235	+	.	16	15	869541_1	62.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AAGAATATCTTTCTTGT;MAPQ=60;MATEID=869541_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_83055001_83080001_132C;SPAN=1380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:60 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:15 DR:16 LR:-62.97 LO:63.12);ALT=T[chr2:83068235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
