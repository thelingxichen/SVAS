chr10	21260555	-	chr10	21261665	+	.	6	2	6131350_1	0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=ACTCCATCTCAAAAAA;MAPQ=27;MATEID=6131350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_21241501_21266501_314C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:106 GQ:8.7 PL:[0.0, 8.7, 273.9] SR:2 DR:6 LR:8.912 LO:10.09);ALT=[chr10:21261665[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	21738872	-	chr10	21739987	+	.	8	0	6133652_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6133652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:21738872(-)-10:21739987(-)__10_21731501_21756501D;SPAN=1115;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:0 DR:8 LR:5.29 LO:14.13);ALT=[chr10:21739987[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	21907820	+	chr10	21788860	+	GG	63	30	6134144_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GG;MAPQ=60;MATEID=6134144_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_21903001_21928001_374C;SPAN=118960;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:30 DR:63 LR:-237.7 LO:237.7);ALT=]chr10:21907820]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	21881510	+	chr10	21882769	-	.	6	2	6134491_1	0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=GGGAGGCTGAGGCAGGAGAAT;MAPQ=0;MATEID=6134491_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_10_21878501_21903501_113C;SECONDARY;SPAN=1259;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:205 GQ:28.9 PL:[0.0, 28.9, 554.5] SR:2 DR:6 LR:29.13 LO:12.14);ALT=C]chr10:21882769];VARTYPE=BND:INV-hh;JOINTYPE=hh
