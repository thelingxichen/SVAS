chr2	113647832	+	chr5	156992421	+	TCTTTCA	10	0	3870213_1	0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=TCTTTCA;MAPQ=60;MATEID=3870213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_156971501_156996501_392C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:220 GQ:26.5 PL:[0.0, 26.5, 587.5] SR:0 DR:10 LR:26.59 LO:15.85);ALT=A[chr5:156992421[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	19793248	+	chrX	63279355	+	AAAAGAG	0	7	1877802_1	6.0	.	EVDNC=ASSMB;INSERTION=AAAAGAG;MAPQ=60;MATEID=1877802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_19771501_19796501_250C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:62 GQ:6.5 PL:[6.5, 0.0, 141.8] SR:7 DR:0 LR:-6.31 LO:13.96);ALT=C[chrX:63279355[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	20447719	-	chr5	156761837	+	.	7	32	3869219_1	91.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTCT;MAPQ=60;MATEID=3869219_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_156751001_156776001_385C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:65 GQ:65 PL:[91.4, 0.0, 65.0] SR:32 DR:7 LR:-91.53 LO:91.53);ALT=[chr5:156761837[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	20988435	+	chr3	20996178	+	.	78	59	1883273_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1883273_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_3_20996501_21021501_341C;SPAN=7743;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:0 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:59 DR:78 LR:-313.6 LO:313.6);ALT=C[chr3:20996178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	21810659	+	chr3	22220997	-	.	7	0	1887451_1	0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=GAAAAC;MAPQ=60;MATEID=1887451_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_22197001_22222001_41C;SPAN=410338;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:7 DP:107 GQ:5.7 PL:[0.0, 5.7, 270.6] SR:0 DR:7 LR:5.882 LO:12.23);ALT=C]chr3:22220997];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	22092361	+	chr3	22097796	+	.	118	60	1887094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAATTCAATGTG;MAPQ=60;MATEID=1887094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_22074501_22099501_107C;SPAN=5435;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:151 DP:90 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:60 DR:118 LR:-445.6 LO:445.6);ALT=G[chr3:22097796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	156381897	-	chr5	156384532	+	GGAAAG	8	7	3867101_1	35.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=GGAAAG;MAPQ=9;MATEID=3867101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_156383501_156408501_182C;SPAN=2635;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:51 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:7 DR:8 LR:-35.7 LO:36.92);ALT=[chr5:156384532[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	156848575	+	chr5	156850881	+	.	24	0	3869988_1	69.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=3869988_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:156848575(+)-5:156850881(-)__5_156849001_156874001D;SPAN=2306;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:37 GQ:19.7 PL:[69.2, 0.0, 19.7] SR:0 DR:24 LR:-70.66 LO:70.66);ALT=T[chr5:156850881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	157101526	-	chr5	157103258	+	.	8	0	3870760_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3870760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:157101526(-)-5:157103258(-)__5_157094001_157119001D;SPAN=1732;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:130 GQ:8.7 PL:[0.0, 8.7, 333.3] SR:0 DR:8 LR:8.812 LO:13.76);ALT=[chr5:157103258[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	72609401	+	chr5	157541721	+	AAACT	59	45	3873171_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=AAACT;MAPQ=60;MATEID=3873171_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_157535001_157560001_463C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:83 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:45 DR:59 LR:-257.5 LO:257.5);ALT=]chr8:72609401]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	157796279	+	chr8	72609406	+	.	25	0	3874533_1	65.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3874533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:157796279(+)-8:72609406(-)__5_157780001_157805001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:63 GQ:65.6 PL:[65.6, 0.0, 85.4] SR:0 DR:25 LR:-65.46 LO:65.63);ALT=A[chr8:72609406[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
