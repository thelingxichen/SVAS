chr13	111258312	+	chr6	129409329	+	.	9	0	8331698_1	3.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=8331698_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:129409329(-)-13:111258312(+)__13_111254501_111279501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:0 DR:9 LR:-3.429 LO:17.14);ALT=]chr13:111258312]A;VARTYPE=BND:TRX-th;JOINTYPE=th
