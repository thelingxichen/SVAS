chr11	125735503	+	chr11	125654235	+	.	27	0	7259203_1	64.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=7259203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:125654235(-)-11:125735503(+)__11_125734001_125759001D;SPAN=81268;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:93 GQ:64.1 PL:[64.1, 0.0, 159.8] SR:0 DR:27 LR:-63.93 LO:66.28);ALT=]chr11:125735503]T;VARTYPE=BND:DUP-th;JOINTYPE=th
