chr2	103017412	+	chr2	102871060	+	.	85	59	1214163_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAGA;MAPQ=60;MATEID=1214163_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_102998001_103023001_83C;SPAN=146352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:122 DP:84 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:59 DR:85 LR:-359.8 LO:359.8);ALT=]chr2:103017412]G;VARTYPE=BND:DUP-th;JOINTYPE=th
