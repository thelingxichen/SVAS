chr3	171757562	+	chr3	171830240	+	.	12	4	1788978_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1788978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_171818501_171843501_114C;SPAN=72678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:4 DR:12 LR:-28.06 LO:32.03);ALT=G[chr3:171830240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
