chr3	19989015	+	chr3	19992295	+	.	11	3	1297274_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=1297274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_19992001_20017001_56C;SPAN=3280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:24 GQ:20 PL:[36.5, 0.0, 20.0] SR:3 DR:11 LR:-36.61 LO:36.61);ALT=T[chr3:19992295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
