chr20	25733134	+	chr20	26084131	+	.	0	8	10461585_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CTTTTTCA;MAPQ=60;MATEID=10461585_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_25725001_25750001_42C;SPAN=350997;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:8 DR:0 LR:-7.443 LO:16.0);ALT=A[chr20:26084131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	26260598	+	chr20	26261779	+	.	93	44	10465125_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GATGTGTGCATTCA;MAPQ=58;MATEID=10465125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_26239501_26264501_227C;SPAN=1181;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:125 DP:29 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:44 DR:93 LR:-369.7 LO:369.7);ALT=A[chr20:26261779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	26297651	+	chr20	26302711	+	.	137	19	10464978_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GAGCAGTTTTGAAACACTCTTTTTGTTGGATCTGCAAGTCGACATTTGGAGCGCTTTGAGGCCT;MAPQ=60;MATEID=10464978_2;MATENM=2;NM=3;NUMPARTS=2;SCTG=c_20_26288501_26313501_229C;SPAN=5060;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:154 DP:18 GQ:41.5 PL:[455.5, 41.5, 0.0] SR:19 DR:137 LR:-455.5 LO:455.5);ALT=T[chr20:26302711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
