chr2	73380753	-	chr2	73382152	+	.	8	0	1087095_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=1087095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:73380753(-)-2:73382152(-)__2_73377501_73402501D;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:143 GQ:12 PL:[0.0, 12.0, 369.6] SR:0 DR:8 LR:12.33 LO:13.42);ALT=[chr2:73382152[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
