chr3	6646214	-	chr3	6654638	+	.	16	43	1820416_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TAATTG;MAPQ=60;MATEID=1820416_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_6639501_6664501_380C;SPAN=8424;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:116 GQ:99 PL:[123.8, 0.0, 156.8] SR:43 DR:16 LR:-123.7 LO:123.9);ALT=[chr3:6654638[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	6646325	+	chr3	6650084	-	.	17	0	1820418_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1820418_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:6646325(+)-3:6650084(+)__3_6639501_6664501D;SPAN=3759;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:117 GQ:24.5 PL:[24.5, 0.0, 258.8] SR:0 DR:17 LR:-24.42 LO:35.92);ALT=A]chr3:6650084];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	6650160	+	chr3	6654638	+	AAATTTACTAGGAAATTTTAAGGAGAAGCAGGACATGTTTATGGTTCTCAGAGTATGTTCTCACAGATTAT	27	79	1820432_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=TAATTG;INSERTION=AAATTTACTAGGAAATTTTAAGGAGAAGCAGGACATGTTTATGGTTCTCAGAGTATGTTCTCACAGATTAT;MAPQ=60;MATEID=1820432_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_6639501_6664501_380C;SPAN=4478;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:82 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:79 DR:27 LR:-283.9 LO:283.9);ALT=T[chr3:6654638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
