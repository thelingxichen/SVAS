chrX	147509696	+	chrX	147511236	+	TG	50	34	7550679_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TG;MAPQ=60;MATEID=7550679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_147490001_147515001_178C;SPAN=1540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:17 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:34 DR:50 LR:-208.0 LO:208.0);ALT=G[chrX:147511236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
