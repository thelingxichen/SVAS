chr7	93327192	+	chr7	93332281	+	.	9	0	5050099_1	11.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=5050099_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:93327192(+)-7:93332281(-)__7_93320501_93345501D;SPAN=5089;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=A[chr7:93332281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31327365	+	chr7	93415631	+	.	6	49	5050614_1	99.0	.	DISC_MAPQ=8;EVDNC=ASDIS;HOMSEQ=ACCCCGTCTCTACTAAAAATACAAAAAA;MAPQ=32;MATEID=5050614_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_7_93394001_93419001_0C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:82 GQ:50.6 PL:[146.3, 0.0, 50.6] SR:49 DR:6 LR:-148.5 LO:148.5);ALT=]chr16:31327365]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	93416941	+	chr7	93422992	+	.	47	31	5050627_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAATCATCATTCTT;MAPQ=60;MATEID=5050627_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_93418501_93443501_375C;SPAN=6051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:32 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:31 DR:47 LR:-184.8 LO:184.8);ALT=T[chr7:93422992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
