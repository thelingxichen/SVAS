chr15	34382658	+	chr15	34388096	+	.	2	2	5921980_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5921980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_34373501_34398501_74C;SPAN=5438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:49 GQ:0 PL:[0.0, 0.0, 118.8] SR:2 DR:2 LR:0.0713 LO:7.387);ALT=T[chr15:34388096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	34388215	+	chr15	34393804	+	.	0	8	5921993_1	11.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5921993_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_34373501_34398501_78C;SPAN=5589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:8 DR:0 LR:-11.78 LO:16.98);ALT=C[chr15:34393804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	34517342	+	chr15	34519891	+	.	11	0	5922439_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5922439_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:34517342(+)-15:34519891(-)__15_34496001_34521001D;SPAN=2549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:0 DR:11 LR:-16.26 LO:23.36);ALT=T[chr15:34519891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	34517851	+	chr15	34519892	+	.	0	16	5922443_1	25.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5922443_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GCTGCT;SCTG=c_15_34496001_34521001_282C;SPAN=2041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:62 GQ:25.1 PL:[25.1, 0.0, 84.9] SR:16 DR:0 LR:-24.84 LO:27.14);ALT=G[chr15:34519892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
