chr8	4122884	+	chr8	4124973	+	TACATAATAATAT	0	37	3719676_1	99.0	.	EVDNC=ASSMB;INSERTION=TACATAATAATAT;MAPQ=60;MATEID=3719676_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_8_4116001_4141001_141C;SPAN=2089;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:22 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:37 DR:0 LR:-108.9 LO:108.9);ALT=T[chr8:4124973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
