chr1	19401391	+	chr1	19403232	+	.	4	3	60175_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=60175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19379501_19404501_28C;SPAN=1841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:85 GQ:0.2 PL:[0.2, 0.0, 204.8] SR:3 DR:4 LR:-0.07842 LO:12.95);ALT=C[chr1:19403232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19404564	+	chr1	19407842	+	.	0	11	59854_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CCTGG;MAPQ=60;MATEID=59854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19404001_19429001_216C;SPAN=3278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:89 GQ:12.2 PL:[12.2, 0.0, 203.6] SR:11 DR:0 LR:-12.2 LO:22.41);ALT=G[chr1:19407842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19537054	+	chr1	19566749	+	.	5	3	60338_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=60338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19551001_19576001_22C;SPAN=29695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:51 GQ:6.2 PL:[6.2, 0.0, 115.1] SR:3 DR:5 LR:-5.989 LO:12.08);ALT=G[chr1:19566749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19635138	+	chr1	19638321	+	.	0	47	60546_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=60546_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19624501_19649501_210C;SPAN=3183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:87 GQ:78.8 PL:[131.6, 0.0, 78.8] SR:47 DR:0 LR:-132.3 LO:132.3);ALT=T[chr1:19638321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19639383	+	chr1	19644093	+	.	0	7	60556_1	4.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=60556_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_19624501_19649501_218C;SPAN=4710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:68 GQ:4.7 PL:[4.7, 0.0, 159.8] SR:7 DR:0 LR:-4.684 LO:13.67);ALT=G[chr1:19644093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19666113	+	chr1	19670850	+	.	0	17	60633_1	34.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=60633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19649001_19674001_58C;SPAN=4737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:82 GQ:34.1 PL:[34.1, 0.0, 162.8] SR:17 DR:0 LR:-33.9 LO:38.83);ALT=T[chr1:19670850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19670930	+	chr1	19683915	+	CTACCAGGCGCCCGATGTTGGCTATGTGTGGGGAGCAGTCACTCACAGTTTCATCCTTCTCCATCTGTCTGGTAAGGCTGCCTCCGAGGTTCATGGTGCCAGAGCCAGATTTGTTGGTCTGCAGCCACAGCATCACCGTGGAGGTCAACTTGTAATGGGCGGTGCGACCGCTGGATTTCT	2	19	60789_1	50.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=CTACCAGGCGCCCGATGTTGGCTATGTGTGGGGAGCAGTCACTCACAGTTTCATCCTTCTCCATCTGTCTGGTAAGGCTGCCTCCGAGGTTCATGGTGCCAGAGCCAGATTTGTTGGTCTGCAGCCACAGCATCACCGTGGAGGTCAACTTGTAATGGGCGGTGCGACCGCTGGATTTCT;MAPQ=60;MATEID=60789_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_19673501_19698501_169C;SPAN=12985;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:45 GQ:50.6 PL:[50.6, 0.0, 57.2] SR:19 DR:2 LR:-50.53 LO:50.56);ALT=T[chr1:19683915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19671749	+	chr1	19683129	+	.	2	10	60649_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=60649_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_19649001_19674001_366C;SPAN=11380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:10 DR:2 LR:-26.02 LO:26.98);ALT=G[chr1:19683129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19683282	+	chr1	19705031	+	.	10	0	60869_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=60869_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19683282(+)-1:19705031(-)__1_19698001_19723001D;SPAN=21749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:32 GQ:24.5 PL:[24.5, 0.0, 50.9] SR:0 DR:10 LR:-24.34 LO:24.94);ALT=A[chr1:19705031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19684057	+	chr1	19705032	+	.	5	19	60823_1	72.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=60823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19673501_19698501_68C;SPAN=20975;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:27 GQ:3.9 PL:[72.6, 3.9, 0.0] SR:19 DR:5 LR:-73.72 LO:73.72);ALT=C[chr1:19705032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19705149	+	chr1	19711997	+	.	2	76	60889_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=60889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19698001_19723001_370C;SPAN=6848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:103 GQ:18.5 PL:[229.7, 0.0, 18.5] SR:76 DR:2 LR:-239.9 LO:239.9);ALT=T[chr1:19711997[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19705195	+	chr1	19811929	+	.	52	0	60891_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=60891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19705195(+)-1:19811929(-)__1_19698001_19723001D;SPAN=106734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:38 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=A[chr1:19811929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19712121	+	chr1	19746153	+	.	0	84	60916_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=60916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19698001_19723001_267C;SPAN=34032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:72 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:84 DR:0 LR:-247.6 LO:247.6);ALT=C[chr1:19746153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19712167	+	chr1	19811928	+	.	103	0	60917_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=60917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19712167(+)-1:19811928(-)__1_19698001_19723001D;SPAN=99761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:43 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:0 DR:103 LR:-303.7 LO:303.7);ALT=A[chr1:19811928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19746297	+	chr1	19811929	+	.	62	0	61010_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=61010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19746297(+)-1:19811929(-)__1_19796001_19821001D;SPAN=65632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:72 GQ:12.6 PL:[198.0, 12.6, 0.0] SR:0 DR:62 LR:-199.6 LO:199.6);ALT=A[chr1:19811929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19923606	+	chr1	19949968	+	TTTTAAAGAAGGTAAGTGAGAAAACAATTCCTAATCCAAAACCAG	33	123	61609_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TACCT;INSERTION=TTTTAAAGAAGGTAAGTGAGAAAACAATTCCTAATCCAAAACCAG;MAPQ=60;MATEID=61609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_19918501_19943501_210C;SECONDARY;SPAN=26362;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:51 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:123 DR:33 LR:-435.7 LO:435.7);ALT=A[chr1:19949968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19923625	+	chr1	19952878	+	.	13	0	61612_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=61612_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19923625(+)-1:19952878(-)__1_19918501_19943501D;SPAN=29253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:0 DR:13 LR:-30.18 LO:31.58);ALT=C[chr1:19952878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	19923696	+	chr17	62743560	-	.	74	0	61613_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=61613_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:19923696(+)-17:62743560(+)__1_19918501_19943501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:50 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:0 DR:74 LR:-217.9 LO:217.9);ALT=G]chr17:62743560];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr17	61628178	+	chr17	61655829	+	.	8	10	6462686_1	42.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6462686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_61617501_61642501_86C;SPAN=27651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:10 DR:8 LR:-42.57 LO:43.16);ALT=T[chr17:61655829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	61843556	+	chr17	61850772	+	.	16	5	6463414_1	28.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6463414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_61838001_61863001_31C;SPAN=7216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:91 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:5 DR:16 LR:-28.16 LO:35.26);ALT=T[chr17:61850772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	61904903	+	chr17	61907260	+	.	8	0	6463239_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6463239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:61904903(+)-17:61907260(-)__17_61887001_61912001D;SPAN=2357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=G[chr17:61907260[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	61904913	+	chr17	61906871	+	.	37	0	6463241_1	93.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6463241_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:61904913(+)-17:61906871(-)__17_61887001_61912001D;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:105 GQ:93.8 PL:[93.8, 0.0, 159.8] SR:0 DR:37 LR:-93.69 LO:94.67);ALT=C[chr17:61906871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	61905569	+	chr17	61906851	+	.	0	39	6463244_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6463244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_61887001_61912001_18C;SPAN=1282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:97 GQ:99 PL:[102.5, 0.0, 132.2] SR:39 DR:0 LR:-102.5 LO:102.7);ALT=G[chr17:61906851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62007747	+	chr17	62009555	+	TTGGGATTCCGGTACCGGTCCTCCGATCTGGCTGCTGGTACTGGCTCAG	8	8	6463842_1	43.0	.	DISC_MAPQ=53;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TTGGGATTCCGGTACCGGTCCTCCGATCTGGCTGCTGGTACTGGCTCAG;MAPQ=60;MATEID=6463842_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_62009501_62034501_173C;SPAN=1808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:36 GQ:43.1 PL:[43.1, 0.0, 43.1] SR:8 DR:8 LR:-43.06 LO:43.06);ALT=T[chr17:62009555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62082738	+	chr17	62083990	+	.	0	35	6464171_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCTGGA;MAPQ=60;MATEID=6464171_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_62083001_62108001_106C;SPAN=1252;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:47 GQ:10.4 PL:[102.8, 0.0, 10.4] SR:35 DR:0 LR:-107.1 LO:107.1);ALT=A[chr17:62083990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62082784	+	chr17	62097799	+	.	29	0	6464172_1	89.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6464172_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:62082784(+)-17:62097799(-)__17_62083001_62108001D;SPAN=15015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:31 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:29 LR:-89.12 LO:89.12);ALT=C[chr17:62097799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62084146	+	chr17	62097814	+	.	25	0	6464177_1	61.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6464177_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:62084146(+)-17:62097814(-)__17_62083001_62108001D;SPAN=13668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:77 GQ:61.7 PL:[61.7, 0.0, 124.4] SR:0 DR:25 LR:-61.66 LO:62.85);ALT=C[chr17:62097814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62474105	+	chr17	62476403	+	.	3	4	6465307_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=6465307_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_62475001_62500001_2C;SPAN=2298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:35 GQ:10.4 PL:[10.4, 0.0, 73.1] SR:4 DR:3 LR:-10.32 LO:13.15);ALT=C[chr17:62476403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62496893	+	chr17	62498128	+	.	9	16	6465367_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6465367_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_62475001_62500001_23C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:116 GQ:44.6 PL:[44.6, 0.0, 236.0] SR:16 DR:9 LR:-44.5 LO:52.03);ALT=T[chr17:62498128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62496893	+	chr17	62498555	+	AGCCCTCTGGAGGCCACATCTGTAGCAATCAGAATAGGAGCTTTTCCATGTTTGAATTCATTTAGAACCCAGTCACGCTCTTGTTGACTCTTGTCACCATGGATACCCATGGCAGGCC	11	21	6465368_1	51.0	.	DISC_MAPQ=54;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGCCCTCTGGAGGCCACATCTGTAGCAATCAGAATAGGAGCTTTTCCATGTTTGAATTCATTTAGAACCCAGTCACGCTCTTGTTGACTCTTGTCACCATGGATACCCATGGCAGGCC;MAPQ=60;MATEID=6465368_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_62475001_62500001_23C;SPAN=1662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:114 GQ:51.8 PL:[51.8, 0.0, 223.4] SR:21 DR:11 LR:-51.64 LO:57.8);ALT=T[chr17:62498555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	62500961	+	chr17	62502192	+	.	0	102	6465176_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=6465176_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_62499501_62524501_291C;SPAN=1231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:144 GQ:50.3 PL:[297.8, 0.0, 50.3] SR:102 DR:0 LR:-307.5 LO:307.5);ALT=C[chr17:62502192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
