chr2	159706408	+	chr2	159743368	+	.	11	0	1061060_1	27.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=1061060_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:159706408(+)-2:159743368(-)__2_159740001_159765001D;SPAN=36960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:34 GQ:27.2 PL:[27.2, 0.0, 53.6] SR:0 DR:11 LR:-27.1 LO:27.63);ALT=G[chr2:159743368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160139607	+	chr2	160143093	+	.	17	8	1062761_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=1062761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160132001_160157001_287C;SPAN=3486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:71 GQ:56.9 PL:[56.9, 0.0, 113.0] SR:8 DR:17 LR:-56.69 LO:57.8);ALT=G[chr2:160143093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160149126	+	chr2	160151649	+	.	50	36	1062789_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAGAATTTC;MAPQ=60;MATEID=1062789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160132001_160157001_316C;SPAN=2523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:134 GQ:99 PL:[188.3, 0.0, 135.5] SR:36 DR:50 LR:-188.6 LO:188.6);ALT=C[chr2:160151649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160569172	+	chr2	160585519	+	.	19	8	1063560_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1063560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160548501_160573501_351C;SPAN=16347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:49 GQ:52.7 PL:[52.7, 0.0, 65.9] SR:8 DR:19 LR:-52.75 LO:52.83);ALT=G[chr2:160585519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160628568	+	chr2	160636516	+	TAAATATTTCCTTTTGTATGGGA	11	12	1063736_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TAAATATTTCCTTTTGTATGGGA;MAPQ=60;MATEID=1063736_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160622001_160647001_174C;SPAN=7948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:90 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:12 DR:11 LR:-41.64 LO:46.37);ALT=A[chr2:160636516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160637510	+	chr2	160639869	+	.	0	68	1063771_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1063771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160622001_160647001_98C;SPAN=2359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:110 GQ:72.5 PL:[194.6, 0.0, 72.5] SR:68 DR:0 LR:-197.7 LO:197.7);ALT=C[chr2:160639869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160637559	+	chr2	160654641	+	.	55	0	1063998_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1063998_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:160637559(+)-2:160654641(-)__2_160646501_160671501D;SPAN=17082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:47 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:55 LR:-161.7 LO:161.7);ALT=A[chr2:160654641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160639981	+	chr2	160654643	+	.	46	13	1063999_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1063999_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_160646501_160671501_311C;SPAN=14662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:48 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:13 DR:46 LR:-145.2 LO:145.2);ALT=C[chr2:160654643[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160755605	+	chr2	160761145	+	.	13	0	1064091_1	21.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1064091_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:160755605(+)-2:160761145(-)__2_160744501_160769501D;SPAN=5540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:80 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:0 DR:13 LR:-21.24 LO:28.16);ALT=T[chr2:160761145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
