chr1	75190519	+	chr1	75198640	+	.	3	4	204919_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=204919_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_75190501_75215501_49C;SPAN=8121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:79 GQ:4.8 PL:[0.0, 4.8, 201.3] SR:4 DR:3 LR:4.898 LO:8.661);ALT=C[chr1:75198640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	75198972	+	chr1	75202224	+	.	8	0	204968_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=204968_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:75198972(+)-1:75202224(-)__1_75190501_75215501D;SPAN=3252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=T[chr1:75202224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	75204472	+	chr1	75214434	+	.	0	8	204976_1	5.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=204976_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_75190501_75215501_225C;SPAN=9962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:8 DR:0 LR:-5.818 LO:15.7);ALT=G[chr1:75214434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	76190524	+	chr1	76198327	+	.	13	0	206451_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=206451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:76190524(+)-1:76198327(-)__1_76195001_76220001D;SPAN=7803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:36 GQ:33.2 PL:[33.2, 0.0, 53.0] SR:0 DR:13 LR:-33.16 LO:33.44);ALT=C[chr1:76198327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	76194173	+	chr1	76198328	+	.	0	8	206453_1	16.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=206453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_76195001_76220001_65C;SPAN=4155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:37 GQ:16.4 PL:[16.4, 0.0, 72.5] SR:8 DR:0 LR:-16.38 LO:18.44);ALT=G[chr1:76198328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	76210423	+	chr14	75348734	-	.	19	0	5802178_1	52.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=5802178_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:76210423(+)-14:75348734(+)__14_75337501_75362501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:38 GQ:39.2 PL:[52.4, 0.0, 39.2] SR:0 DR:19 LR:-52.52 LO:52.52);ALT=G]chr14:75348734];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	76253290	+	chr1	76254844	+	.	18	7	206609_1	58.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=206609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_76244001_76269001_314C;SPAN=1554;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:64 GQ:58.7 PL:[58.7, 0.0, 95.0] SR:7 DR:18 LR:-58.58 LO:59.1);ALT=G[chr1:76254844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74946991	+	chr14	74951118	+	GATCTGTACTGGGATTTCCCAGCAGAAGAGACTTTGGTTTTTGTCATCCTGAAGTTGCCACTCCACCACCAGTTTTAT	8	60	5801006_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=GATCTGTACTGGGATTTCCCAGCAGAAGAGACTTTGGTTTTTGTCATCCTGAAGTTGCCACTCCACCACCAGTTTTAT;MAPQ=60;MATEID=5801006_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_74945501_74970501_186C;SPAN=4127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:104 GQ:64.4 PL:[186.5, 0.0, 64.4] SR:60 DR:8 LR:-189.5 LO:189.5);ALT=C[chr14:74951118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74951290	+	chr14	74953032	+	.	5	123	5801022_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;MAPQ=60;MATEID=5801022_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74945501_74970501_247C;SPAN=1742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:128 DP:164 GQ:18.4 PL:[378.2, 0.0, 18.4] SR:123 DR:5 LR:-397.4 LO:397.4);ALT=T[chr14:74953032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74951343	+	chr14	74959893	+	.	103	0	5801023_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5801023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:74951343(+)-14:74959893(-)__14_74945501_74970501D;SPAN=8550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:93 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:0 DR:103 LR:-303.7 LO:303.7);ALT=T[chr14:74959893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	74953140	+	chr14	74959894	+	.	105	34	5801031_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=5801031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_74945501_74970501_29C;SPAN=6754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:119 DP:138 GQ:20.7 PL:[376.2, 20.7, 0.0] SR:34 DR:105 LR:-383.4 LO:383.4);ALT=C[chr14:74959894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	75520411	+	chr14	75530654	+	.	33	0	5802778_1	81.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5802778_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:75520411(+)-14:75530654(-)__14_75509001_75534001D;SPAN=10243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:102 GQ:81.5 PL:[81.5, 0.0, 164.0] SR:0 DR:33 LR:-81.3 LO:82.9);ALT=A[chr14:75530654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	75618848	+	chr14	75643058	+	.	0	46	5803094_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5803094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_75631501_75656501_45C;SPAN=24210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:57 GQ:1.1 PL:[136.4, 0.0, 1.1] SR:46 DR:0 LR:-144.4 LO:144.4);ALT=T[chr14:75643058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	76121320	+	chr14	76123713	+	.	0	14	5804539_1	35.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5804539_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_76097001_76122001_360C;SPAN=2393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:40 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:14 DR:0 LR:-35.38 LO:35.77);ALT=C[chr14:76123713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	76123878	+	chr14	76127117	+	.	29	4	5804408_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5804408_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_76121501_76146501_311C;SPAN=3239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:91 GQ:71.3 PL:[71.3, 0.0, 147.2] SR:4 DR:29 LR:-71.08 LO:72.62);ALT=T[chr14:76127117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	76452209	+	chr14	76488667	+	.	10	0	5805339_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5805339_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:76452209(+)-14:76488667(-)__14_76464501_76489501D;SPAN=36458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:0 DR:10 LR:-20.82 LO:23.18);ALT=G[chr14:76488667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	76618371	+	chr14	76620695	+	.	9	0	5805608_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5805608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:76618371(+)-14:76620695(-)__14_76611501_76636501D;SPAN=2324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:0 DR:9 LR:-6.139 LO:17.59);ALT=T[chr14:76620695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
