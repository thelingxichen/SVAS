chr4	181876802	+	chr4	181878289	+	.	123	70	2365718_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTCTACAGCACTTTCT;MAPQ=60;MATEID=2365718_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_181863501_181888501_254C;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:64 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:70 DR:123 LR:-458.8 LO:458.8);ALT=T[chr4:181878289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
