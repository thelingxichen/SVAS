chr17	69791899	+	chr17	69793366	-	.	8	0	9794998_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=9794998_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:69791899(+)-17:69793366(+)__17_69776001_69801001D;SPAN=1467;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:139 GQ:11.1 PL:[0.0, 11.1, 359.7] SR:0 DR:8 LR:11.25 LO:13.52);ALT=G]chr17:69793366];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	126979420	+	chr17	69996998	+	.	7	58	9796009_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATAGATAGATAGATAGATAGAT;MAPQ=60;MATEID=9796009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_69996501_70021501_49C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:45 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:58 DR:7 LR:-171.6 LO:171.6);ALT=]chrX:126979420]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	70635365	+	chr17	70506244	+	.	56	58	9798538_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=9798538_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_70633501_70658501_428C;SPAN=129121;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:101 GQ:13.8 PL:[270.6, 13.8, 0.0] SR:58 DR:56 LR:-275.6 LO:275.6);ALT=]chr17:70635365]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	70680629	+	chr17	70520588	+	T	53	31	9799733_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=9799733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_70658001_70683001_143C;SPAN=160041;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:74 DP:103 GQ:31.7 PL:[216.5, 0.0, 31.7] SR:31 DR:53 LR:-224.0 LO:224.0);ALT=]chr17:70680629]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	126144028	+	chrX	126124709	+	GTGAAAA	48	36	11375786_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=GTGAAAA;MAPQ=60;MATEID=11375786_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_126101501_126126501_77C;SPAN=19319;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:40 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:36 DR:48 LR:-208.0 LO:208.0);ALT=]chrX:126144028]A;VARTYPE=BND:DUP-th;JOINTYPE=th
