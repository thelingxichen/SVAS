chr7	77705958	+	chr7	77707317	-	.	9	0	4989011_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4989011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:77705958(+)-7:77707317(+)__7_77689501_77714501D;SPAN=1359;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:123 GQ:3.3 PL:[0.0, 3.3, 303.6] SR:0 DR:9 LR:3.615 LO:16.17);ALT=T]chr7:77707317];VARTYPE=BND:INV-hh;JOINTYPE=hh
