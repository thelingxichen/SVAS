chr12	19373868	+	chr5	44529751	+	.	0	26	5255583_1	71.0	.	BX=CTCTGTGGTCGCGGTT-1_1,TGTCTCGGTCCTCCAT-1_1,GGCAATTAGGTAACGC-1_3,ACCTTCGGTACGGTGA-1_1,CCAACTCTCGGGCACT-1_1,TTTGAGGAGGGAACGG-1_1,CCAGGGTTCTATCCAT-1_1,GATTCAGTCAACAGTC-1_1,TCGTAGATCAAGATCC-1_1,TTTGTCATCCTTAATC-1_1,TGCAACATCGGCACCA-1_2,CTGCGAGCATATGCGT-1_1,GAGCCGTGTCGTTGGC-1_1,CAGCCGAAGGACACCA-1_1,GGACTTATCCTCGCAT-1_2,ATCACTTCATGACATC-1_1,GAGCAGATCGACGGAA-1_1,TGGAGCCCAATGGGAC-1_2,GGAAAGCCAGAACAGC-1_1,ATGTGTGAGAGAGAGT-1_1,CTGGTCTGTACTACAC-1_1;EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=5255583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_44516501_44541501_73C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:24 GQ:6.6 PL:[0.0, 6.6, 72.6] SR:0 DR:0 LR:6.743 LO:0.0),OC001T.bam(GT:0/1 AD:26 DP:52 GQ:58.1 PL:[71.3, 0.0, 58.1] SR:26 DR:0 LR:-71.27 LO:71.27);ALT=]chr12:19373868]a;VARTYPE=BND:TRX-ht;JOINTYPE=ht	.
chr5	44532859	+	chr12	19373619	+	.	0	29	10751927_1	79.0	.	BX=TGCAACATCGGCACCA-1_1,CATCAAGTCCAAACTG-1_1,CGTCCATTCTAATGGC-1_1,GAAGTCTAGGCAGTCA-1_2,CTACCTGCATGTAAGA-1_1,TCGTAGATCAAGATCC-1_1,GGACTTATCCTCGCAT-1_2,TCGACGGAGGGTGAAA-1_1,CGATAACGTCCAGTAT-1_1,TGTAGTGGTAGGGATC-1_1,CGACTCTCAAGCCATT-1_2,ACCACCTAGAACTCCT-1_1,GGAAAGCCAGAACAGC-1_1,CGCTATCCAAGAAAGG-1_1,TTTGAGGAGGGAACGG-1_1,CTGGTCTGTACTACAC-1_1,GATTCAGTCAACAGTC-1_1,TCGGAATTCTGCTGTC-1_1,AGCGGTCAGGCTAGCA-1_1,AGGAAGCCAGAACAGC-1_1,CCAACTCTCGGGCACT-1_1,CATCGTCGTCACCAGC-1_2,AAGCTACGTTTCCTGC-1_1,CTGCGAGCATATGCGT-1_1;EVDNC=ASSMB;HOMSEQ=TATT;MAPQ=60;MATEID=10751927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_19355001_19380001_17C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:35 GQ:9.6 PL:[0.0, 9.6, 105.6] SR:0 DR:0 LR:9.834 LO:0.0),OC001T.bam(GT:0/1 AD:29 DP:57 GQ:63.2 PL:[79.7, 0.0, 63.2] SR:29 DR:0 LR:-79.81 LO:79.81);ALT=T[chr12:19373619[;VARTYPE=BND:TRX-th;JOINTYPE=th	.
chr5	44532859	+	chr12	19373619	+	.	0	29	10751927_1	79.0	.	BX=TGCAACATCGGCACCA-1_1,CATCAAGTCCAAACTG-1_1,CGTCCATTCTAATGGC-1_1,GAAGTCTAGGCAGTCA-1_2,CTACCTGCATGTAAGA-1_1,TCGTAGATCAAGATCC-1_1,GGACTTATCCTCGCAT-1_2,TCGACGGAGGGTGAAA-1_1,CGATAACGTCCAGTAT-1_1,TGTAGTGGTAGGGATC-1_1,CGACTCTCAAGCCATT-1_2,ACCACCTAGAACTCCT-1_1,GGAAAGCCAGAACAGC-1_1,CGCTATCCAAGAAAGG-1_1,TTTGAGGAGGGAACGG-1_1,CTGGTCTGTACTACAC-1_1,GATTCAGTCAACAGTC-1_1,TCGGAATTCTGCTGTC-1_1,AGCGGTCAGGCTAGCA-1_1,AGGAAGCCAGAACAGC-1_1,CCAACTCTCGGGCACT-1_1,CATCGTCGTCACCAGC-1_2,AAGCTACGTTTCCTGC-1_1,CTGCGAGCATATGCGT-1_1;EVDNC=ASSMB;HOMSEQ=TATT;MAPQ=60;MATEID=10751927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_19355001_19380001_17C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:35 GQ:9.6 PL:[0.0, 9.6, 105.6] SR:0 DR:0 LR:9.834 LO:0.0),OC001T.bam(GT:0/1 AD:29 DP:57 GQ:63.2 PL:[79.7, 0.0, 63.2] SR:29 DR:0 LR:-79.81 LO:79.81);ALT=T[chr12:19373619[;VARTYPE=BND:TRX-th;JOINTYPE=th	.
chr12	19373868	+	chr5	44529751	+	.	0	26	5255583_1	71.0	.	BX=CTCTGTGGTCGCGGTT-1_1,TGTCTCGGTCCTCCAT-1_1,GGCAATTAGGTAACGC-1_3,ACCTTCGGTACGGTGA-1_1,CCAACTCTCGGGCACT-1_1,TTTGAGGAGGGAACGG-1_1,CCAGGGTTCTATCCAT-1_1,GATTCAGTCAACAGTC-1_1,TCGTAGATCAAGATCC-1_1,TTTGTCATCCTTAATC-1_1,TGCAACATCGGCACCA-1_2,CTGCGAGCATATGCGT-1_1,GAGCCGTGTCGTTGGC-1_1,CAGCCGAAGGACACCA-1_1,GGACTTATCCTCGCAT-1_2,ATCACTTCATGACATC-1_1,GAGCAGATCGACGGAA-1_1,TGGAGCCCAATGGGAC-1_2,GGAAAGCCAGAACAGC-1_1,ATGTGTGAGAGAGAGT-1_1,CTGGTCTGTACTACAC-1_1;EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=5255583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_44516501_44541501_73C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:24 GQ:6.6 PL:[0.0, 6.6, 72.6] SR:0 DR:0 LR:6.743 LO:0.0),OC001T.bam(GT:0/1 AD:26 DP:52 GQ:58.1 PL:[71.3, 0.0, 58.1] SR:26 DR:0 LR:-71.27 LO:71.27);ALT=]chr12:19373868]a;VARTYPE=BND:TRX-ht;JOINTYPE=ht	.
