chr12	12562192	+	chr12	101274977	+	.	0	16	7403548_1	33.0	.	EVDNC=ASSMB;HOMSEQ=GGGTACA;MAPQ=60;MATEID=7403548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_12544001_12569001_396C;SPAN=88712785;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:71 GQ:33.8 PL:[33.8, 0.0, 136.1] SR:16 DR:0 LR:-33.58 LO:37.21);ALT=A[chr12:101274977[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	13303668	-	chr12	13304737	+	.	9	0	7409280_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7409280_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:13303668(-)-12:13304737(-)__12_13279001_13304001D;SPAN=1069;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:0 DR:9 LR:-4.242 LO:17.27);ALT=[chr12:13304737[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
