chr6	11882569	+	chr6	12144133	+	.	30	0	4028876_1	79.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=4028876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:11882569(+)-6:12144133(-)__6_12127501_12152501D;SPAN=261564;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:74 GQ:79.1 PL:[79.1, 0.0, 98.9] SR:0 DR:30 LR:-78.98 LO:79.13);ALT=A[chr6:12144133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	12144599	+	chr6	11883055	+	.	37	0	4028877_1	99.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=4028877_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:11883055(-)-6:12144599(+)__6_12127501_12152501D;SPAN=261544;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:71 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.2 LO:103.2);ALT=]chr6:12144599]A;VARTYPE=BND:DUP-th;JOINTYPE=th
