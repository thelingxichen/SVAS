chr14	78864270	+	chr14	78867030	+	.	74	22	8626175_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGT;MAPQ=60;MATEID=8626175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_78865501_78890501_231C;SPAN=2760;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:46 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:22 DR:74 LR:-257.5 LO:257.5);ALT=T[chr14:78867030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
