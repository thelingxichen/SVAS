chr11	89047641	+	chr6	65967557	+	.	8	0	4953255_1	15.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=4953255_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:65967557(-)-11:89047641(+)__11_89033001_89058001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:0 DR:8 LR:-15.84 LO:18.23);ALT=]chr11:89047641]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	66260039	+	chr6	66262022	+	.	71	13	2884261_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AAAGATATAGTA;MAPQ=60;MATEID=2884261_2;MATENM=1;NM=1;NUMPARTS=3;REPSEQ=AA;SCTG=c_6_66248001_66273001_327C;SPAN=1983;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:69 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:13 DR:71 LR:-237.7 LO:237.7);ALT=T[chr6:66262022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	90770461	+	chr8	90777567	+	.	6	4	3964422_1	13.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3964422_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAA;SCTG=c_8_90772501_90797501_234C;SPAN=7106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:37 GQ:13.1 PL:[13.1, 0.0, 75.8] SR:4 DR:6 LR:-13.08 LO:15.67);ALT=G[chr8:90777567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	90995115	+	chr8	90996759	+	.	11	0	3965103_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3965103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:90995115(+)-8:90996759(-)__8_90993001_91018001D;SPAN=1644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:0 DR:11 LR:-13.28 LO:22.64);ALT=G[chr8:90996759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91013789	+	chr8	91029351	+	.	30	4	3965168_1	94.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3965168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_91017501_91042501_98C;SPAN=15562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:43 GQ:8.3 PL:[94.1, 0.0, 8.3] SR:4 DR:30 LR:-97.88 LO:97.88);ALT=G[chr8:91029351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91031400	+	chr8	91033137	+	.	0	7	3965198_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3965198_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_91017501_91042501_230C;SPAN=1737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:7 DR:0 LR:-0.6203 LO:13.03);ALT=T[chr8:91033137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91057225	+	chr8	91064064	+	CATTAAATTTGACGGTGGAGAGGAAGTACTTATTTCAGGGGAATTCAACGACCTGAGAA	2	47	3965318_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=CATTAAATTTGACGGTGGAGAGGAAGTACTTATTTCAGGGGAATTCAACGACCTGAGAA;MAPQ=60;MATEID=3965318_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_91042001_91067001_338C;SPAN=6839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:88 GQ:81.8 PL:[131.3, 0.0, 81.8] SR:47 DR:2 LR:-131.9 LO:131.9);ALT=T[chr8:91064064[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91404361	-	chr8	91406052	+	.	9	0	3966557_1	9.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=3966557_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:91404361(-)-8:91406052(-)__8_91385001_91410001D;SPAN=1691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=[chr8:91406052[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	91933624	-	chr8	91935001	+	.	3	2	3967562_1	0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=GTGAGCCACCA;MAPQ=32;MATEID=3967562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_91924001_91949001_356C;SPAN=1377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:108 GQ:15.9 PL:[0.0, 15.9, 293.7] SR:2 DR:3 LR:16.06 LO:5.98);ALT=[chr8:91935001[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	91990883	+	chr8	91992590	+	.	0	7	3967712_1	0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=3967712_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_91973001_91998001_154C;SPAN=1707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:85 GQ:0.2 PL:[0.2, 0.0, 204.8] SR:7 DR:0 LR:-0.07842 LO:12.95);ALT=G[chr8:91992590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91992690	+	chr8	91997342	+	.	7	4	3967716_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3967716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_91973001_91998001_26C;SPAN=4652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:4 DR:7 LR:-17.84 LO:22.11);ALT=C[chr8:91997342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	92033634	+	chr8	92052872	+	.	14	11	3967831_1	49.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3967831_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_92046501_92071501_263C;SPAN=19238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:48 GQ:49.7 PL:[49.7, 0.0, 66.2] SR:11 DR:14 LR:-49.72 LO:49.85);ALT=T[chr8:92052872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	92186284	+	chr11	90133210	+	.	4	23	3968373_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TTTTCT;MAPQ=60;MATEID=3968373_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTTTTTTTTTTTTT;SCTG=c_8_92169001_92194001_321C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:39 GQ:2.5 PL:[25.9, 0.0, 2.5] SR:23 DR:4 LR:-27.33 LO:27.33);ALT=T[chr11:90133210[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	88068251	+	chr11	88070668	+	.	0	57	4951029_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4951029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_88053001_88078001_298C;SPAN=2417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:104 GQ:90.8 PL:[160.1, 0.0, 90.8] SR:57 DR:0 LR:-161.0 LO:161.0);ALT=C[chr11:88070668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	88964485	+	chr11	88967931	+	.	0	85	4952907_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TGT;MAPQ=60;MATEID=4952907_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_88959501_88984501_244C;SPAN=3446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:43 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:85 DR:0 LR:-250.9 LO:250.9);ALT=T[chr11:88967931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	89507200	-	chr11	89810561	+	.	36	19	4954284_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTGGGTGACAGAGC;MAPQ=0;MATEID=4954284_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_89498501_89523501_113C;SPAN=303361;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:42 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:19 DR:36 LR:-148.5 LO:148.5);ALT=[chr11:89810561[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	90421832	-	chr11	91808875	+	.	12	0	4960025_1	33.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4960025_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:90421832(-)-11:91808875(-)__11_91801501_91826501D;SPAN=1387043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:24 GQ:23.3 PL:[33.2, 0.0, 23.3] SR:0 DR:12 LR:-33.17 LO:33.17);ALT=[chr11:91808875[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
