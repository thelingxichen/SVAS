chr7	114563183	+	chr7	114582329	+	.	5	3	3535793_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3535793_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_7_114562001_114587001_78C;SPAN=19146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:3 DR:5 LR:0.4634 LO:12.88);ALT=G[chr7:114582329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
