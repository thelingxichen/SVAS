chr9	20973939	+	chr9	20972549	+	.	11	0	5798749_1	17.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5798749_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:20972549(-)-9:20973939(+)__9_20972001_20997001D;SPAN=1390;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:72 GQ:17 PL:[17.0, 0.0, 155.6] SR:0 DR:11 LR:-16.8 LO:23.5);ALT=]chr9:20973939]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	21025578	+	chr9	24390962	-	.	59	60	5802155_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=5802155_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_24377501_24402501_89C;SPAN=3365384;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:13 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:60 DR:59 LR:-303.7 LO:303.7);ALT=A]chr9:24390962];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	22233015	-	chr9	25350745	+	.	66	57	5802398_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=5802398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_25333001_25358001_75C;SPAN=3117730;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:12 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:57 DR:66 LR:-316.9 LO:316.9);ALT=[chr9:25350745[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
