chr5	143515053	+	chr5	143512489	+	.	80	47	3814586_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3814586_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_143496501_143521501_310C;SPAN=2564;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:125 GQ:7.2 PL:[316.8, 7.2, 0.0] SR:47 DR:80 LR:-330.2 LO:330.2);ALT=]chr5:143515053]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	143512867	+	chr5	143515048	+	GAATAAGCTC	0	47	3814588_1	99.0	.	EVDNC=ASSMB;INSERTION=GAATAAGCTC;MAPQ=60;MATEID=3814588_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_143496501_143521501_23C;SPAN=2181;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:129 GQ:99 PL:[120.2, 0.0, 192.8] SR:47 DR:0 LR:-120.2 LO:121.1);ALT=G[chr5:143515048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
