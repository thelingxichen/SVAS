chr18	72163701	+	chr18	72168561	+	.	9	0	6674636_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6674636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:72163701(+)-18:72168561(-)__18_72152501_72177501D;SPAN=4860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=G[chr18:72168561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	72167268	+	chr18	72168562	+	.	8	6	6674640_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6674640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_72152501_72177501_308C;SPAN=1294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:6 DR:8 LR:-17.89 LO:23.8);ALT=G[chr18:72168562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
