chr5	145199583	+	chr5	145202640	+	.	0	10	2604677_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2604677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_145187001_145212001_64C;SPAN=3057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:10 DR:0 LR:-21.63 LO:23.53);ALT=T[chr5:145202640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145547830	+	chr5	145551472	+	.	0	19	2605265_1	45.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2605265_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_145530001_145555001_91C;SPAN=3642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:65 GQ:45.2 PL:[45.2, 0.0, 111.2] SR:19 DR:0 LR:-45.11 LO:46.71);ALT=T[chr5:145551472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145552387	+	chr5	145562106	+	.	9	0	2605390_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2605390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:145552387(+)-5:145562106(-)__5_145554501_145579501D;SPAN=9719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=T[chr5:145562106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145557275	+	chr5	145562106	+	.	32	0	2605398_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2605398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:145557275(+)-5:145562106(-)__5_145554501_145579501D;SPAN=4831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:61 GQ:56.3 PL:[89.3, 0.0, 56.3] SR:0 DR:32 LR:-89.43 LO:89.43);ALT=G[chr5:145562106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145583272	+	chr5	145598547	+	.	8	0	2605345_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2605345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:145583272(+)-5:145598547(-)__5_145579001_145604001D;SPAN=15275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:69 GQ:7.7 PL:[7.7, 0.0, 159.5] SR:0 DR:8 LR:-7.714 LO:16.06);ALT=T[chr5:145598547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145583387	+	chr5	145602964	+	ATGTGATGCTGATCCTTCAGCCTTAGCCAACTATGTTGTAGCACTGGTCAAGAAGGACAAACCTGAGAAAGAATTAAAAGCCTTTTGTGCTGATCAACTTGATGTCTTTTTACAAAA	2	46	2605347_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATGTGATGCTGATCCTTCAGCCTTAGCCAACTATGTTGTAGCACTGGTCAAGAAGGACAAACCTGAGAAAGAATTAAAAGCCTTTTGTGCTGATCAACTTGATGTCTTTTTACAAAA;MAPQ=60;MATEID=2605347_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_145579001_145604001_110C;SPAN=19577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:71 GQ:37.1 PL:[132.8, 0.0, 37.1] SR:46 DR:2 LR:-135.4 LO:135.4);ALT=T[chr5:145602964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145598666	+	chr5	145602964	+	.	2	16	2605373_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2605373_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_5_145579001_145604001_110C;SPAN=4298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:56 GQ:44.3 PL:[44.3, 0.0, 90.5] SR:16 DR:2 LR:-44.25 LO:45.16);ALT=G[chr5:145602964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145826983	+	chr5	145834615	+	.	29	0	2605788_1	80.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2605788_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:145826983(+)-5:145834615(-)__5_145824001_145849001D;SPAN=7632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:58 GQ:60.2 PL:[80.0, 0.0, 60.2] SR:0 DR:29 LR:-80.16 LO:80.16);ALT=T[chr5:145834615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	145843358	+	chr5	145849105	+	.	3	4	2605825_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2605825_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_145848501_145873501_215C;SPAN=5747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:29 GQ:11.9 PL:[11.9, 0.0, 58.1] SR:4 DR:3 LR:-11.95 LO:13.7);ALT=T[chr5:145849105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
