chr2	226854066	+	chr2	226860379	-	.	47	34	1725305_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=1725305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_226845501_226870501_227C;SPAN=6313;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:69 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:34 DR:47 LR:-217.9 LO:217.9);ALT=A]chr2:226860379];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	226860092	-	chr2	226864447	+	.	49	47	1725315_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTAAGACT;MAPQ=60;MATEID=1725315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_226845501_226870501_219C;SPAN=4355;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:76 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:47 DR:49 LR:-237.7 LO:237.7);ALT=[chr2:226864447[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
