chr18	63723838	+	chr18	63732362	+	.	93	66	6656441_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AGATTGC;MAPQ=60;MATEID=6656441_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_18_63700001_63725001_171C;SPAN=8524;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:31 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:66 DR:93 LR:-399.4 LO:399.4);ALT=C[chr18:63732362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	63907136	+	chr18	63911761	+	GGTTTTATTTA	60	33	6656705_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;INSERTION=GGTTTTATTTA;MAPQ=0;MATEID=6656705_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_63896001_63921001_212C;SPAN=4625;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:44 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:33 DR:60 LR:-234.4 LO:234.4);ALT=C[chr18:63911761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	64219707	+	chr18	64221254	+	.	56	40	6657396_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTTT;MAPQ=60;MATEID=6657396_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_18_64214501_64239501_190C;SPAN=1547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:44 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:40 DR:56 LR:-227.8 LO:227.8);ALT=T[chr18:64221254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
