chr1	174232543	+	chr1	174073192	+	.	62	46	643211_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=643211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_174219501_174244501_43C;SPAN=159351;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:62 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:46 DR:62 LR:-257.5 LO:257.5);ALT=]chr1:174232543]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	174796560	+	chr1	174801845	+	.	75	59	645743_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=645743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_174783001_174808001_322C;SPAN=5285;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:104 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:59 DR:75 LR:-307.0 LO:307.0);ALT=G[chr1:174801845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
