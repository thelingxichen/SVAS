chr3	176166428	+	chr3	175733328	+	.	20	0	1802624_1	59.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1802624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:175733328(-)-3:176166428(+)__3_176155001_176180001D;SPAN=433100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:14 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:20 LR:-59.41 LO:59.41);ALT=]chr3:176166428]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	175733467	+	chr3	176166530	+	.	12	0	1802625_1	26.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1802625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:175733467(+)-3:176166530(-)__3_176155001_176180001D;SPAN=433063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:47 GQ:26.9 PL:[26.9, 0.0, 86.3] SR:0 DR:12 LR:-26.88 LO:28.66);ALT=A[chr3:176166530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
