chr2	61700774	-	chr2	61703160	+	.	58	19	1035376_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCCCAGCTACTGGGGAGGCTGAGG;MAPQ=60;MATEID=1035376_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_61691001_61716001_188C;SPAN=2386;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:72 DP:106 GQ:47.3 PL:[209.0, 0.0, 47.3] SR:19 DR:58 LR:-214.6 LO:214.6);ALT=[chr2:61703160[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	61925924	-	chr8	96738679	+	.	2	4	5560114_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=5560114_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_96726001_96751001_384C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:53 GQ:0.9 PL:[0.0, 0.9, 128.7] SR:4 DR:2 LR:1.155 LO:7.245);ALT=[chr8:96738679[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	62844191	-	chr2	62866175	+	.	17	24	1041577_1	83.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AAAAGTCAGGAAACAACAGATGCTGGAGAGGA;MAPQ=60;MATEID=1041577_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_62842501_62867501_510C;SPAN=21984;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:108 GQ:83 PL:[83.0, 0.0, 178.7] SR:24 DR:17 LR:-82.97 LO:84.92);ALT=[chr2:62866175[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	62844312	+	chr2	62866123	-	.	16	16	1041578_1	66.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=AAAAAAAGCTCATCATCACTGCTCATTAGAGAAATGCAAA;MAPQ=60;MATEID=1041578_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_2_62842501_62867501_31C;SPAN=21811;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:107 GQ:66.8 PL:[66.8, 0.0, 192.2] SR:16 DR:16 LR:-66.74 LO:70.15);ALT=T]chr2:62866123];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	63002951	+	chr2	63010274	+	.	69	54	1041937_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGCC;MAPQ=60;MATEID=1041937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62989501_63014501_316C;SPAN=7323;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:83 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:54 DR:69 LR:-307.0 LO:307.0);ALT=C[chr2:63010274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18835664	+	chr8	96265721	+	.	30	0	10201538_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10201538_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:96265721(-)-19:18835664(+)__19_18816001_18841001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:82 GQ:77 PL:[77.0, 0.0, 119.9] SR:0 DR:30 LR:-76.81 LO:77.38);ALT=]chr19:18835664]A;VARTYPE=BND:TRX-th;JOINTYPE=th
