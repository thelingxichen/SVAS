chr6	56757777	-	chr21	18408566	+	.	22	0	4227336_1	52.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4227336_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:56757777(-)-21:18408566(-)__6_56742001_56767001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:75 GQ:52.4 PL:[52.4, 0.0, 128.3] SR:0 DR:22 LR:-52.3 LO:54.12);ALT=[chr21:18408566[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	56758363	+	chr6	56760947	+	.	102	75	4227342_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CCTACTTTTAGTTCTTT;MAPQ=0;MATEID=4227342_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TTT;SCTG=c_6_56742001_56767001_113C;SECONDARY;SPAN=2584;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:172 DP:751 GQ:99 PL:[364.6, 0.0, 1457.0] SR:75 DR:102 LR:-364.3 LO:401.4);ALT=T[chr6:56760947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	56761005	+	chr21	18408584	-	.	15	53	4227349_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=4227349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_56742001_56767001_46C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:81 GQ:31.1 PL:[163.1, 0.0, 31.1] SR:53 DR:15 LR:-167.7 LO:167.7);ALT=T]chr21:18408584];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	57284911	+	chr6	57289366	+	TTACAGCTTCG	40	73	4229382_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TTACAGCTTCG;MAPQ=60;MATEID=4229382_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_6_57281001_57306001_532C;SPAN=4455;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:107 DP:186 GQ:99 PL:[302.9, 0.0, 147.8] SR:73 DR:40 LR:-305.7 LO:305.7);ALT=T[chr6:57289366[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	57572700	+	chr6	57585284	-	.	24	0	4231222_1	59.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=4231222_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:57572700(+)-6:57585284(+)__6_57575001_57600001D;SPAN=12584;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:72 GQ:59.9 PL:[59.9, 0.0, 112.7] SR:0 DR:24 LR:-59.72 LO:60.68);ALT=C]chr6:57585284];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	57572822	-	chr6	57585123	+	.	18	0	4231223_1	40.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=4231223_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:57572822(-)-6:57585123(-)__6_57575001_57600001D;SPAN=12301;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:72 GQ:40.1 PL:[40.1, 0.0, 132.5] SR:0 DR:18 LR:-39.91 LO:42.8);ALT=[chr6:57585123[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	58076948	+	chr6	62128256	-	.	10	0	4237289_1	20.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=4237289_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:58076948(+)-6:62128256(+)__6_62107501_62132501D;SPAN=4051308;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=A]chr6:62128256];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	58360885	+	chr6	58362626	-	.	12	0	4234161_1	5.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=4234161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:58360885(+)-6:58362626(+)__6_58359001_58384001D;SPAN=1741;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:128 GQ:5 PL:[5.0, 0.0, 305.3] SR:0 DR:12 LR:-4.934 LO:22.91);ALT=A]chr6:58362626];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	61897088	+	chr6	61896042	+	.	4	9	4236600_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAGAATGCTTCTGTCTAGTTTT;MAPQ=60;MATEID=4236600_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_61887001_61912001_280C;SPAN=1046;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:132 GQ:7.4 PL:[7.4, 0.0, 311.0] SR:9 DR:4 LR:-7.151 LO:25.12);ALT=]chr6:61897088]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	61928298	-	chr6	61931261	+	.	8	0	4236751_1	0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=4236751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:61928298(-)-6:61931261(-)__6_61911501_61936501D;SPAN=2963;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:123 GQ:6.6 PL:[0.0, 6.6, 310.2] SR:0 DR:8 LR:6.916 LO:13.95);ALT=[chr6:61931261[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr21	18457512	+	chr21	21822281	+	.	0	23	10715672_1	66.0	.	EVDNC=ASSMB;HOMSEQ=ATATATATATATATATATATATATA;MAPQ=60;MATEID=10715672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_18448501_18473501_42C;SPAN=3364769;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:23 DP:6 GQ:6 PL:[66.0, 6.0, 0.0] SR:23 DR:0 LR:-66.02 LO:66.02);ALT=A[chr21:21822281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	18612332	+	chr21	18613634	+	.	100	73	10715746_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATA;MAPQ=60;MATEID=10715746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_18595501_18620501_45C;SPAN=1302;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:25 GQ:36 PL:[396.0, 36.0, 0.0] SR:73 DR:100 LR:-396.1 LO:396.1);ALT=A[chr21:18613634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
