chr4	172374412	+	chr4	172379426	+	.	106	66	2336957_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2336957_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_4_172357501_172382501_108C;SPAN=5014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:141 DP:33 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:66 DR:106 LR:-415.9 LO:415.9);ALT=G[chr4:172379426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	172988639	+	chr4	172992932	+	C	117	85	2338459_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=2338459_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_4_172970001_172995001_250C;SPAN=4293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:42 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:85 DR:117 LR:-452.2 LO:452.2);ALT=A[chr4:172992932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	173425032	+	chr4	173433521	+	A	39	36	2339837_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=2339837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_173411001_173436001_306C;SPAN=8489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:67 GQ:18 PL:[198.0, 18.0, 0.0] SR:36 DR:39 LR:-198.0 LO:198.0);ALT=A[chr4:173433521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	174254399	+	chr4	174255426	+	.	26	0	2342496_1	56.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2342496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:174254399(+)-4:174255426(-)__4_174244001_174269001D;SPAN=1027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:107 GQ:56.9 PL:[56.9, 0.0, 202.1] SR:0 DR:26 LR:-56.84 LO:61.44);ALT=A[chr4:174255426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	174533067	+	chr4	174535912	+	.	32	31	2343835_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=ACTTTAAA;MAPQ=0;MATEID=2343835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_174513501_174538501_363C;SECONDARY;SPAN=2845;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:56 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:31 DR:32 LR:-178.2 LO:178.2);ALT=T[chr4:174535912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
