chr10	69321659	+	chr10	69341590	-	.	30	0	6330546_1	86.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6330546_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:69321659(+)-10:69341590(+)__10_69335001_69360001D;SPAN=19931;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:46 GQ:23.9 PL:[86.6, 0.0, 23.9] SR:0 DR:30 LR:-88.45 LO:88.45);ALT=A]chr10:69341590];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	70126353	+	chr10	70127381	-	.	9	0	6334191_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6334191_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:70126353(+)-10:70127381(+)__10_70119001_70144001D;SPAN=1028;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:114 GQ:0.9 PL:[0.0, 0.9, 277.2] SR:0 DR:9 LR:1.176 LO:16.48);ALT=G]chr10:70127381];VARTYPE=BND:INV-hh;JOINTYPE=hh
