chr13	25156801	-	chr13	25540421	+	.	9	0	5424833_1	17.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5424833_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:25156801(-)-13:25540421(-)__13_25529001_25554001D;SPAN=383620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:0 DR:9 LR:-17.25 LO:20.3);ALT=[chr13:25540421[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	25170039	-	chr13	25527098	+	.	11	6	5424409_1	38.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGAAGGTGCTGAGCAGAC;MAPQ=60;MATEID=5424409_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_25504501_25529501_259C;SPAN=357059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:54 GQ:38.3 PL:[38.3, 0.0, 91.1] SR:6 DR:11 LR:-38.19 LO:39.45);ALT=[chr13:25527098[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	25487230	+	chr13	25496897	+	.	8	4	5424294_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=5424294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_25480001_25505001_359C;SPAN=9667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:4 DR:8 LR:-8.898 LO:19.93);ALT=C[chr13:25496897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
