chr13	26754439	-	chr13	26755462	+	.	12	0	7963360_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7963360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:26754439(-)-13:26755462(-)__13_26729501_26754501D;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:0 DR:12 LR:-20.92 LO:26.38);ALT=[chr13:26755462[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
