chr19	58018448	+	chr19	58005436	+	.	3	2	10390743_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCACACTGGAGAAA;MAPQ=60;MATEID=10390743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_57991501_58016501_34C;SPAN=13012;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:2 DR:3 LR:6.844 LO:6.647);ALT=]chr19:58018448]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	58934311	-	chr19	58935465	+	.	9	0	10395208_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=10395208_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:58934311(-)-19:58935465(-)__19_58922501_58947501D;SPAN=1154;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:162 GQ:13.9 PL:[0.0, 13.9, 419.2] SR:0 DR:9 LR:14.18 LO:15.07);ALT=[chr19:58935465[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
