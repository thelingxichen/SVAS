chrX	152087627	+	chrX	152088870	+	.	2	3	7557121_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=7557121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_152071501_152096501_123C;SPAN=1243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:43 GQ:1.7 PL:[1.7, 0.0, 100.7] SR:3 DR:2 LR:-1.554 LO:7.624);ALT=T[chrX:152088870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152655501	+	chrX	152648071	+	.	29	0	7558583_1	50.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7558583_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:152648071(-)-23:152655501(+)__23_152635001_152660001D;SPAN=7430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:167 GQ:50.6 PL:[50.6, 0.0, 354.2] SR:0 DR:29 LR:-50.49 LO:63.73);ALT=]chrX:152655501]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	152713369	+	chrX	152719852	+	.	0	19	7558097_1	47.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7558097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_152708501_152733501_274C;SPAN=6483;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:55 GQ:47.9 PL:[47.9, 0.0, 84.2] SR:19 DR:0 LR:-47.82 LO:48.41);ALT=T[chrX:152719852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152734721	+	chrX	152735907	+	.	0	7	7558026_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7558026_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_152733001_152758001_142C;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=T[chrX:152735907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152966433	+	chrX	152967461	+	.	0	8	7558703_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=7558703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_152953501_152978501_248C;SPAN=1028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:8 DR:0 LR:-12.05 LO:17.05);ALT=G[chrX:152967461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152969532	+	chrX	152981001	+	.	8	0	7558710_1	18.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7558710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:152969532(+)-23:152981001(-)__23_152953501_152978501D;SPAN=11469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:0 DR:8 LR:-18.55 LO:19.42);ALT=A[chrX:152981001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152981145	+	chrX	152986327	+	.	3	38	7558469_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7558469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_152978001_153003001_175C;SPAN=5182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:86 GQ:95.6 PL:[112.1, 0.0, 95.6] SR:38 DR:3 LR:-112.1 LO:112.1);ALT=C[chrX:152986327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152981197	+	chrX	152989749	+	.	17	0	7558470_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7558470_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:152981197(+)-23:152989749(-)__23_152978001_153003001D;SPAN=8552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:0 DR:17 LR:-42.84 LO:43.35);ALT=T[chrX:152989749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152986429	+	chrX	152989788	+	TTTAGGAGAAATGAAGGGAATGCAGAGAAGCAACACAACAAAGACCTCCGCATAGAGGAAGGTGGCAACTGCAGTCCACTGCAGACTCATCCTGTTGCTAGAAGGTTTCCCACAGGAAGATGTGAGCTTGTTT	63	91	7558487_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TTTAGGAGAAATGAAGGGAATGCAGAGAAGCAACACAACAAAGACCTCCGCATAGAGGAAGGTGGCAACTGCAGTCCACTGCAGACTCATCCTGTTGCTAGAAGGTTTCCCACAGGAAGATGTGAGCTTGTTT;MAPQ=60;MATEID=7558487_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_152978001_153003001_167C;SPAN=3359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:83 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:91 DR:63 LR:-340.0 LO:340.0);ALT=T[chrX:152989788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152986476	+	chrX	152988699	+	.	12	0	7558488_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7558488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:152986476(+)-23:152988699(-)__23_152978001_153003001D;SPAN=2223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:63 GQ:22.7 PL:[22.7, 0.0, 128.3] SR:0 DR:12 LR:-22.54 LO:26.91);ALT=G[chrX:152988699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	152988744	+	chrX	152989788	+	.	62	15	7558494_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=7558494_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_23_152978001_153003001_167C;SPAN=1044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:75 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:15 DR:62 LR:-221.2 LO:221.2);ALT=C[chrX:152989788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153055329	+	chrX	153059704	+	.	15	0	7558845_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7558845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153055329(+)-23:153059704(-)__23_153051501_153076501D;SPAN=4375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:0 DR:15 LR:-35.16 LO:36.62);ALT=C[chrX:153059704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153055802	+	chrX	153059725	+	.	31	0	7558851_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7558851_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153055802(+)-23:153059725(-)__23_153051501_153076501D;SPAN=3923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:46 GQ:20.6 PL:[89.9, 0.0, 20.6] SR:0 DR:31 LR:-92.19 LO:92.19);ALT=T[chrX:153059725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153056368	+	chrX	153059734	+	.	15	0	7558854_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7558854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153056368(+)-23:153059734(-)__23_153051501_153076501D;SPAN=3366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:0 DR:15 LR:-31.91 LO:35.06);ALT=G[chrX:153059734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153060209	+	chrX	153063177	+	CCGAGGCCTGCCTGGAGCCCCAGATCACCCCTTCCTACTACACCACTTCTGACGCTGTCATTTCCACTGAGACCGTCTTCATTGTGGAGATCTCCCTGACATGCAAGAACAGGGTCCAGAACATGGCTCTCTATGCTGACGTCGGTGGAAAACAATTCCCTGTCACTCGAGGCCAGGATGTGGGGCGTTAT	0	122	7558862_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGGTG;INSERTION=CCGAGGCCTGCCTGGAGCCCCAGATCACCCCTTCCTACTACACCACTTCTGACGCTGTCATTTCCACTGAGACCGTCTTCATTGTGGAGATCTCCCTGACATGCAAGAACAGGGTCCAGAACATGGCTCTCTATGCTGACGTCGGTGGAAAACAATTCCCTGTCACTCGAGGCCAGGATGTGGGGCGTTAT;MAPQ=60;MATEID=7558862_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_153051501_153076501_158C;SPAN=2968;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:100 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:122 DR:0 LR:-359.8 LO:359.8);ALT=G[chrX:153063177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153060214	+	chrX	153061956	+	.	53	0	7558863_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7558863_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153060214(+)-23:153061956(-)__23_153051501_153076501D;SPAN=1742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:201 GQ:99 PL:[120.7, 0.0, 365.0] SR:0 DR:53 LR:-120.5 LO:127.5);ALT=C[chrX:153061956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153060214	+	chrX	153062938	+	.	18	0	7558864_1	5.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7558864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153060214(+)-23:153062938(-)__23_153051501_153076501D;SPAN=2724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:200 GQ:5.2 PL:[5.2, 0.0, 480.5] SR:0 DR:18 LR:-5.233 LO:34.04);ALT=C[chrX:153062938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153187264	+	chrX	153191590	+	.	84	14	7559073_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7559073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_153174001_153199001_134C;SPAN=4326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:47 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:14 DR:84 LR:-267.4 LO:267.4);ALT=T[chrX:153191590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153197885	+	chrX	153199395	+	AATGAGGTGATATGTCCATGGGGCACATCATCTGGGTCCTCTTC	2	26	7559094_1	78.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AATGAGGTGATATGTCCATGGGGCACATCATCTGGGTCCTCTTC;MAPQ=60;MATEID=7559094_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_153174001_153199001_15C;SPAN=1510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:38 GQ:12.8 PL:[78.8, 0.0, 12.8] SR:26 DR:2 LR:-81.48 LO:81.48);ALT=C[chrX:153199395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153197929	+	chrX	153200336	+	.	10	0	7559106_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7559106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153197929(+)-23:153200336(-)__23_153198501_153223501D;SPAN=2407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:0 DR:10 LR:-26.78 LO:26.78);ALT=A[chrX:153200336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153201033	+	chrX	153205555	+	.	0	17	7559115_1	42.0	.	EVDNC=ASSMB;HOMSEQ=CTGG;MAPQ=60;MATEID=7559115_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_153198501_153223501_133C;SPAN=4522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:17 DR:0 LR:-42.57 LO:43.16);ALT=G[chrX:153205555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153205689	+	chrX	153206931	+	.	0	9	7559119_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7559119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_153198501_153223501_255C;SPAN=1242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:9 DR:0 LR:-18.87 LO:20.92);ALT=G[chrX:153206931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153357765	+	chrX	153363060	+	.	11	8	7559405_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7559405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_153345501_153370501_159C;SPAN=5295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:8 DR:11 LR:-39.54 LO:40.27);ALT=C[chrX:153363060[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153633999	+	chrX	153637448	+	.	15	4	7560314_1	40.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7560314_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_153615001_153640001_176C;SPAN=3449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:58 GQ:40.4 PL:[40.4, 0.0, 99.8] SR:4 DR:15 LR:-40.4 LO:41.81);ALT=G[chrX:153637448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153657107	+	chrX	153660173	+	.	9	0	7560358_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7560358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153657107(+)-23:153660173(-)__23_153639501_153664501D;SPAN=3066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:0 DR:9 LR:-14.0 LO:19.3);ALT=G[chrX:153660173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153657200	+	chrX	153660610	+	GACTTGTGGGCTCCTGCGGCCGACACTCATGAAGGCCACATCACCAGCGACTTGCAGCTCTCTACCTACTTAGATCCCGCCCTGGAGCTGGGTCCCAGGAATGTGCTGCTGTTCCTGCAGGACAAGCTGAGCATTGAGGATTTCACAGCATATGGCGGTGTGTTTGGAAACAAGCAGGACAGCGCCTTTTCTAACCTAG	0	64	7560360_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GACTTGTGGGCTCCTGCGGCCGACACTCATGAAGGCCACATCACCAGCGACTTGCAGCTCTCTACCTACTTAGATCCCGCCCTGGAGCTGGGTCCCAGGAATGTGCTGCTGTTCCTGCAGGACAAGCTGAGCATTGAGGATTTCACAGCATATGGCGGTGTGTTTGGAAACAAGCAGGACAGCGCCTTTTCTAACCTAG;MAPQ=60;MATEID=7560360_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_153639501_153664501_244C;SPAN=3410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:78 GQ:1.2 PL:[191.4, 1.2, 0.0] SR:64 DR:0 LR:-202.1 LO:202.1);ALT=G[chrX:153660610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153665594	+	chrX	153666868	+	.	8	0	7560510_1	14.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7560510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153665594(+)-23:153666868(-)__23_153664001_153689001D;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=C[chrX:153666868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153672694	+	chrX	153673979	+	.	41	35	7560522_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7560522_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_153664001_153689001_87C;SPAN=1285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:50 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:35 DR:41 LR:-171.6 LO:171.6);ALT=G[chrX:153673979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153763602	+	chrX	153774250	+	TGAAGAAGGGCTCACTCTGTTTGCGGATGTCAGCCACTGTGAGGCGGGAACGGGCATAGCCCACGATGAAGGTGTTTTCGGGCAGAAGGCCATCCCGGAACAGCCACCAGATGGTGGGGTAGATCTTCTTCTTGGCCAGGTCAC	0	37	7560612_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGAAGAAGGGCTCACTCTGTTTGCGGATGTCAGCCACTGTGAGGCGGGAACGGGCATAGCCCACGATGAAGGTGTTTTCGGGCAGAAGGCCATCCCGGAACAGCCACCAGATGGTGGGGTAGATCTTCTTCTTGGCCAGGTCAC;MAPQ=60;MATEID=7560612_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_153762001_153787001_54C;SPAN=10648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:61 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:37 DR:0 LR:-107.1 LO:107.1);ALT=T[chrX:153774250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153764453	+	chrX	153775003	+	.	23	0	7560615_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7560615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153764453(+)-23:153775003(-)__23_153762001_153787001D;SPAN=10550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:68 GQ:57.5 PL:[57.5, 0.0, 107.0] SR:0 DR:23 LR:-57.5 LO:58.33);ALT=C[chrX:153775003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153775977	+	chrX	153780200	+	.	9	0	7560627_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7560627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:153775977(+)-23:153780200(-)__23_153762001_153787001D;SPAN=4223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:0 DR:9 LR:-17.25 LO:20.3);ALT=C[chrX:153780200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153991256	+	chrX	153993719	+	TAATTATTTTGCCAAAGAAACATAAGAAGAAAAAGGAGCGGAAGTCATTGCCAGAAGAAGATGTAGCC	8	12	7561004_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TAATTATTTTGCCAAAGAAACATAAGAAGAAAAAGGAGCGGAAGTCATTGCCAGAAGAAGATGTAGCC;MAPQ=60;MATEID=7561004_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_153982501_154007501_264C;SPAN=2463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:57 GQ:37.4 PL:[37.4, 0.0, 100.1] SR:12 DR:8 LR:-37.37 LO:38.99);ALT=G[chrX:153993719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	153991256	+	chrX	153993172	+	.	5	5	7561003_1	10.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=7561003_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_23_153982501_154007501_264C;SPAN=1916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:5 DR:5 LR:-10.69 LO:16.71);ALT=G[chrX:153993172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154001525	+	chrX	154003467	+	CAAGTCAGAAGAAGCTGATGATCAAGCAGGGCCTTCTGGACAAGCATGGGAAGCCCACAGACAGCACACCTGCCACCTGGAAGCAGGAGTATGTTGACTA	3	21	7561022_1	54.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=CAAGTCAGAAGAAGCTGATGATCAAGCAGGGCCTTCTGGACAAGCATGGGAAGCCCACAGACAGCACACCTGCCACCTGGAAGCAGGAGTATGTTGACTA;MAPQ=60;MATEID=7561022_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_153982501_154007501_113C;SPAN=1942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:54 GQ:54.8 PL:[54.8, 0.0, 74.6] SR:21 DR:3 LR:-54.69 LO:54.89);ALT=G[chrX:154003467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154019345	+	chrX	154020416	+	TGTCTATGGATCATGCCACCATGAAGAATTCTGGCCACCGTACAGGACTGTTTTTCATTCAGCTTCAGAGTGATTC	3	23	7561067_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TGTCTATGGATCATGCCACCATGAAGAATTCTGGCCACCGTACAGGACTGTTTTTCATTCAGCTTCAGAGTGATTC;MAPQ=60;MATEID=7561067_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_154007001_154032001_186C;SPAN=1071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:81 GQ:57.5 PL:[57.5, 0.0, 136.7] SR:23 DR:3 LR:-57.28 LO:59.17);ALT=T[chrX:154020416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154020169	+	chrX	154033579	+	.	9	0	7561097_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7561097_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154020169(+)-23:154033579(-)__23_154031501_154056501D;SPAN=13410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=T[chrX:154033579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154020562	+	chrX	154033546	+	.	0	41	7561098_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7561098_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_154031501_154056501_163C;SPAN=12984;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:33 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:41 DR:0 LR:-118.8 LO:118.8);ALT=T[chrX:154033546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154444834	+	chrX	154455512	+	.	11	0	7561759_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7561759_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154444834(+)-23:154455512(-)__23_154423501_154448501D;SPAN=10678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:32 GQ:27.8 PL:[27.8, 0.0, 47.6] SR:0 DR:11 LR:-27.64 LO:28.0);ALT=T[chrX:154455512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154444848	+	chrX	154448458	+	.	33	0	7561682_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7561682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154444848(+)-23:154448458(-)__23_154448001_154473001D;SPAN=3610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:26 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:0 DR:33 LR:-95.72 LO:95.72);ALT=T[chrX:154448458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154444853	+	chrX	154456666	+	AAGATGTAGATTCCTTCATGAAACAGCCTGGGAATGAGACTGCAGATACAGTATTAAAGAAGCTGGATGAACAGTACCAGAAGTATAAGTTTATGGAACTCAACCTTGCTCAAAAGAAAAGAAGGCTAAAAGGTCAGATTCCTGAAATTAAACAGACTTTGGAAATTCTAAAATACATGCAGAAGAAAAAA	4	15	7561761_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AAGATGTAGATTCCTTCATGAAACAGCCTGGGAATGAGACTGCAGATACAGTATTAAAGAAGCTGGATGAACAGTACCAGAAGTATAAGTTTATGGAACTCAACCTTGCTCAAAAGAAAAGAAGGCTAAAAGGTCAGATTCCTGAAATTAAACAGACTTTGGAAATTCTAAAATACATGCAGAAGAAAAAA;MAPQ=60;MATEID=7561761_2;MATENM=1;NM=0;NUMPARTS=4;SCTG=c_23_154423501_154448501_143C;SPAN=11813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:34 GQ:37.1 PL:[43.7, 0.0, 37.1] SR:15 DR:4 LR:-43.62 LO:43.62);ALT=G[chrX:154456666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154448585	+	chrX	154456666	+	CTAAAAGGTCAGATTCCTGAAATTAAACAGACTTTGGAAATTCTAAAATACATGCAGAAGAAAAAA	0	34	7561686_1	96.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTAAAAGGTCAGATTCCTGAAATTAAACAGACTTTGGAAATTCTAAAATACATGCAGAAGAAAAAA;MAPQ=60;MATEID=7561686_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_23_154448001_154473001_38C;SPAN=8081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:59 GQ:46.7 PL:[96.2, 0.0, 46.7] SR:34 DR:0 LR:-97.17 LO:97.17);ALT=G[chrX:154456666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	154774962	+	chrX	154842507	+	.	14	0	7562176_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7562176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154774962(+)-23:154842507(-)__23_154840001_154865001D;SPAN=67545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:37 GQ:36.2 PL:[36.2, 0.0, 52.7] SR:0 DR:14 LR:-36.19 LO:36.38);ALT=T[chrX:154842507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	155216658	+	chrX	155033244	+	.	20	0	7562837_1	57.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=7562837_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:155033244(-)-23:155216658(+)__23_155207501_155232501D;SPAN=183414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:31 GQ:14.9 PL:[57.8, 0.0, 14.9] SR:0 DR:20 LR:-58.8 LO:58.8);ALT=]chrX:155216658]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	155033271	+	chrX	155213887	+	.	31	0	7562838_1	91.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=7562838_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:155033271(+)-23:155213887(-)__23_155207501_155232501D;SPAN=180616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:39 GQ:2.6 PL:[91.7, 0.0, 2.6] SR:0 DR:31 LR:-96.83 LO:96.83);ALT=C[chrX:155213887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	155111110	+	chrX	155119115	+	.	9	0	7562525_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7562525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:155111110(+)-23:155119115(-)__23_155109501_155134501D;SPAN=8005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:0 DR:9 LR:-14.27 LO:19.37);ALT=A[chrX:155119115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
