chr6	5037249	+	chr6	5039187	+	AAAATCTGCTTC	0	75	3998391_1	99.0	.	EVDNC=ASSMB;INSERTION=AAAATCTGCTTC;MAPQ=60;MATEID=3998391_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_5022501_5047501_101C;SPAN=1938;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:40 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:75 DR:0 LR:-221.2 LO:221.2);ALT=T[chr6:5039187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
