chr2	239500398	+	chr2	239501733	+	.	58	39	1778960_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAT;MAPQ=60;MATEID=1778960_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_239487501_239512501_332C;SPAN=1335;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:85 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:39 DR:58 LR:-257.5 LO:257.5);ALT=T[chr2:239501733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
