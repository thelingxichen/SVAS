chr14	65360396	+	chr14	65363541	+	.	67	53	8560754_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAATTTTC;MAPQ=60;MATEID=8560754_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_65341501_65366501_420C;SPAN=3145;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:88 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:53 DR:67 LR:-270.7 LO:270.7);ALT=C[chr14:65363541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65842187	+	chr14	65843223	-	.	19	0	8563178_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=8563178_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65842187(+)-14:65843223(+)__14_65831501_65856501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:113 GQ:32.3 PL:[32.3, 0.0, 240.2] SR:0 DR:19 LR:-32.1 LO:41.46);ALT=A]chr14:65843223];VARTYPE=BND:INV-hh;JOINTYPE=hh
