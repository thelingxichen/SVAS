chr16	77756514	+	chr16	77759326	+	.	3	2	6255550_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6255550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_77738501_77763501_262C;SPAN=2812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:67 GQ:4.8 PL:[0.0, 4.8, 171.6] SR:2 DR:3 LR:4.948 LO:6.824);ALT=G[chr16:77759326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78371638	+	chr16	78384899	+	.	51	49	6256618_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6256618_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_78375501_78400501_60C;SPAN=13261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:9 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:49 DR:51 LR:-234.4 LO:234.4);ALT=A[chr16:78384899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	78928639	+	chr16	79095001	+	.	27	17	6257609_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATTGGG;MAPQ=60;MATEID=6257609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_79086001_79111001_207C;SPAN=166362;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:17 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:17 DR:27 LR:-105.6 LO:105.6);ALT=G[chr16:79095001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
