chr7	106820507	+	chr7	106822817	+	.	0	7	3511528_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3511528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_106820001_106845001_340C;SPAN=2310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:104 GQ:4.8 PL:[0.0, 4.8, 260.7] SR:7 DR:0 LR:5.069 LO:12.32);ALT=G[chr7:106822817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107220800	+	chr7	107224324	+	.	21	0	3512676_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3512676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:107220800(+)-7:107224324(-)__7_107212001_107237001D;SPAN=3524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:73 GQ:49.7 PL:[49.7, 0.0, 125.6] SR:0 DR:21 LR:-49.54 LO:51.45);ALT=C[chr7:107224324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107221309	+	chr7	107224325	+	.	2	13	3512678_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3512678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_107212001_107237001_214C;SPAN=3016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:80 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:13 DR:2 LR:-24.54 LO:30.82);ALT=G[chr7:107224325[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107531734	+	chr7	107542183	+	AGAGGCCATTTCAATCGAATATCTCATGGCCTACAGGGACTTTCTGCAGTGCCTCTGAGAACTTACGCAGATCAGCCGA	9	19	3513935_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGAGGCCATTTCAATCGAATATCTCATGGCCTACAGGGACTTTCTGCAGTGCCTCTGAGAACTTACGCAGATCAGCCGA;MAPQ=60;MATEID=3513935_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_107530501_107555501_172C;SPAN=10449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:126 GQ:35.3 PL:[35.3, 0.0, 269.6] SR:19 DR:9 LR:-35.18 LO:45.74);ALT=G[chr7:107542183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107531734	+	chr7	107533643	+	.	10	6	3513934_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3513934_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_107530501_107555501_172C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:117 GQ:8 PL:[8.0, 0.0, 275.3] SR:6 DR:10 LR:-7.914 LO:23.41);ALT=G[chr7:107533643[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107531768	+	chr7	107542767	+	.	9	0	3513936_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3513936_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:107531768(+)-7:107542767(-)__7_107530501_107555501D;SPAN=10999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:137 GQ:7.2 PL:[0.0, 7.2, 346.5] SR:0 DR:9 LR:7.408 LO:15.74);ALT=A[chr7:107542767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	107556141	+	chr7	107557239	+	.	3	6	3513860_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3513860_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_107555001_107580001_139C;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:108 GQ:9.3 PL:[0.0, 9.3, 280.5] SR:6 DR:3 LR:9.454 LO:10.04);ALT=C[chr7:107557239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85211624	+	chr7	107829249	+	.	14	43	3515475_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TAAA;MAPQ=60;MATEID=3515475_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_107824501_107849501_349C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:61 GQ:3.5 PL:[142.1, 0.0, 3.5] SR:43 DR:14 LR:-149.4 LO:149.4);ALT=]chr11:85211624]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	85217464	-	chr11	86255084	+	.	36	0	4947110_1	99.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=4947110_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85217464(-)-11:86255084(-)__11_86240001_86265001D;SPAN=1037620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:5 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=[chr11:86255084[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	85217696	+	chr11	86254971	-	.	31	0	4947111_1	89.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=4947111_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85217696(+)-11:86254971(+)__11_86240001_86265001D;SPAN=1037275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:10 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=T]chr11:86254971];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	85339729	+	chr11	85345127	+	.	12	0	4944464_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4944464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85339729(+)-11:85345127(-)__11_85333501_85358501D;SPAN=5398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:0 DR:12 LR:-15.23 LO:24.87);ALT=C[chr11:85345127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85339729	+	chr11	85342727	+	.	9	0	4944463_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4944463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85339729(+)-11:85342727(-)__11_85333501_85358501D;SPAN=2998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:96 GQ:3.8 PL:[3.8, 0.0, 228.2] SR:0 DR:9 LR:-3.7 LO:17.19);ALT=C[chr11:85342727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85339733	+	chr11	85342187	+	.	34	3	4944465_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4944465_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_85333501_85358501_191C;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:102 GQ:84.8 PL:[84.8, 0.0, 160.7] SR:3 DR:34 LR:-84.6 LO:85.96);ALT=G[chr11:85342187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85342853	+	chr11	85345130	+	.	0	12	4944469_1	18.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4944469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_85333501_85358501_260C;SPAN=2277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:12 DR:0 LR:-18.21 LO:25.61);ALT=G[chr11:85345130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85359134	+	chr11	85365105	+	.	53	7	4944572_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4944572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_85358001_85383001_186C;SPAN=5971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:67 GQ:8.1 PL:[178.2, 8.1, 0.0] SR:7 DR:53 LR:-182.6 LO:182.6);ALT=G[chr11:85365105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85359134	+	chr11	85361289	+	.	11	8	4944570_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TAAGG;MAPQ=60;MATEID=4944570_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_85358001_85383001_343C;SPAN=2155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:70 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:8 DR:11 LR:-30.55 LO:34.51);ALT=G[chr11:85361289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85361386	+	chr11	85365105	+	.	3	14	4944576_1	36.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=4944576_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_85358001_85383001_343C;SPAN=3719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:73 GQ:36.5 PL:[36.5, 0.0, 138.8] SR:14 DR:3 LR:-36.34 LO:39.81);ALT=G[chr11:85365105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85365302	+	chr11	85366636	+	.	0	8	4944590_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=4944590_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_85358001_85383001_338C;SPAN=1334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:81 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:8 DR:0 LR:-4.463 LO:15.47);ALT=T[chr11:85366636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	85550690	-	chr11	85552115	+	.	11	0	4945086_1	19.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4945086_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:85550690(-)-11:85552115(-)__11_85529501_85554501D;SPAN=1425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=[chr11:85552115[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	86013523	+	chr11	86017286	+	.	0	23	4946200_1	43.0	.	EVDNC=ASSMB;HOMSEQ=GGTG;MAPQ=60;MATEID=4946200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_85995001_86020001_121C;SPAN=3763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:122 GQ:43.1 PL:[43.1, 0.0, 251.0] SR:23 DR:0 LR:-42.87 LO:51.46);ALT=G[chr11:86017286[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
