chr5	52394499	+	chr5	52396240	+	.	5	3	2471121_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2471121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_52381001_52406001_211C;SPAN=1741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:55 GQ:5 PL:[5.0, 0.0, 127.1] SR:3 DR:5 LR:-4.905 LO:11.87);ALT=T[chr5:52396240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	52403052	+	chr5	52404352	+	.	0	7	2471141_1	9.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2471141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_52381001_52406001_240C;SPAN=1300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:51 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:7 DR:0 LR:-9.29 LO:14.6);ALT=C[chr5:52404352[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	52403084	+	chr5	52405538	+	.	8	0	2471148_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2471148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:52403084(+)-5:52405538(-)__5_52405501_52430501D;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=A[chr5:52405538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	52856570	+	chr5	52942059	+	.	25	0	2471820_1	75.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2471820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:52856570(+)-5:52942059(-)__5_52920001_52945001D;SPAN=85489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:31 GQ:1.5 PL:[75.9, 1.5, 0.0] SR:0 DR:25 LR:-78.48 LO:78.48);ALT=C[chr5:52942059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	52856592	+	chr5	52899279	+	.	16	12	2471852_1	65.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CAGGT;MAPQ=60;MATEID=2471852_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_5_52895501_52920501_41C;SPAN=42687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:28 GQ:2.3 PL:[65.0, 0.0, 2.3] SR:12 DR:16 LR:-68.45 LO:68.45);ALT=T[chr5:52899279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
