chr5	121576131	+	chr5	121580809	+	.	49	36	2568386_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGAGATACAATTTCA;MAPQ=60;MATEID=2568386_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_5_121569001_121594001_83C;SPAN=4678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:27 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:36 DR:49 LR:-188.1 LO:188.1);ALT=A[chr5:121580809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122110906	+	chr5	122135385	+	TCAAGTCCATCATCTCCAGAACCAGCTAGTCTTCCTGCAGAAGATATTAGTGCAAACTCCAATGGCCCAAAACCCACAGAAGTTGTATTAGATGATGACAGAGAAGATCTTTTTGC	26	55	2569054_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TCAAGTCCATCATCTCCAGAACCAGCTAGTCTTCCTGCAGAAGATATTAGTGCAAACTCCAATGGCCCAAAACCCACAGAAGTTGTATTAGATGATGACAGAGAAGATCTTTTTGC;MAPQ=60;MATEID=2569054_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_122132501_122157501_17C;SPAN=24479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:32 GQ:18 PL:[198.0, 18.0, 0.0] SR:55 DR:26 LR:-198.0 LO:198.0);ALT=G[chr5:122135385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122110906	+	chr5	122130959	+	.	47	18	2568953_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2568953_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_5_122108001_122133001_195C;SPAN=20053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:67 GQ:11.6 PL:[150.2, 0.0, 11.6] SR:18 DR:47 LR:-157.1 LO:157.1);ALT=G[chr5:122130959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122154719	+	chr5	122161745	+	.	6	8	2569094_1	29.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2569094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_122132501_122157501_82C;SPAN=7026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:25 GQ:29.6 PL:[29.6, 0.0, 29.6] SR:8 DR:6 LR:-29.54 LO:29.54);ALT=G[chr5:122161745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122161888	+	chr5	122165289	+	TGGGAGGCGAAAGTGCAACAAGGGGAAAGAGATTTTGAACAGATATCTAAAACGATTCGAAAAGAAGTGGGAAGATTTGAGAAAGAACGAGTGAAGGATTTTAAAACCGTTATCATCAAGTACTTAGAATCACTAGTTCAAACACAACA	0	21	2568999_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACAG;INSERTION=TGGGAGGCGAAAGTGCAACAAGGGGAAAGAGATTTTGAACAGATATCTAAAACGATTCGAAAAGAAGTGGGAAGATTTGAGAAAGAACGAGTGAAGGATTTTAAAACCGTTATCATCAAGTACTTAGAATCACTAGTTCAAACACAACA;MAPQ=60;MATEID=2568999_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_122157001_122182001_195C;SPAN=3401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:47 GQ:56.6 PL:[56.6, 0.0, 56.6] SR:21 DR:0 LR:-56.59 LO:56.59);ALT=G[chr5:122165289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122163341	+	chr5	122165289	+	.	2	11	2569002_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACAG;MAPQ=60;MATEID=2569002_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_122157001_122182001_195C;SPAN=1948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:11 DR:2 LR:-28.83 LO:30.91);ALT=G[chr5:122165289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	122582810	+	chr9	40135784	+	.	3	32	2570062_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAATG;MAPQ=60;MATEID=2570062_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_122573501_122598501_63C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:23 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:32 DR:3 LR:-95.72 LO:95.72);ALT=G[chr9:40135784[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	123013680	+	chr5	123696644	-	.	16	0	2571224_1	44.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=2571224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:123013680(+)-5:123696644(+)__5_123676001_123701001D;SPAN=682964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:30 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:0 DR:16 LR:-44.89 LO:44.89);ALT=G]chr5:123696644];VARTYPE=BND:INV-hh;JOINTYPE=hh
