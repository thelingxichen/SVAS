chr10	20011418	+	chr10	20017385	+	.	10	0	4535013_1	23.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4535013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:20011418(+)-10:20017385(-)__10_19992001_20017001D;SPAN=5967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=C[chr10:20017385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	20106120	+	chr10	20290703	+	.	4	2	4535682_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4535682_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_20286001_20311001_118C;SPAN=184583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:39 GQ:5.9 PL:[5.9, 0.0, 88.4] SR:2 DR:4 LR:-5.939 LO:10.27);ALT=G[chr10:20290703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
