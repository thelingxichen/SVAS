chr4	142230783	+	chr4	142233063	+	.	67	51	2958275_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGCC;MAPQ=60;MATEID=2958275_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_4_142222501_142247501_302C;SPAN=2280;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:90 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:51 DR:67 LR:-267.4 LO:267.4);ALT=C[chr4:142233063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
