chr18	63766873	+	chr18	63769203	+	.	45	47	10045370_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTGG;MAPQ=60;MATEID=10045370_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_18_63749001_63774001_100C;SPAN=2330;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:16 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:47 DR:45 LR:-224.5 LO:224.5);ALT=G[chr18:63769203[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
