chr8	17780698	+	chr8	17793095	+	AAACAGCTTTGAAGTGTGGAGCGGGAAAGGAGCAGTTTCTGAGCTGCAAAAACTAGTTTCTAAA	3	30	3764380_1	91.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AAACAGCTTTGAAGTGTGGAGCGGGAAAGGAGCAGTTTCTGAGCTGCAAAAACTAGTTTCTAAA;MAPQ=60;MATEID=3764380_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_17762501_17787501_104C;SPAN=12397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:52 GQ:32.3 PL:[91.7, 0.0, 32.3] SR:30 DR:3 LR:-92.95 LO:92.95);ALT=G[chr8:17793095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17780698	+	chr8	17782220	+	.	11	24	3764379_1	73.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3764379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_17762501_17787501_166C;SPAN=1522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:94 GQ:73.7 PL:[73.7, 0.0, 152.9] SR:24 DR:11 LR:-73.56 LO:75.15);ALT=G[chr8:17782220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17924808	+	chr8	17928809	+	AATTTTTCATCCACCACCTGCATAATTTTTCCACTTGGCACGAATGTATTTATCATATTCTTCAGAGAATTCACTATAACCTTTAG	0	58	3764889_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AATTTTTCATCCACCACCTGCATAATTTTTCCACTTGGCACGAATGTATTTATCATATTCTTCAGAGAATTCACTATAACCTTTAG;MAPQ=60;MATEID=3764889_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_17909501_17934501_246C;SPAN=4001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:91 GQ:51.5 PL:[167.0, 0.0, 51.5] SR:58 DR:0 LR:-170.0 LO:170.0);ALT=C[chr8:17928809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17927388	+	chr8	17928812	+	AT	0	43	3764903_1	99.0	.	EVDNC=ASSMB;INSERTION=AT;MAPQ=60;MATEID=3764903_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_17909501_17934501_111C;SPAN=1424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:101 GQ:99 PL:[114.8, 0.0, 128.0] SR:43 DR:0 LR:-114.6 LO:114.6);ALT=C[chr8:17928812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17927433	+	chr8	17941522	+	.	20	0	3764998_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3764998_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:17927433(+)-8:17941522(-)__8_17934001_17959001D;SPAN=14089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:0 DR:20 LR:-52.2 LO:52.37);ALT=G[chr8:17941522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17928899	+	chr8	17941490	+	GTTGGTCCTGAAGGAGGATAGGTTGATTTTCTGCAGTCCTCTGTCCA	66	66	3765000_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTGGTCCTGAAGGAGGATAGGTTGATTTTCTGCAGTCCTCTGTCCA;MAPQ=60;MATEID=3765000_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_17934001_17959001_372C;SPAN=12591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:49 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:66 DR:66 LR:-277.3 LO:277.3);ALT=C[chr8:17941490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	17933149	+	chr8	17941526	+	.	26	0	3765002_1	71.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3765002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:17933149(+)-8:17941526(-)__8_17934001_17959001D;SPAN=8377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:53 GQ:55.1 PL:[71.6, 0.0, 55.1] SR:0 DR:26 LR:-71.55 LO:71.55);ALT=A[chr8:17941526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	18454620	+	chr8	18455945	+	.	44	28	3766641_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAGGATC;MAPQ=60;MATEID=3766641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_18448501_18473501_189C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:90 GQ:38.3 PL:[180.2, 0.0, 38.3] SR:28 DR:44 LR:-185.5 LO:185.5);ALT=C[chr8:18455945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
