chr18	158714	+	chr18	163307	+	.	11	6	6523552_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6523552_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_147001_172001_225C;SPAN=4593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:6 DR:11 LR:-28.83 LO:30.91);ALT=G[chr18:163307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	657947	+	chr18	659639	+	.	0	47	6524614_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6524614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_637001_662001_301C;SPAN=1692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:59 GQ:3.8 PL:[139.1, 0.0, 3.8] SR:47 DR:0 LR:-146.9 LO:146.9);ALT=G[chr18:659639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	659715	+	chr18	662144	+	.	0	10	6524616_1	24.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6524616_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_637001_662001_204C;SPAN=2429;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:32 GQ:24.5 PL:[24.5, 0.0, 50.9] SR:10 DR:0 LR:-24.34 LO:24.94);ALT=G[chr18:662144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	662355	+	chr18	670689	+	.	11	0	6524721_1	20.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6524721_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:662355(+)-18:670689(-)__18_661501_686501D;SPAN=8334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:0 DR:11 LR:-20.87 LO:24.74);ALT=G[chr18:670689[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	669185	+	chr18	670689	+	.	14	0	6524728_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6524728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:669185(+)-18:670689(-)__18_661501_686501D;SPAN=1504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:63 GQ:29.3 PL:[29.3, 0.0, 121.7] SR:0 DR:14 LR:-29.15 LO:32.46);ALT=C[chr18:670689[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	697356	+	chr18	706470	+	.	0	11	6524664_1	23.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6524664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_686001_711001_280C;SPAN=9114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:11 DR:0 LR:-23.85 LO:25.91);ALT=C[chr18:706470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	706579	+	chr18	712504	+	.	17	6	6524768_1	57.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6524768_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_710501_735501_52C;SPAN=5925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:31 GQ:14.9 PL:[57.8, 0.0, 14.9] SR:6 DR:17 LR:-58.8 LO:58.8);ALT=C[chr18:712504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
