chr7	25057461	+	chr7	25059854	+	.	31	24	3213570_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAAATATATAAAGTC;MAPQ=60;MATEID=3213570_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_25039001_25064001_365C;SPAN=2393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:62 GQ:13.1 PL:[135.2, 0.0, 13.1] SR:24 DR:31 LR:-140.6 LO:140.6);ALT=C[chr7:25059854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	25163747	+	chr7	25164817	+	.	116	0	3214125_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=3214125_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:25163747(+)-7:25164817(-)__7_25161501_25186501D;SPAN=1070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:124 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:0 DR:116 LR:-366.4 LO:366.4);ALT=C[chr7:25164817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	33827299	+	chr7	25164818	+	.	45	0	3813456_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=3813456_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:25164818(-)-8:33827299(+)__8_33810001_33835001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:49 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:45 LR:-145.2 LO:145.2);ALT=]chr8:33827299]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	32680009	+	chr8	32691262	+	.	95	62	3810027_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3810027_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_8_32658501_32683501_291C;SPAN=11253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:130 DP:18 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:62 DR:95 LR:-386.2 LO:386.2);ALT=G[chr8:32691262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	32785602	+	chr8	32899149	+	.	9	0	3810379_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3810379_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:32785602(+)-8:32899149(-)__8_32879001_32904001D;SPAN=113547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=C[chr8:32899149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
