chr6	86623833	+	chr6	86625833	+	CATGGGG	69	38	4312775_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CATGGGG;MAPQ=60;MATEID=4312775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_86607501_86632501_199C;SPAN=2000;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:15 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:38 DR:69 LR:-260.8 LO:260.8);ALT=C[chr6:86625833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	86708754	+	chr6	86714792	+	.	36	50	4313157_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=GTGCCACATTTTCTT;MAPQ=60;MATEID=4313157_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_6_86705501_86730501_164C;SPAN=6038;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:17 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:50 DR:36 LR:-250.9 LO:250.9);ALT=T[chr6:86714792[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
