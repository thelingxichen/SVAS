chr20	13160730	+	chr20	13164100	+	.	44	39	6927654_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTC;MAPQ=60;MATEID=6927654_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_13156501_13181501_132C;SPAN=3370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:68 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:44 LR:-201.3 LO:201.3);ALT=C[chr20:13164100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	13605901	+	chr20	13610579	+	.	0	7	6929076_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6929076_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_13597501_13622501_366C;SPAN=4678;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=T[chr20:13610579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	13878381	-	chr20	13879653	+	.	2	3	6930102_1	0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=GCTGGGATTACAGGCATG;MAPQ=55;MATEID=6930102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_13867001_13892001_67C;SPAN=1272;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:127 GQ:21 PL:[0.0, 21.0, 349.8] SR:3 DR:2 LR:21.2 LO:5.697);ALT=[chr20:13879653[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
