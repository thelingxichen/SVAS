chr5	111066768	+	chr5	111092829	+	.	11	0	2554065_1	30.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=2554065_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:111066768(+)-5:111092829(-)__5_111083001_111108001D;SPAN=26061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:22 GQ:20.6 PL:[30.5, 0.0, 20.6] SR:0 DR:11 LR:-30.4 LO:30.4);ALT=C[chr5:111092829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	111093073	-	chr7	23520284	+	.	10	0	3208710_1	17.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3208710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:111093073(-)-7:23520284(-)__7_23520001_23545001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:0 DR:10 LR:-17.57 LO:22.03);ALT=[chr7:23520284[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	21948126	+	chr7	21951233	+	.	0	7	3201815_1	0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=3201815_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_21927501_21952501_258C;SPAN=3107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:7 DR:0 LR:2.902 LO:12.57);ALT=C[chr7:21951233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	21948127	+	chr7	21956370	+	.	2	3	3201816_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=3201816_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_21927501_21952501_146C;SPAN=8243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:50 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:3 DR:2 LR:-2.959 LO:9.695);ALT=T[chr7:21956370[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	21951374	+	chr7	21956372	+	.	0	11	3201914_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3201914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_21952001_21977001_447C;SPAN=4998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:11 DR:0 LR:-21.68 LO:25.03);ALT=T[chr7:21956372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	21951422	+	chr7	21985435	+	.	9	0	3202006_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3202006_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:21951422(+)-7:21985435(-)__7_21976501_22001501D;SPAN=34013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=A[chr7:21985435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	21956515	+	chr7	21985399	+	.	19	5	3202007_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=3202007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_21976501_22001501_383C;SPAN=28884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:47 GQ:53.3 PL:[53.3, 0.0, 59.9] SR:5 DR:19 LR:-53.29 LO:53.31);ALT=G[chr7:21985399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	22434803	+	chr7	22436761	+	.	76	46	3203661_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=3203661_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_22417501_22442501_173C;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:73 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:46 DR:76 LR:-307.0 LO:307.0);ALT=C[chr7:22436761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23221827	+	chr7	23224687	+	.	8	7	3206417_1	1.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3206417_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_23201501_23226501_304C;SPAN=2860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:117 GQ:1.4 PL:[1.4, 0.0, 281.9] SR:7 DR:8 LR:-1.312 LO:18.67);ALT=T[chr7:23224687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23339227	+	chr7	23340455	+	.	0	4	3207080_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=3207080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_23324001_23349001_348C;SPAN=1228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:118 GQ:18.6 PL:[0.0, 18.6, 323.4] SR:4 DR:0 LR:18.77 LO:5.825);ALT=G[chr7:23340455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23347569	+	chr7	23348974	+	.	0	9	3207323_1	9.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3207323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_23348501_23373501_61C;SPAN=1405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:9 DR:0 LR:-9.119 LO:18.15);ALT=G[chr7:23348974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23556149	+	chr7	23571407	+	GGATTTTGATCTTGATCGAGAATGGGATTCAGAGTGTTTGGAAACCCTTGATGGACTACGAGATCCTGACCTGCTCTCCGATTTTACACGAGCAGGAGTTCCCGTTGGAGATTTTGACTGAGAGCGAGACT	3	15	3208051_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGATTTTGATCTTGATCGAGAATGGGATTCAGAGTGTTTGGAAACCCTTGATGGACTACGAGATCCTGACCTGCTCTCCGATTTTACACGAGCAGGAGTTCCCGTTGGAGATTTTGACTGAGAGCGAGACT;MAPQ=60;MATEID=3208051_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_23544501_23569501_93C;SPAN=15258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:61 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:15 DR:3 LR:-36.29 LO:38.43);ALT=T[chr7:23571407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23561502	+	chr7	23571527	+	.	15	0	3208081_1	35.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3208081_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:23561502(+)-7:23571527(-)__7_23544501_23569501D;SPAN=10025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:50 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.97 LO:37.08);ALT=A[chr7:23571527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	23815639	-	chr7	23838145	+	.	30	0	3209311_1	89.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3209311_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:23815639(-)-7:23838145(-)__7_23838501_23863501D;SPAN=22506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:0 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=[chr7:23838145[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	23815822	+	chr7	23837989	-	.	21	0	3209224_1	45.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=3209224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:23815822(+)-7:23837989(+)__7_23814001_23839001D;SPAN=22167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:88 GQ:45.5 PL:[45.5, 0.0, 167.6] SR:0 DR:21 LR:-45.48 LO:49.44);ALT=T]chr7:23837989];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	24038165	+	chr7	24040071	+	.	49	35	3210279_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATAT;MAPQ=60;MATEID=3210279_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_24034501_24059501_97C;SPAN=1906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:66 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:35 DR:49 LR:-211.3 LO:211.3);ALT=T[chr7:24040071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
