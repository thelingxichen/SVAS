chr8	29962621	+	chr8	28072387	+	.	0	8	5431274_1	16.0	.	EVDNC=ASSMB;HOMSEQ=GAA;MAPQ=60;MATEID=5431274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_29939001_29964001_105C;SPAN=1890234;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:8 DR:0 LR:-16.11 LO:18.33);ALT=]chr8:29962621]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	30604000	+	chr8	30605600	+	.	24	0	5432885_1	69.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5432885_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:30604000(+)-8:30605600(-)__8_30600501_30625501D;SPAN=1600;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:24 DP:19 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=T[chr8:30605600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
