chr1	63944505	+	chr1	63988800	+	ATTTGATAGTCCATTTCTGTGCTTTTGCTCTTCAGAACTTGTGGGAGAAGCAAATAGACTCATTTGACAAGTTCCAGTTGTTGGAGAATAAGTTATAACACTTTTCTTCCTTGTGATTTTTGAAGGATCAAATGAATTTTCTTCTAACAGACCATCCAACTTCAGTGATCTTTTAACA	4	12	180092_1	32.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATTTGATAGTCCATTTCTGTGCTTTTGCTCTTCAGAACTTGTGGGAGAAGCAAATAGACTCATTTGACAAGTTCCAGTTGTTGGAGAATAAGTTATAACACTTTTCTTCCTTGTGATTTTTGAAGGATCAAATGAATTTTCTTCTAACAGACCATCCAACTTCAGTGATCTTTTAACA;MAPQ=60;MATEID=180092_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_63969501_63994501_27C;SPAN=44295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:40 GQ:32 PL:[32.0, 0.0, 65.0] SR:12 DR:4 LR:-32.08 LO:32.69);ALT=C[chr1:63988800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	63955932	+	chr1	63988797	+	.	22	0	180094_1	61.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=180094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:63955932(+)-1:63988797(-)__1_63969501_63994501D;SPAN=32865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:40 GQ:35.3 PL:[61.7, 0.0, 35.3] SR:0 DR:22 LR:-62.17 LO:62.17);ALT=G[chr1:63988797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	64839515	-	chr1	64854716	+	.	23	0	182587_1	66.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=182587_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:64839515(-)-1:64854716(-)__1_64827001_64852001D;SPAN=15201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:7 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:23 LR:-66.02 LO:66.02);ALT=[chr1:64854716[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	65339208	+	chr1	65348958	+	CATCCGGTAGTGGAGCCGGAGGGACATCTTGTCATCAACGGTGATGGTGCGATTTGGAGCATACCAGAGCTTGGTGTTCTCGTCATACAGGGCAAAGAGGTTGTGACAAAGAGGAGAGAT	3	21	183429_1	60.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=CATCCGGTAGTGGAGCCGGAGGGACATCTTGTCATCAACGGTGATGGTGCGATTTGGAGCATACCAGAGCTTGGTGTTCTCGTCATACAGGGCAAAGAGGTTGTGACAAAGAGGAGAGAT;MAPQ=60;MATEID=183429_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_65341501_65366501_68C;SPAN=9750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:57 GQ:60.5 PL:[60.5, 0.0, 77.0] SR:21 DR:3 LR:-60.48 LO:60.6);ALT=T[chr1:65348958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65344831	+	chr1	65348958	+	.	0	11	183439_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AC;MAPQ=60;MATEID=183439_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_65341501_65366501_68C;SPAN=4127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:11 DR:0 LR:-8.677 LO:21.71);ALT=C[chr1:65348958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65349161	+	chr1	65432016	+	CATTTATTCAGCTGTCCAGTGTTCTCCAAGAAGCAAACTGGATTTTCTTCTCTACTTTCCAAAGCTACTTCAGAGAAGCG	0	39	183698_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATTTATTCAGCTGTCCAGTGTTCTCCAAGAAGCAAACTGGATTTTCTTCTCTACTTTCCAAAGCTACTTCAGAGAAGCG;MAPQ=60;MATEID=183698_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_65415001_65440001_64C;SPAN=82855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:17 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:39 DR:0 LR:-115.5 LO:115.5);ALT=G[chr1:65432016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65352069	+	chr1	65432120	+	.	15	0	183701_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=183701_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:65352069(+)-1:65432120(-)__1_65415001_65440001D;SPAN=80051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:19 GQ:1.4 PL:[44.3, 0.0, 1.4] SR:0 DR:15 LR:-46.75 LO:46.75);ALT=C[chr1:65432120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65886423	+	chr1	65890984	+	.	6	3	184985_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=184985_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_65880501_65905501_61C;SPAN=4561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:97 GQ:3 PL:[0.0, 3.0, 240.9] SR:3 DR:6 LR:3.173 LO:12.54);ALT=G[chr1:65890984[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65886476	+	chr1	65895543	+	.	16	0	184988_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=184988_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:65886476(+)-1:65895543(-)__1_65880501_65905501D;SPAN=9067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:98 GQ:26.3 PL:[26.3, 0.0, 211.1] SR:0 DR:16 LR:-26.27 LO:34.69);ALT=T[chr1:65895543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65891061	+	chr1	65897485	+	.	6	3	185002_1	8.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=185002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_65880501_65905501_267C;SPAN=6424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:3 DR:6 LR:-8.035 LO:17.94);ALT=G[chr1:65897485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65891061	+	chr1	65893464	+	.	3	6	185000_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=185000_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_65880501_65905501_187C;SPAN=2403;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:6 DR:3 LR:-11.02 LO:18.56);ALT=G[chr1:65893464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	65891061	+	chr1	65895544	+	.	5	3	185001_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=185001_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_65880501_65905501_315C;SPAN=4483;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:3 DR:5 LR:0.1925 LO:12.92);ALT=G[chr1:65895544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	66024188	+	chr1	66030268	+	.	61	37	185480_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTTTCTTAATGTTTT;MAPQ=60;MATEID=185480_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_66003001_66028001_222C;SPAN=6080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:16 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:37 DR:61 LR:-227.8 LO:227.8);ALT=T[chr1:66030268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	66654829	+	chr1	66668990	+	.	8	0	186632_1	20.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=186632_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:66654829(+)-1:66668990(-)__1_66664501_66689501D;SPAN=14161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:0 DR:8 LR:-19.91 LO:20.23);ALT=A[chr1:66668990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	67390778	+	chr1	67391825	+	.	6	3	188049_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=188049_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_67375001_67400001_129C;SPAN=1047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:91 GQ:4.5 PL:[0.0, 4.5, 227.7] SR:3 DR:6 LR:4.848 LO:10.5);ALT=T[chr1:67391825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	67411979	+	chr1	67423741	+	.	4	9	188167_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=188167_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_1_67399501_67424501_155C;SPAN=11762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:78 GQ:15.2 PL:[15.2, 0.0, 173.6] SR:9 DR:4 LR:-15.18 LO:23.09);ALT=G[chr1:67423741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	68366032	-	chr1	68367217	+	.	8	0	190570_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=190570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:68366032(-)-1:68367217(-)__1_68355001_68380001D;SPAN=1185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=[chr1:68367217[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	68472903	+	chr18	13691676	-	.	9	0	6548738_1	24.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6548738_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:68472903(+)-18:13691676(+)__18_13671001_13696001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:20 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.29 LO:24.29);ALT=A]chr18:13691676];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr13	27050095	+	chr13	27052214	+	.	84	0	5429335_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5429335_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:27050095(+)-13:27052214(-)__13_27048001_27073001D;SPAN=2119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:18 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=G[chr13:27052214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	27999075	+	chr13	28001227	+	.	29	101	5431779_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5431779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_27979001_28004001_97C;SPAN=2152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:113 DP:145 GQ:17 PL:[333.8, 0.0, 17.0] SR:101 DR:29 LR:-350.7 LO:350.7);ALT=G[chr13:28001227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28001329	+	chr13	28004007	+	.	3	30	5432137_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5432137_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28003501_28028501_163C;SPAN=2678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:39 GQ:0.6 PL:[95.7, 0.6, 0.0] SR:30 DR:3 LR:-101.1 LO:101.1);ALT=T[chr13:28004007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28001330	+	chr13	28003309	+	.	3	12	5431787_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5431787_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_27979001_28004001_360C;SPAN=1979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:98 GQ:23 PL:[23.0, 0.0, 214.4] SR:12 DR:3 LR:-22.96 LO:32.06);ALT=G[chr13:28003309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28004103	+	chr13	28008940	+	TGCAGTTTTGAAGACTGTAAGAAGACCTTTAAGAAACATCAGCAGCTGAAAATCCATCAGTGCCAGCATACCAATGAACCTCTATTCAAGTGTACCCAGGAAGGATGTGGGAAACACTTTGCATCACCCAGCAAGCTGAAACGACATGCCAAGGCCCACGAGGGCTATGTATGTCAAAAAGGATGTTCCTTTGTGGCAAAAACATGGACGGAACTTCTGAAACATGTGAGAGAAACCCATAA	0	42	5432143_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGCAGTTTTGAAGACTGTAAGAAGACCTTTAAGAAACATCAGCAGCTGAAAATCCATCAGTGCCAGCATACCAATGAACCTCTATTCAAGTGTACCCAGGAAGGATGTGGGAAACACTTTGCATCACCCAGCAAGCTGAAACGACATGCCAAGGCCCACGAGGGCTATGTATGTCAAAAAGGATGTTCCTTTGTGGCAAAAACATGGACGGAACTTCTGAAACATGTGAGAGAAACCCATAA;MAPQ=60;MATEID=5432143_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_13_28003501_28028501_220C;SPAN=4837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:91 GQ:99 PL:[114.2, 0.0, 104.3] SR:42 DR:0 LR:-114.0 LO:114.0);ALT=A[chr13:28008940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28004760	+	chr13	28006868	+	.	2	15	5432146_1	24.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=5432146_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_13_28003501_28028501_220C;SPAN=2108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:94 GQ:24.2 PL:[24.2, 0.0, 202.4] SR:15 DR:2 LR:-24.05 LO:32.36);ALT=T[chr13:28006868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28004793	+	chr13	28008939	+	.	10	0	5432147_1	6.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5432147_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28004793(+)-13:28008939(-)__13_28003501_28028501D;SPAN=4146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:98 GQ:6.5 PL:[6.5, 0.0, 230.9] SR:0 DR:10 LR:-6.459 LO:19.48);ALT=C[chr13:28008939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28004811	+	chr13	28008273	+	.	19	0	5432148_1	41.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5432148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28004811(+)-13:28008273(-)__13_28003501_28028501D;SPAN=3462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:78 GQ:41.6 PL:[41.6, 0.0, 147.2] SR:0 DR:19 LR:-41.59 LO:44.92);ALT=G[chr13:28008273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28006942	+	chr13	28008275	+	.	2	7	5432156_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=5432156_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=TATGTATG;SCTG=c_13_28003501_28028501_220C;SPAN=1333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:97 GQ:7.8 PL:[0.0, 7.8, 137.6] SR:7 DR:2 LR:8.28 LO:5.709);ALT=G[chr13:28008275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28006994	+	chr13	28008938	+	.	9	0	5432157_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5432157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28006994(+)-13:28008938(-)__13_28003501_28028501D;SPAN=1944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:109 GQ:0.2 PL:[0.2, 0.0, 264.2] SR:0 DR:9 LR:-0.1782 LO:16.67);ALT=C[chr13:28008938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28011411	+	chr13	28014125	+	.	2	5	5432184_1	0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5432184_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28003501_28028501_298C;SPAN=2714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:86 GQ:3.3 PL:[0.0, 3.3, 214.5] SR:5 DR:2 LR:3.494 LO:10.65);ALT=C[chr13:28014125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28014634	+	chr13	28024645	+	.	18	0	5432198_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5432198_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28014634(+)-13:28024645(-)__13_28003501_28028501D;SPAN=10011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:94 GQ:34.1 PL:[34.1, 0.0, 192.5] SR:0 DR:18 LR:-33.95 LO:40.41);ALT=C[chr13:28024645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28015382	+	chr13	28019225	+	.	2	6	5432203_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=5432203_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28003501_28028501_292C;SPAN=3843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:6 DR:2 LR:-2.025 LO:15.08);ALT=T[chr13:28019225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28015414	+	chr13	28024644	+	.	9	0	5432204_1	4.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5432204_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28015414(+)-13:28024644(-)__13_28003501_28028501D;SPAN=9230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:0 DR:9 LR:-4.242 LO:17.27);ALT=A[chr13:28024644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28196147	+	chr13	28222514	+	.	11	12	5432326_1	49.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=5432326_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_13_28175001_28200001_152C;SPAN=26367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:48 GQ:49.7 PL:[49.7, 0.0, 66.2] SR:12 DR:11 LR:-49.72 LO:49.85);ALT=G[chr13:28222514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28196147	+	chr13	28239822	+	AAAGCAATAGAAGAACTGCTTAAGGAGGCAAAACGTGGGAAAACTAGAGCTGAAACAATGGGACCCATGGGTT	14	41	5432327_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AAAGCAATAGAAGAACTGCTTAAGGAGGCAAAACGTGGGAAAACTAGAGCTGAAACAATGGGACCCATGGGTT;MAPQ=60;MATEID=5432327_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_28175001_28200001_152C;SPAN=43675;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:41 DR:14 LR:-141.9 LO:141.9);ALT=G[chr13:28239822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28222591	+	chr13	28239822	+	.	5	32	5432489_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5432489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28224001_28249001_51C;SPAN=17231;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:59 GQ:43.4 PL:[99.5, 0.0, 43.4] SR:32 DR:5 LR:-100.7 LO:100.7);ALT=G[chr13:28239822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28528709	+	chr13	28508271	+	TAGAGATA	43	20	5433347_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TAGAGATA;MAPQ=60;MATEID=5433347_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28493501_28518501_266C;SPAN=20438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:44 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:20 DR:43 LR:-148.5 LO:148.5);ALT=]chr13:28528709]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	28578312	+	chr13	28588589	+	.	9	4	5433507_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5433507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28567001_28592001_84C;SPAN=10277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:101 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:4 DR:9 LR:-12.25 LO:24.22);ALT=C[chr13:28588589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28592727	+	chr13	28597487	+	.	0	9	5433673_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5433673_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28591501_28616501_212C;SPAN=4760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:9 DR:0 LR:-5.868 LO:17.54);ALT=C[chr13:28597487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28602427	+	chr13	28608024	+	.	0	8	5433715_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5433715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28591501_28616501_393C;SPAN=5597;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-1.754 LO:15.04);ALT=T[chr13:28608024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28636207	+	chr13	28644625	+	.	2	12	5433854_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACC;MAPQ=60;MATEID=5433854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28616001_28641001_173C;SPAN=8418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:44 GQ:34.4 PL:[34.4, 0.0, 70.7] SR:12 DR:2 LR:-34.29 LO:35.04);ALT=C[chr13:28644625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28636250	+	chr13	28674604	+	.	29	0	5433855_1	84.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5433855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28636250(+)-13:28674604(-)__13_28616001_28641001D;SPAN=38354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:40 GQ:12.2 PL:[84.8, 0.0, 12.2] SR:0 DR:29 LR:-88.02 LO:88.02);ALT=T[chr13:28674604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28644750	+	chr13	28674605	+	.	24	9	5434460_1	53.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5434460_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=CAACAA;SCTG=c_13_28665001_28690001_168C;SPAN=29855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:45 GQ:27 PL:[53.0, 0.0, 27.0] SR:9 DR:24 LR:-53.34 LO:53.34);ALT=C[chr13:28674605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28650935	+	chr13	28674635	+	.	34	0	5434461_1	96.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5434461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:28650935(+)-13:28674635(-)__13_28665001_28690001D;SPAN=23700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:58 GQ:43.7 PL:[96.5, 0.0, 43.7] SR:0 DR:34 LR:-97.57 LO:97.57);ALT=G[chr13:28674635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	28712565	+	chr13	28748409	+	.	2	2	5434221_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5434221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_28738501_28763501_343C;SPAN=35844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:44 GQ:1.4 PL:[1.4, 0.0, 103.7] SR:2 DR:2 LR:-1.283 LO:7.582);ALT=A[chr13:28748409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29233324	+	chr13	29236546	+	.	5	11	5435637_1	7.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5435637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_29228501_29253501_347C;SPAN=3222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:155 GQ:7.6 PL:[7.6, 0.0, 367.4] SR:11 DR:5 LR:-7.522 LO:28.86);ALT=G[chr13:29236546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29233366	+	chr13	29238644	+	.	48	0	5435638_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5435638_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:29233366(+)-13:29238644(-)__13_29228501_29253501D;SPAN=5278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:114 GQ:99 PL:[127.7, 0.0, 147.5] SR:0 DR:48 LR:-127.6 LO:127.7);ALT=G[chr13:29238644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29233377	+	chr13	29242609	+	.	52	0	5435640_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5435640_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:29233377(+)-13:29242609(-)__13_29228501_29253501D;SPAN=9232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:132 GQ:99 PL:[136.1, 0.0, 182.3] SR:0 DR:52 LR:-135.9 LO:136.3);ALT=C[chr13:29242609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29233377	+	chr13	29246473	+	.	11	0	5435641_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5435641_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:29233377(+)-13:29246473(-)__13_29228501_29253501D;SPAN=13096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:122 GQ:3.5 PL:[3.5, 0.0, 290.6] SR:0 DR:11 LR:-3.258 LO:20.81);ALT=C[chr13:29246473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29236629	+	chr13	29246473	+	.	9	0	5435652_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5435652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:29236629(+)-13:29246473(-)__13_29228501_29253501D;SPAN=9844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:123 GQ:3.3 PL:[0.0, 3.3, 303.6] SR:0 DR:9 LR:3.615 LO:16.17);ALT=A[chr13:29246473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29236644	+	chr13	29238645	+	.	14	79	5435653_1	99.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5435653_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_13_29228501_29253501_364C;SPAN=2001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:104 GQ:1.5 PL:[254.1, 1.5, 0.0] SR:79 DR:14 LR:-268.1 LO:268.1);ALT=G[chr13:29238645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29236644	+	chr13	29242610	+	TTTTTCTTGTGTGAAAAATGAACTTTTGCCTAGTCATCCCCTTGAATTATCAGAAAAAAAT	28	155	5435654_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTTTCTTGTGTGAAAAATGAACTTTTGCCTAGTCATCCCCTTGAATTATCAGAAAAAAAT;MAPQ=60;MATEID=5435654_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_29228501_29253501_364C;SPAN=5966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:171 DP:124 GQ:46 PL:[505.0, 46.0, 0.0] SR:155 DR:28 LR:-505.0 LO:505.0);ALT=G[chr13:29242610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29242713	+	chr13	29246474	+	.	2	69	5435668_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5435668_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_29228501_29253501_265C;SPAN=3761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:124 GQ:98.6 PL:[200.9, 0.0, 98.6] SR:69 DR:2 LR:-202.6 LO:202.6);ALT=T[chr13:29246474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	29246569	+	chr13	29252171	+	.	0	107	5435684_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5435684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_29228501_29253501_238C;SPAN=5602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:107 DP:136 GQ:12.8 PL:[316.4, 0.0, 12.8] SR:107 DR:0 LR:-333.1 LO:333.1);ALT=G[chr13:29252171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	30215837	+	chr13	30221845	+	.	21	19	5438617_1	95.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GAGAACTACTTTTT;MAPQ=60;MATEID=5438617_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_30208501_30233501_58C;SPAN=6008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:63 GQ:55.7 PL:[95.3, 0.0, 55.7] SR:19 DR:21 LR:-95.66 LO:95.66);ALT=T[chr13:30221845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	31127882	-	chr18	12884124	+	.	14	0	6546250_1	32.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6546250_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:31127882(-)-18:12884124(-)__18_12862501_12887501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:53 GQ:32 PL:[32.0, 0.0, 94.7] SR:0 DR:14 LR:-31.86 LO:33.68);ALT=[chr18:12884124[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr13	31309802	+	chr13	31330078	+	.	12	0	5441992_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5441992_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:31309802(+)-13:31330078(-)__13_31286501_31311501D;SPAN=20276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=G[chr13:31330078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	31309806	+	chr13	31326185	+	.	21	0	5441993_1	57.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5441993_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:31309806(+)-13:31326185(-)__13_31286501_31311501D;SPAN=16379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:44 GQ:47.6 PL:[57.5, 0.0, 47.6] SR:0 DR:21 LR:-57.43 LO:57.43);ALT=C[chr13:31326185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	31309813	+	chr13	31318196	+	.	25	15	5441994_1	87.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5441994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_31286501_31311501_38C;SPAN=8383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:42 GQ:11.9 PL:[87.8, 0.0, 11.9] SR:15 DR:25 LR:-90.67 LO:90.67);ALT=G[chr13:31318196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	31318296	+	chr13	31326189	+	.	2	28	5441816_1	67.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=5441816_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_13_31311001_31336001_125C;SPAN=7893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:106 GQ:67.1 PL:[67.1, 0.0, 189.2] SR:28 DR:2 LR:-67.01 LO:70.29);ALT=A[chr13:31326189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	31318296	+	chr13	31330079	+	CCAGAACTGTGTAGATGCGTACCCCACTTTCCTCGCTGTGCTCTGGTCTGCGGGGCTACTTTGCAGCCA	2	49	5441817_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCAGAACTGTGTAGATGCGTACCCCACTTTCCTCGCTGTGCTCTGGTCTGCGGGGCTACTTTGCAGCCA;MAPQ=60;MATEID=5441817_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_31311001_31336001_125C;SPAN=11783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:103 GQ:99 PL:[137.3, 0.0, 110.9] SR:49 DR:2 LR:-137.3 LO:137.3);ALT=A[chr13:31330079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	11973033	-	chr18	11974170	+	.	8	0	6543868_1	13.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6543868_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:11973033(-)-18:11974170(-)__18_11956001_11981001D;SPAN=1137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=[chr18:11974170[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	11981764	+	chr18	11999050	+	.	0	11	6543565_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6543565_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_11980501_12005501_81C;SPAN=17286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:11 DR:0 LR:-15.72 LO:23.22);ALT=G[chr18:11999050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12308362	+	chr18	12310941	+	.	13	0	6544398_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6544398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:12308362(+)-18:12310941(-)__18_12299001_12324001D;SPAN=2579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:51 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:0 DR:13 LR:-29.1 LO:31.04);ALT=G[chr18:12310941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12308794	+	chr18	12310942	+	.	0	13	6544400_1	22.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6544400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_12299001_12324001_202C;SPAN=2148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:75 GQ:22.7 PL:[22.7, 0.0, 158.0] SR:13 DR:0 LR:-22.59 LO:28.56);ALT=T[chr18:12310942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12703163	+	chr18	12706548	+	.	79	19	6545731_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6545731_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_12691001_12716001_71C;SPAN=3385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:85 GQ:24 PL:[264.0, 24.0, 0.0] SR:19 DR:79 LR:-264.1 LO:264.1);ALT=G[chr18:12706548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12703190	+	chr18	12712698	+	.	10	0	6545732_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6545732_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:12703190(+)-18:12712698(-)__18_12691001_12716001D;SPAN=9508;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:63 GQ:16.1 PL:[16.1, 0.0, 134.9] SR:0 DR:10 LR:-15.94 LO:21.55);ALT=G[chr18:12712698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	12718634	+	chr18	12720506	+	.	6	7	6545552_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAG;MAPQ=60;MATEID=6545552_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_12715501_12740501_144C;SPAN=1872;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:65 GQ:22.1 PL:[22.1, 0.0, 134.3] SR:7 DR:6 LR:-22.0 LO:26.73);ALT=G[chr18:12720506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	13682106	+	chr18	13726328	+	.	0	7	6548788_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6548788_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_13671001_13696001_220C;SPAN=44222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:36 GQ:13.4 PL:[13.4, 0.0, 72.8] SR:7 DR:0 LR:-13.35 LO:15.77);ALT=T[chr18:13726328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	13726768	+	chr18	13731472	+	.	27	0	6548453_1	67.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6548453_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:13726768(+)-18:13731472(-)__18_13720001_13745001D;SPAN=4704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:81 GQ:67.4 PL:[67.4, 0.0, 126.8] SR:0 DR:27 LR:-67.18 LO:68.26);ALT=G[chr18:13731472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
