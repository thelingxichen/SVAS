chr12	33689912	-	chr12	33692963	+	.	9	0	7539910_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7539910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:33689912(-)-12:33692963(-)__12_33687501_33712501D;SPAN=3051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:210 GQ:27.1 PL:[0.0, 27.1, 564.4] SR:0 DR:9 LR:27.19 LO:14.03);ALT=[chr12:33692963[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	34617603	+	chr12	34634570	-	.	9	0	7545421_1	5.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7545421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:34617603(+)-12:34634570(+)__12_34594001_34619001D;SPAN=16967;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:0 DR:9 LR:-5.868 LO:17.54);ALT=T]chr12:34634570];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	34618009	-	chr12	34634409	+	.	14	0	7545422_1	28.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=7545422_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:34618009(-)-12:34634409(-)__12_34594001_34619001D;SPAN=16400;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:0 DR:14 LR:-28.06 LO:32.03);ALT=[chr12:34634409[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
