chr13	72843037	+	chr13	72846925	+	AAATTGCAG	0	94	8147024_1	99.0	.	EVDNC=ASSMB;INSERTION=AAATTGCAG;MAPQ=60;MATEID=8147024_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_13_72838501_72863501_44C;SPAN=3888;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:44 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:94 DR:0 LR:-277.3 LO:277.3);ALT=T[chr13:72846925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
