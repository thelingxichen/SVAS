chr4	152680075	+	chr4	152681959	+	.	0	8	2274722_1	2.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2274722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_152659501_152684501_168C;SPAN=1884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:8 DR:0 LR:-2.567 LO:15.16);ALT=C[chr4:152681959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
