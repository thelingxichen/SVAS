chr5	19375269	+	chr5	19376397	+	TGG	48	34	2428201_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TGG;MAPQ=60;MATEID=2428201_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_19355001_19380001_136C;SPAN=1128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:17 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:34 DR:48 LR:-188.1 LO:188.1);ALT=A[chr5:19376397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
