chr10	58894812	+	chr10	58937152	+	.	85	82	6288258_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;MAPQ=60;MATEID=6288258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_58922501_58947501_314C;SPAN=42340;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:133 DP:44 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:82 DR:85 LR:-392.8 LO:392.8);ALT=A[chr10:58937152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
