chr7	113416176	+	chr7	113422208	+	.	100	65	3532589_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CATAATGGCATTTTT;MAPQ=60;MATEID=3532589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_113410501_113435501_100C;SPAN=6032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:142 DP:74 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:65 DR:100 LR:-419.2 LO:419.2);ALT=T[chr7:113422208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
