chr9	88307775	+	chr9	88356718	+	.	12	0	4312521_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4312521_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:88307775(+)-9:88356718(-)__9_88298001_88323001D;SPAN=48943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=A[chr9:88356718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	89201789	+	chr18	40322295	-	.	17	0	6602204_1	45.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6602204_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:89201789(+)-18:40322295(+)__18_40302501_40327501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:0 DR:17 LR:-45.01 LO:45.06);ALT=A]chr18:40322295];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr18	38259893	+	chr18	38266750	+	.	22	19	6597774_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6597774_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_38244501_38269501_156C;SPAN=6857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:61 GQ:43.1 PL:[102.5, 0.0, 43.1] SR:19 DR:22 LR:-103.5 LO:103.5);ALT=T[chr18:38266750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	38864779	+	chr18	38868344	+	TAAAACTCTTAAG	51	26	6599232_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TAAAACTCTTAAG;MAPQ=60;MATEID=6599232_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_38857001_38882001_230C;SPAN=3565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:18 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:26 DR:51 LR:-184.8 LO:184.8);ALT=T[chr18:38868344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	39535371	+	chr18	39537534	+	.	10	0	6600492_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6600492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:39535371(+)-18:39537534(-)__18_39518501_39543501D;SPAN=2163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:0 DR:10 LR:-10.79 LO:20.31);ALT=A[chr18:39537534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	39537723	+	chr18	39542454	+	.	3	6	6600498_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6600498_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_39518501_39543501_157C;SPAN=4731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:68 GQ:4.7 PL:[4.7, 0.0, 159.8] SR:6 DR:3 LR:-4.684 LO:13.67);ALT=A[chr18:39542454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
