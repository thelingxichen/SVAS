chr13	54670445	+	chr13	54678812	+	TATGGTAAAG	0	41	5505506_1	99.0	.	EVDNC=ASSMB;INSERTION=TATGGTAAAG;MAPQ=60;MATEID=5505506_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_54659501_54684501_196C;SPAN=8367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:72 GQ:56.6 PL:[116.0, 0.0, 56.6] SR:41 DR:0 LR:-116.8 LO:116.8);ALT=G[chr13:54678812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
