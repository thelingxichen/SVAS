chr5	178109066	+	chr5	178113412	+	.	32	39	3963581_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GAGAT;MAPQ=60;MATEID=3963581_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_178090501_178115501_358C;SPAN=4346;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:65 DP:80 GQ:1.4 PL:[192.8, 0.0, 1.4] SR:39 DR:32 LR:-204.6 LO:204.6);ALT=T[chr5:178113412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
