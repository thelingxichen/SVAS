chrX	130813253	+	chrX	130974276	-	.	12	30	7526951_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TAGACACACAC;MAPQ=60;MATEID=7526951_2;MATENM=2;NM=5;NUMPARTS=2;SCTG=c_23_130952501_130977501_257C;SPAN=161023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:13 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:30 DR:12 LR:-115.5 LO:115.5);ALT=C]chrX:130974276];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	131205246	+	chrX	131206296	+	.	2	3	7527152_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7527152_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_131197501_131222501_134C;SPAN=1050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:50 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:3 DR:2 LR:0.3422 LO:7.35);ALT=G[chrX:131206296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
