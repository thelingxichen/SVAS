chrY	15019505	+	chrY	15021271	+	.	0	7	7564911_1	20.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7564911_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_24_15018501_15043501_3C;SPAN=1766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:9 GQ:0.8 PL:[20.6, 0.0, 0.8] SR:7 DR:0 LR:-21.71 LO:21.71);ALT=A[chrY:15021271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
