chr13	107196509	+	chr13	107209395	+	.	11	10	5636320_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=5636320_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_13_107187501_107212501_59C;SPAN=12886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:72 GQ:36.8 PL:[36.8, 0.0, 135.8] SR:10 DR:11 LR:-36.61 LO:39.93);ALT=C[chr13:107209395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	107212005	+	chr13	107219921	+	.	14	25	5636446_1	72.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=5636446_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_107212001_107237001_194C;SPAN=7916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:97 GQ:72.8 PL:[72.8, 0.0, 161.9] SR:25 DR:14 LR:-72.75 LO:74.64);ALT=A[chr13:107219921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
