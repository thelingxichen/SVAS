chr6	52242022	+	chr6	52075273	+	.	8	5	4208106_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4208106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_52234001_52259001_68C;SPAN=166749;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:5 DR:8 LR:-16.75 LO:21.78);ALT=]chr6:52242022]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	52651110	+	chr6	52652674	+	TAGATTAAGTAAAATGACATCATGACTATTATTTCCCCTCATGAC	29	111	4210320_1	99.0	.	DISC_MAPQ=44;EVDNC=TSI_L;INSERTION=TAGATTAAGTAAAATGACATCATGACTATTATTTCCCCTCATGAC;MAPQ=60;MATEID=4210320_2;MATENM=8;NM=8;NUMPARTS=3;SCTG=c_6_52650501_52675501_179C;SPAN=1564;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:126 DP:176 GQ:58 PL:[368.3, 0.0, 58.0] SR:111 DR:29 LR:-381.1 LO:381.1);ALT=T[chr6:52652674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
