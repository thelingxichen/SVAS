chr1	38432782	+	chr6	28863899	-	.	57	59	193709_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;MAPQ=60;MATEID=193709_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_38416001_38441001_385C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:45 GQ:27 PL:[297.0, 27.0, 0.0] SR:59 DR:57 LR:-297.1 LO:297.1);ALT=G]chr6:28863899];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	38095059	-	chr6	29863616	+	.	8	73	1953661_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=GGGAGGTGGGGGGCAGCCCC;MAPQ=41;MATEID=1953661_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_38073001_38098001_71C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:88 GQ:13.8 PL:[240.9, 13.8, 0.0] SR:73 DR:8 LR:-245.0 LO:245.0);ALT=[chr6:29863616[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	29685488	+	chr6	29688081	+	.	126	39	4105487_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAGAAAGACCCAAGCCT;MAPQ=60;MATEID=4105487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_29669501_29694501_170C;SPAN=2593;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:140 DP:837 GQ:99 PL:[235.6, 0.0, 1797.0] SR:39 DR:126 LR:-235.4 LO:305.2);ALT=T[chr6:29688081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29766211	+	chr6	29922619	+	.	60	0	4106421_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4106421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29766211(+)-6:29922619(-)__6_29914501_29939501D;SPAN=156408;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:12 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=T[chr6:29922619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29876631	+	chr6	29832275	+	.	9	0	4106185_1	17.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=4106185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29832275(-)-6:29876631(+)__6_29816501_29841501D;SPAN=44356;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=]chr6:29876631]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	29910758	+	chr6	29855942	+	.	22	92	4106031_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CACAGACTGACCGAG;MAPQ=37;MATEID=4106031_2;MATENM=4;NM=2;NUMPARTS=2;SCTG=c_6_29890001_29915001_52C;SPAN=54816;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:101 DP:15 GQ:27 PL:[297.0, 27.0, 0.0] SR:92 DR:22 LR:-297.1 LO:297.1);ALT=]chr6:29910758]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	29914600	+	chr6	29899648	+	.	16	0	4106040_1	31.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=4106040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29899648(-)-6:29914600(+)__6_29890001_29915001D;SPAN=14952;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:78 GQ:31.7 PL:[31.7, 0.0, 157.1] SR:0 DR:16 LR:-31.68 LO:36.46);ALT=]chr6:29914600]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	29899785	+	chr6	29914896	+	.	14	0	4106041_1	26.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=4106041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29899785(+)-6:29914896(-)__6_29890001_29915001D;SPAN=15111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:73 GQ:26.6 PL:[26.6, 0.0, 148.7] SR:0 DR:14 LR:-26.44 LO:31.44);ALT=T[chr6:29914896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30486061	+	chr10	116796712	+	.	0	9	6541559_1	7.0	.	EVDNC=ASSMB;HOMSEQ=TGTGTCTAGCTAAAGGATTGTAAA;MAPQ=60;MATEID=6541559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_116791501_116816501_303C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:9 DR:0 LR:-7.222 LO:17.79);ALT=A[chr10:116796712[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	30718984	+	chr6	30720392	+	.	67	39	4109661_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4109661_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30698501_30723501_275C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:67 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:39 DR:67 LR:-244.3 LO:244.3);ALT=T[chr6:30720392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31210339	+	chr6	31287118	+	.	9	0	4118269_1	12.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=4118269_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31210339(+)-6:31287118(-)__6_31286501_31311501D;SPAN=76779;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:0 DR:9 LR:-12.1 LO:18.81);ALT=T[chr6:31287118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31211630	+	chr6	31213117	+	.	168	84	4112585_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AATACCCACCACCC;MAPQ=60;MATEID=4112585_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_6_31188501_31213501_74C;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:212 DP:83 GQ:57.1 PL:[627.1, 57.1, 0.0] SR:84 DR:168 LR:-627.2 LO:627.2);ALT=C[chr6:31213117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31235303	-	chr6	31236724	+	.	9	0	4112816_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=4112816_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31235303(-)-6:31236724(-)__6_31213001_31238001D;SPAN=1421;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:128 GQ:4.8 PL:[0.0, 4.8, 320.1] SR:0 DR:9 LR:4.969 LO:16.01);ALT=[chr6:31236724[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	31296275	+	chr6	31304750	+	.	32	0	4118341_1	77.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=4118341_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31296275(+)-6:31304750(-)__6_31286501_31311501D;SPAN=8475;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:103 GQ:77.9 PL:[77.9, 0.0, 170.3] SR:0 DR:32 LR:-77.73 LO:79.7);ALT=A[chr6:31304750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31776260	+	chr6	31544164	+	.	60	16	4115946_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=4115946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31752001_31777001_79C;SPAN=232096;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:50 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:16 DR:60 LR:-194.7 LO:194.7);ALT=]chr6:31776260]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	117006342	+	chrX	128670974	-	.	29	49	11380376_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=11380376_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_128649501_128674501_167C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:37 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:49 DR:29 LR:-208.0 LO:208.0);ALT=T]chrX:128670974];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	117847133	+	chr10	118538221	+	.	72	47	6545199_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6545199_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_117845001_117870001_2C;SPAN=691088;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:40 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:47 DR:72 LR:-277.3 LO:277.3);ALT=T[chr10:118538221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
