chr13	101205427	+	chr13	101208764	+	.	78	61	8276761_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATGG;MAPQ=60;MATEID=8276761_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_101185001_101210001_219C;SPAN=3337;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:111 DP:156 GQ:53.6 PL:[324.2, 0.0, 53.6] SR:61 DR:78 LR:-335.1 LO:335.1);ALT=G[chr13:101208764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	101894146	+	chr13	101896425	+	.	75	21	8280974_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CAT;MAPQ=60;MATEID=8280974_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_101871001_101896001_8C;SPAN=2279;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:76 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:21 DR:75 LR:-270.7 LO:270.7);ALT=T[chr13:101896425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
