chr5	76808191	-	chr12	51017186	+	.	4	45	3549733_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACACACACACACACACACACACACACACACACACAC;MAPQ=60;MATEID=3549733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_76807501_76832501_306C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:52 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:45 DR:4 LR:-151.8 LO:151.8);ALT=[chr12:51017186[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	50973716	+	chr12	50975506	+	.	59	38	7603424_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCCACT;MAPQ=60;MATEID=7603424_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_12_50960001_50985001_118C;SPAN=1790;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:73 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:38 DR:59 LR:-221.2 LO:221.2);ALT=T[chr12:50975506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
