chr14	91963666	-	chr14	91965728	+	.	8	0	8678161_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=8678161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:91963666(-)-14:91965728(-)__14_91948501_91973501D;SPAN=2062;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:139 GQ:11.1 PL:[0.0, 11.1, 359.7] SR:0 DR:8 LR:11.25 LO:13.52);ALT=[chr14:91965728[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
