chr7	117824309	+	chr7	117825708	+	.	6	12	3546258_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3546258_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_117820501_117845501_239C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:116 GQ:11.6 PL:[11.6, 0.0, 269.0] SR:12 DR:6 LR:-11.49 LO:25.89);ALT=G[chr7:117825708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	117824309	+	chr7	117831966	+	AACTGTTGCCGTTATTACATCAGATGGGAGAATGATTGTGGGAACACTGAAAGGTTTTGACCAGACCATTAATTTGATTTTGGATGAAAGCCATGAACGAGTATTCAGCTCTTCACAGGGGGTAGAACAAGTGGTACTAGGATTATACATTGTAAGAGGTGACAACGT	10	48	3546259_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AACTGTTGCCGTTATTACATCAGATGGGAGAATGATTGTGGGAACACTGAAAGGTTTTGACCAGACCATTAATTTGATTTTGGATGAAAGCCATGAACGAGTATTCAGCTCTTCACAGGGGGTAGAACAAGTGGTACTAGGATTATACATTGTAAGAGGTGACAACGT;MAPQ=60;MATEID=3546259_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_117820501_117845501_239C;SPAN=7657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:123 GQ:99 PL:[131.9, 0.0, 164.9] SR:48 DR:10 LR:-131.7 LO:132.0);ALT=G[chr7:117831966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	117824331	+	chr7	117828330	+	.	48	0	3546260_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3546260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:117824331(+)-7:117828330(-)__7_117820501_117845501D;SPAN=3999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:120 GQ:99 PL:[125.9, 0.0, 165.5] SR:0 DR:48 LR:-125.9 LO:126.2);ALT=G[chr7:117828330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
