chr2	150436162	+	chr2	150444178	+	ATATATCTGGAGGTGCAGCAGCCACATGAGACTCATCCGAACCTGATGATCCTGCAGTCGAAAAGGCTTTGGGATTGACAACCCTTTTAACTAAAGAGCAAAATCCTGGGAGATAGGAAACCAGTCTGGCTCTGTTACAAAGCACATTGGCCATCTCCGCTGGAGAAGATAGTTCGCAAAATAGCTTTCCTTTGGTAAAGTTATTT	13	42	1039516_1	99.0	.	DISC_MAPQ=25;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATATATCTGGAGGTGCAGCAGCCACATGAGACTCATCCGAACCTGATGATCCTGCAGTCGAAAAGGCTTTGGGATTGACAACCCTTTTAACTAAAGAGCAAAATCCTGGGAGATAGGAAACCAGTCTGGCTCTGTTACAAAGCACATTGGCCATCTCCGCTGGAGAAGATAGTTCGCAAAATAGCTTTCCTTTGGTAAAGTTATTT;MAPQ=60;MATEID=1039516_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_150430001_150455001_29C;SPAN=8016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:103 GQ:99 PL:[117.5, 0.0, 130.7] SR:42 DR:13 LR:-117.3 LO:117.4);ALT=C[chr2:150444178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	150438828	+	chr2	150444177	+	.	77	0	1039533_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=1039533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:150438828(+)-2:150444177(-)__2_150430001_150455001D;SPAN=5349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:94 GQ:2.1 PL:[231.0, 2.1, 0.0] SR:0 DR:77 LR:-243.1 LO:243.1);ALT=A[chr2:150444177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
