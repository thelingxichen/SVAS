chr12	47979593	-	chr12	47981822	+	.	9	0	7588840_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=7588840_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:47979593(-)-12:47981822(-)__12_47971001_47996001D;SPAN=2229;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:185 GQ:20.2 PL:[0.0, 20.2, 488.5] SR:0 DR:9 LR:20.41 LO:14.54);ALT=[chr12:47981822[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
