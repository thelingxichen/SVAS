chr3	98410686	+	chr3	98414783	+	.	63	0	2190312_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2190312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:98410686(+)-3:98414783(-)__3_98392001_98417001D;SPAN=4097;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:15 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:0 DR:63 LR:-184.8 LO:184.8);ALT=A[chr3:98414783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	98754923	+	chr8	138827171	-	.	11	0	2191776_1	26.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2191776_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:98754923(+)-8:138827171(+)__3_98735001_98760001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:0 DR:11 LR:-26.29 LO:27.14);ALT=T]chr8:138827171];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	98899063	+	chr3	98902390	+	.	72	63	2191944_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=2191944_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_98882001_98907001_481C;SPAN=3327;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:84 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:63 DR:72 LR:-310.3 LO:310.3);ALT=T[chr3:98902390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	99298388	+	chr3	99299429	-	.	3	1	2193400_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=2193400_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_99274001_99299001_248C;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:1 DR:3 LR:6.844 LO:6.647);ALT=A]chr3:99299429];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	99817368	+	chr3	99536534	+	.	39	35	2195334_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAT;MAPQ=60;MATEID=2195334_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_99813001_99838001_344C;SPAN=280834;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:64 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:35 DR:39 LR:-188.1 LO:188.1);ALT=]chr3:99817368]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	51541549	+	chr5	51543168	-	.	9	0	3419367_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3419367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:51541549(+)-5:51543168(+)__5_51523501_51548501D;SPAN=1619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:113 GQ:0.6 PL:[0.0, 0.6, 273.9] SR:0 DR:9 LR:0.9055 LO:16.52);ALT=A]chr5:51543168];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	52473558	+	chr8	138259033	-	GTATATA	4	27	3422799_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTATATA;MAPQ=60;MATEID=3422799_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_52454501_52479501_360C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:27 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:27 DR:4 LR:-82.52 LO:82.52);ALT=A]chr8:138259033];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	52805997	+	chr5	52716477	+	.	65	63	3424182_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTTG;MAPQ=60;MATEID=3424182_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_52797501_52822501_368C;SPAN=89520;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:73 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:63 DR:65 LR:-313.6 LO:313.6);ALT=]chr5:52805997]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	53122614	-	chr5	53125512	+	TAAT	46	90	3425665_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TAAT;MAPQ=60;MATEID=3425665_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_53116001_53141001_79C;SPAN=2898;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:125 DP:127 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:90 DR:46 LR:-376.3 LO:376.3);ALT=[chr5:53125512[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	53122763	+	chr5	53125485	-	TTCAGTTAG	43	99	3425667_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTCAGTTAG;MAPQ=60;MATEID=3425667_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_53116001_53141001_163C;SPAN=2722;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:130 DP:115 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:99 DR:43 LR:-386.2 LO:386.2);ALT=G]chr5:53125485];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	53142469	+	chr5	53144942	-	.	13	0	3426164_1	12.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=3426164_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:53142469(+)-5:53144942(+)__5_53140501_53165501D;SPAN=2473;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:112 GQ:12.8 PL:[12.8, 0.0, 257.0] SR:0 DR:13 LR:-12.57 LO:26.1);ALT=C]chr5:53144942];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	137945250	-	chr8	137946688	+	.	11	0	5725101_1	7.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5725101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:137945250(-)-8:137946688(-)__8_137935001_137960001D;SPAN=1438;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:0 DR:11 LR:-7.051 LO:21.42);ALT=[chr8:137946688[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	138125855	+	chr8	138127582	+	TTTAATTTCCTC	59	27	5725739_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TTTAATTTCCTC;MAPQ=60;MATEID=5725739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_138106501_138131501_325C;SPAN=1727;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:63 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:27 DR:59 LR:-227.8 LO:227.8);ALT=C[chr8:138127582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
