chr8	67344822	+	chr8	67356599	+	.	10	0	3897634_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3897634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67344822(+)-8:67356599(-)__8_67350501_67375501D;SPAN=11777;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:44 GQ:21.2 PL:[21.2, 0.0, 83.9] SR:0 DR:10 LR:-21.09 LO:23.3);ALT=G[chr8:67356599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67579934	+	chr8	67588976	+	.	9	0	3898447_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3898447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67579934(+)-8:67588976(-)__8_67571001_67596001D;SPAN=9042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:100 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.617 LO:17.02);ALT=A[chr8:67588976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67625106	+	chr8	67705848	+	.	10	0	3898795_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3898795_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67625106(+)-8:67705848(-)__8_67693501_67718501D;SPAN=80742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:44 GQ:21.2 PL:[21.2, 0.0, 83.9] SR:0 DR:10 LR:-21.09 LO:23.3);ALT=G[chr8:67705848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67834405	+	chr8	67837679	+	.	38	0	3899348_1	92.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3899348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67834405(+)-8:67837679(-)__8_67816001_67841001D;SPAN=3274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:120 GQ:92.9 PL:[92.9, 0.0, 198.5] SR:0 DR:38 LR:-92.93 LO:95.02);ALT=T[chr8:67837679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67834677	+	chr8	67837691	+	.	49	0	3899353_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3899353_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67834677(+)-8:67837691(-)__8_67816001_67841001D;SPAN=3014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:114 GQ:99 PL:[131.0, 0.0, 144.2] SR:0 DR:49 LR:-130.9 LO:130.9);ALT=T[chr8:67837691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67834962	+	chr8	67837669	+	.	71	22	3899357_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=3899357_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_67816001_67841001_48C;SPAN=2707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:84 DP:123 GQ:52.7 PL:[244.1, 0.0, 52.7] SR:22 DR:71 LR:-250.7 LO:250.7);ALT=T[chr8:67837669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	67971735	+	chr8	67974095	+	.	14	0	3899832_1	21.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3899832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:67971735(+)-8:67974095(-)__8_67963001_67988001D;SPAN=2360;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:0 DR:14 LR:-21.29 LO:29.89);ALT=A[chr8:67974095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	68578998	-	chr8	68580168	+	.	8	0	3901446_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3901446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:68578998(-)-8:68580168(-)__8_68575501_68600501D;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=[chr8:68580168[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
