chr12	98955403	+	chr12	98959001	+	.	37	46	5305006_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5305006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_98955501_98980501_86C;SPAN=3598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:23 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:46 DR:37 LR:-204.7 LO:204.7);ALT=G[chr12:98959001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98987551	+	chr12	98991631	+	.	10	0	5305197_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5305197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:98987551(+)-12:98991631(-)__12_98980001_99005001D;SPAN=4080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:0 DR:10 LR:-6.73 LO:19.53);ALT=T[chr12:98991631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98987551	+	chr12	98989501	+	.	46	0	5305196_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5305196_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:98987551(+)-12:98989501(-)__12_98980001_99005001D;SPAN=1950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:139 GQ:99 PL:[114.2, 0.0, 223.1] SR:0 DR:46 LR:-114.2 LO:116.1);ALT=T[chr12:98989501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98987913	+	chr12	98992298	+	AGTACAGTTGTGAATTTGGCTCCGCGAAGTATTATGCACTGTGTGGCTTTGGTGGGGTCTTAAGTTGTGGTCTGACACACACTGCTGTGGTTCCCCTGGATTTAGTGAAATGCCGTATGCAGGTGGACCCCCAAAAGTACAAGGGCATATTTAACGGATTCTCAGTTACACTTAAAGAGGATGGTGTTCGTGGTTTGGCTAAAGGATGGGCTCCGACTTTCCTTGGCTACTCCATGCAGGGACTCTGCAAGTTTGGCTTTTATGAAGTCTTTAAAGTCTTGTATAGCAATATGCTTGGAG	0	156	5305202_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AGTACAGTTGTGAATTTGGCTCCGCGAAGTATTATGCACTGTGTGGCTTTGGTGGGGTCTTAAGTTGTGGTCTGACACACACTGCTGTGGTTCCCCTGGATTTAGTGAAATGCCGTATGCAGGTGGACCCCCAAAAGTACAAGGGCATATTTAACGGATTCTCAGTTACACTTAAAGAGGATGGTGTTCGTGGTTTGGCTAAAGGATGGGCTCCGACTTTCCTTGGCTACTCCATGCAGGGACTCTGCAAGTTTGGCTTTTATGAAGTCTTTAAAGTCTTGTATAGCAATATGCTTGGAG;MAPQ=60;MATEID=5305202_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_98980001_99005001_226C;SPAN=4385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:156 DP:120 GQ:42.1 PL:[462.1, 42.1, 0.0] SR:156 DR:0 LR:-462.1 LO:462.1);ALT=G[chr12:98992298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98987913	+	chr12	98989503	+	.	7	146	5305201_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5305201_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_98980001_99005001_226C;SPAN=1590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:174 GQ:27.1 PL:[475.3, 27.1, 0.0] SR:146 DR:7 LR:-483.2 LO:483.2);ALT=G[chr12:98989503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98989628	+	chr12	98991632	+	.	2	45	5305208_1	99.0	.	DISC_MAPQ=42;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=5305208_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_98980001_99005001_226C;SPAN=2004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:83 GQ:70.1 PL:[129.5, 0.0, 70.1] SR:45 DR:2 LR:-130.2 LO:130.2);ALT=T[chr12:98991632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98992507	+	chr12	98993731	+	.	11	0	5305219_1	16.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5305219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:98992507(+)-12:98993731(-)__12_98980001_99005001D;SPAN=1224;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:0 DR:11 LR:-16.26 LO:23.36);ALT=C[chr12:98993731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	98993905	+	chr12	98994947	+	.	13	20	5305224_1	85.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=25;MATEID=5305224_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_98980001_99005001_246C;SPAN=1042;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:75 GQ:85.4 PL:[85.4, 0.0, 95.3] SR:20 DR:13 LR:-85.31 LO:85.35);ALT=G[chr12:98994947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
