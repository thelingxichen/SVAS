chr19	382342	+	chr19	381011	+	.	16	0	10102941_1	20.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=10102941_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:381011(-)-19:382342(+)__19_367501_392501D;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:119 GQ:20.6 PL:[20.6, 0.0, 268.1] SR:0 DR:16 LR:-20.58 LO:33.22);ALT=]chr19:382342]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	396115	+	chr19	394906	+	.	34	0	10102576_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=10102576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:394906(-)-19:396115(+)__19_392001_417001D;SPAN=1209;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:0 DR:34 LR:-110.1 LO:110.1);ALT=]chr19:396115]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	668190	-	chr19	669809	+	.	8	0	10104048_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=10104048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:668190(-)-19:669809(-)__19_661501_686501D;SPAN=1619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:0 DR:8 LR:5.29 LO:14.13);ALT=[chr19:669809[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	1093675	-	chr19	1227293	+	.	5	13	10106146_1	28.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=10106146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1078001_1103001_0C;SPAN=133618;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:91 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:13 DR:5 LR:-28.16 LO:35.26);ALT=[chr19:1227293[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	1950289	+	chr19	1951814	+	.	34	0	10110082_1	94.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=10110082_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1950289(+)-19:1951814(-)__19_1935501_1960501D;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:65 GQ:61.7 PL:[94.7, 0.0, 61.7] SR:0 DR:34 LR:-94.96 LO:94.96);ALT=C[chr19:1951814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2909528	+	chr19	2910826	+	AGTCTTGACC	25	40	10116187_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=TCGTGATCCGCCCGCCTCGGCCTCC;INSERTION=AGTCTTGACC;MAPQ=0;MATEID=10116187_2;MATENM=2;NM=5;NUMPARTS=2;REPSEQ=CC;SCTG=c_19_2891001_2916001_420C;SECONDARY;SPAN=1298;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:107 GQ:96.5 PL:[162.5, 0.0, 96.5] SR:40 DR:25 LR:-163.3 LO:163.3);ALT=C[chr19:2910826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
