chr2	15694265	+	chr2	15698704	+	TACCAGATGTATTGGCGTAAAAATAATAAACGAT	0	11	698587_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TACCAGATGTATTGGCGTAAAAATAATAAACGAT;MAPQ=60;MATEID=698587_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_15680001_15705001_325C;SPAN=4439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:70 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:11 DR:0 LR:-17.35 LO:23.65);ALT=G[chr2:15698704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	15732073	+	chr2	15735614	+	AGATGGGTGTAATGCCTGAGATTGCACAAGCTGTGGAAGAGATGGATTGGCT	4	5	698897_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AGATGGGTGTAATGCCTGAGATTGCACAAGCTGTGGAAGAGATGGATTGGCT;MAPQ=60;MATEID=698897_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_15729001_15754001_110C;SPAN=3541;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:5 DR:4 LR:-2.296 LO:15.12);ALT=G[chr2:15735614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	15732073	+	chr2	15735268	+	.	2	5	698896_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=698896_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_15729001_15754001_110C;SPAN=3195;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:89 GQ:4.2 PL:[0.0, 4.2, 224.4] SR:5 DR:2 LR:4.306 LO:10.56);ALT=G[chr2:15735268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	16407988	+	chr2	16406393	+	CAGGCCC	46	42	700651_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=CAGGCCC;MAPQ=60;MATEID=700651_2;MATENM=13;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_2_16390501_16415501_123C;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:95 GQ:0.8 PL:[228.5, 0.0, 0.8] SR:42 DR:46 LR:-242.1 LO:242.1);ALT=]chr2:16407988]A;VARTYPE=BND:DUP-th;JOINTYPE=th
