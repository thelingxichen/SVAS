chr7	123185731	+	chr7	123190523	+	.	0	9	3562124_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=3562124_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_123186001_123211001_5C;SPAN=4792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:9 DR:0 LR:-15.89 LO:19.85);ALT=C[chr7:123190523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
