chr14	88391701	+	chr14	88393397	+	.	49	52	8662090_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTT;MAPQ=60;MATEID=8662090_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_14_88371501_88396501_369C;SPAN=1696;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:88 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:52 DR:49 LR:-260.8 LO:260.8);ALT=T[chr14:88393397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
