chr7	26163495	+	chr7	25823213	+	GA	81	26	4635943_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GA;MAPQ=60;MATEID=4635943_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26141501_26166501_479C;SPAN=340282;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:90 DP:149 GQ:99 PL:[256.7, 0.0, 104.9] SR:26 DR:81 LR:-260.2 LO:260.2);ALT=]chr7:26163495]T;VARTYPE=BND:DUP-th;JOINTYPE=th
