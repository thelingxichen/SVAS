chr20	19902780	-	chr20	19903794	+	.	4	2	10442678_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GATTACAGGCGTGAGC;MAPQ=60;MATEID=10442678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_19894001_19919001_30C;SPAN=1014;SUBN=10;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:6 DP:64 GQ:2.6 PL:[2.6, 0.0, 151.1] SR:2 DR:4 LR:-2.467 LO:11.46);ALT=[chr20:19903794[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
