chr5	4793562	-	chr5	4794774	+	.	8	0	3168931_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3168931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:4793562(-)-5:4794774(-)__5_4777501_4802501D;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:176 GQ:21.1 PL:[0.0, 21.1, 468.7] SR:0 DR:8 LR:21.27 LO:12.68);ALT=[chr5:4794774[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
