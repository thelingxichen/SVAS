chr12	133049439	+	chr12	133050780	+	.	8	0	7923347_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7923347_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:133049439(+)-12:133050780(-)__12_133035001_133060001D;SPAN=1341;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:0 DR:8 LR:-6.901 LO:15.9);ALT=C[chr12:133050780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133141112	+	chr12	133344211	-	.	31	46	7923836_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAGACTCCGTCTCCAAAAAAAAAA;MAPQ=60;MATEID=7923836_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_133133001_133158001_404C;SPAN=203099;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:21 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:46 DR:31 LR:-194.7 LO:194.7);ALT=C]chr12:133344211];VARTYPE=BND:INV-hh;JOINTYPE=hh
