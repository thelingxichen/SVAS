chr5	151456430	+	chr5	151462448	+	.	105	65	3847803_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAAAATTACATGGTGGA;MAPQ=60;MATEID=3847803_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_151459001_151484001_378C;SPAN=6018;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:148 DP:85 GQ:40 PL:[439.0, 40.0, 0.0] SR:65 DR:105 LR:-439.0 LO:439.0);ALT=A[chr5:151462448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
