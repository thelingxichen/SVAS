chr16	27236557	+	chr16	27238040	+	TTGGGATCTCGTGGGGCCAGTAGTCGTTGCAGTGGGGGCAGCGCGGTTCAGCATTCGACTGGAAGTACTTGGCCACGCAGGGTAAGTGCATCCTGATCCCACAGGTTTCGCAGCTTTGAC	2	33	6169795_1	87.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=TTGGGATCTCGTGGGGCCAGTAGTCGTTGCAGTGGGGGCAGCGCGGTTCAGCATTCGACTGGAAGTACTTGGCCACGCAGGGTAAGTGCATCCTGATCCCACAGGTTTCGCAGCTTTGAC;MAPQ=60;MATEID=6169795_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_27219501_27244501_20C;SPAN=1483;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:90 GQ:87.8 PL:[87.8, 0.0, 130.7] SR:33 DR:2 LR:-87.85 LO:88.31);ALT=T[chr16:27238040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	27238159	+	chr16	27244322	+	.	2	3	6169828_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6169828_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_27244001_27269001_289C;SPAN=6163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:41 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:3 DR:2 LR:-5.397 LO:10.15);ALT=T[chr16:27244322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	27244468	+	chr16	27246495	+	AGCCTTTCTAAACAAATCCAGTTCATTCTCTGCAAAATCCGTAGCCATTTTGGAAATTGAAGTTGTAGCAAGAT	2	22	6169832_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TCACC;INSERTION=AGCCTTTCTAAACAAATCCAGTTCATTCTCTGCAAAATCCGTAGCCATTTTGGAAATTGAAGTTGTAGCAAGAT;MAPQ=60;MATEID=6169832_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_27244001_27269001_334C;SPAN=2027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:81 GQ:57.5 PL:[57.5, 0.0, 136.7] SR:22 DR:2 LR:-57.28 LO:59.17);ALT=G[chr16:27246495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	27246620	+	chr16	27268755	+	.	0	50	6169922_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6169922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_27268501_27293501_0C;SPAN=22135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:50 DR:0 LR:-155.1 LO:155.1);ALT=C[chr16:27268755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	27246666	+	chr16	27280024	+	.	40	0	6169924_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6169924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:27246666(+)-16:27280024(-)__16_27268501_27293501D;SPAN=33358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:80 GQ:83.9 PL:[110.3, 0.0, 83.9] SR:0 DR:40 LR:-110.6 LO:110.6);ALT=A[chr16:27280024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	27268890	+	chr16	27280024	+	.	34	0	6169926_1	76.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6169926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:27268890(+)-16:27280024(-)__16_27268501_27293501D;SPAN=11134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:133 GQ:76.4 PL:[76.4, 0.0, 244.7] SR:0 DR:34 LR:-76.2 LO:81.23);ALT=A[chr16:27280024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
