chr6	70462248	+	chr6	70506704	+	TATAGTAACCGTATAATACAGTGTCCTCAATCTGTCTGCTGACATTAGCATTAGCCCAGTCCTTAAATGTACCATTTTGATTTTTCATGTAAGAAACCAAAAATATATCCACTGGTAGAAGTGCTGATGTGATAAGTGCAATTGCTAGAGAAAAAATTGCTGTTATGGTGGAGACAACTTCACTTTCCCGCCGACTTTGGTATTTACGAACATATATCCAGCAGAATGCCAAAATAG	0	12	2893260_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TATAGTAACCGTATAATACAGTGTCCTCAATCTGTCTGCTGACATTAGCATTAGCCCAGTCCTTAAATGTACCATTTTGATTTTTCATGTAAGAAACCAAAAATATATCCACTGGTAGAAGTGCTGATGTGATAAGTGCAATTGCTAGAGAAAAAATTGCTGTTATGGTGGAGACAACTTCACTTTCCCGCCGACTTTGGTATTTACGAACATATATCCAGCAGAATGCCAAAATAG;MAPQ=60;MATEID=2893260_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_70486501_70511501_35C;SPAN=44456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:37 GQ:29.6 PL:[29.6, 0.0, 59.3] SR:12 DR:0 LR:-29.59 LO:30.16);ALT=G[chr6:70506704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	70500365	+	chr6	70506704	+	.	25	5	2893293_1	50.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=2893293_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GTAGTA;SCTG=c_6_70486501_70511501_35C;SPAN=6339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:84 GQ:50.3 PL:[50.3, 0.0, 99.7] SR:5 DR:25 LR:-50.1 LO:51.24);ALT=C[chr6:70506704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	71377846	+	chr6	71442079	+	.	0	22	2895369_1	61.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=2895369_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_71442001_71467001_2C;SPAN=64233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:43 GQ:41.3 PL:[61.1, 0.0, 41.3] SR:22 DR:0 LR:-61.13 LO:61.13);ALT=T[chr6:71442079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	71442214	+	chr6	71464681	+	.	0	15	2895370_1	27.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2895370_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_71442001_71467001_234C;SPAN=22467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:80 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:15 DR:0 LR:-27.84 LO:33.52);ALT=G[chr6:71464681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	71874808	-	chr8	55014310	+	.	16	0	3864540_1	44.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=3864540_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:71874808(-)-8:55014310(-)__8_55002501_55027501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:33 GQ:34.1 PL:[44.0, 0.0, 34.1] SR:0 DR:16 LR:-43.91 LO:43.91);ALT=[chr8:55014310[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	54745646	+	chr8	54755594	+	TGAAGATAGGATTGCCAGTTGACTTTGTTTGCACGAACTTCTGCAGCCTTGGCAGCAATAATATTGGTGGGGACAGCAGCATCCACAGCACCTCGGATATCCATTTTGGTCATCTAAACTTCGTAATCTTGAATGTCTTTCAACAAAT	0	24	3863598_1	54.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGAAGATAGGATTGCCAGTTGACTTTGTTTGCACGAACTTCTGCAGCCTTGGCAGCAATAATATTGGTGGGGACAGCAGCATCCACAGCACCTCGGATATCCATTTTGGTCATCTAAACTTCGTAATCTTGAATGTCTTTCAACAAAT;MAPQ=60;MATEID=3863598_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_54733001_54758001_241C;SPAN=9948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:92 GQ:54.5 PL:[54.5, 0.0, 166.7] SR:24 DR:0 LR:-54.3 LO:57.58);ALT=C[chr8:54755594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	54754333	+	chr8	54755507	+	.	20	0	3863632_1	43.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3863632_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:54754333(+)-8:54755507(-)__8_54733001_54758001D;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:83 GQ:43.7 PL:[43.7, 0.0, 155.9] SR:0 DR:20 LR:-43.53 LO:47.18);ALT=T[chr8:54755507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	55047952	+	chr8	55049070	+	.	20	7	3864702_1	57.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3864702_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_55027001_55052001_120C;SPAN=1118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:81 GQ:57.5 PL:[57.5, 0.0, 136.7] SR:7 DR:20 LR:-57.28 LO:59.17);ALT=G[chr8:55049070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
