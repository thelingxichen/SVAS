chr4	56720119	+	chr4	56724479	+	.	0	7	1977360_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1977360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_56717501_56742501_76C;SPAN=4360;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:107 GQ:5.7 PL:[0.0, 5.7, 270.6] SR:7 DR:0 LR:5.882 LO:12.23);ALT=G[chr4:56724479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	56768706	+	chr4	56770507	+	.	3	2	1977581_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1977581_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_56766501_56791501_363C;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:94 GQ:12 PL:[0.0, 12.0, 250.8] SR:2 DR:3 LR:12.26 LO:6.224);ALT=T[chr4:56770507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57302494	+	chr4	57307828	+	.	38	8	1979427_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1979427_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57281001_57306001_271C;SPAN=5334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:52 GQ:3.9 PL:[132.0, 3.9, 0.0] SR:8 DR:38 LR:-136.2 LO:136.2);ALT=G[chr4:57307828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57333882	+	chr4	57337885	+	.	16	0	1979636_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1979636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:57333882(+)-4:57337885(-)__4_57330001_57355001D;SPAN=4003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:110 GQ:23 PL:[23.0, 0.0, 244.1] SR:0 DR:16 LR:-23.01 LO:33.81);ALT=C[chr4:57337885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57333910	+	chr4	57335819	+	.	37	15	1979637_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1979637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57330001_57355001_139C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:103 GQ:99 PL:[117.5, 0.0, 130.7] SR:15 DR:37 LR:-117.3 LO:117.4);ALT=A[chr4:57335819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57335939	+	chr4	57337886	+	.	0	43	1979641_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1979641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57330001_57355001_314C;SPAN=1947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:118 GQ:99 PL:[110.0, 0.0, 176.0] SR:43 DR:0 LR:-110.0 LO:110.8);ALT=A[chr4:57337886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57340557	+	chr4	57344545	+	AGTGTCTTCTGATAATGAACGGCGGCAAAGAT	2	10	1979662_1	13.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AGCCTCCTCTGTTCGACCCTGAAGCTGCAGAATATAAGCCATCTGACCATGAATGATGGCCAGTTCTGCCTGTGGGTCTTCCTCAGTCCCATCAGTGTCTTCTGATAATGAACGGCGGCAAAGATCT;INSERTION=AGTGTCTTCTGATAATGAACGGCGGCAAAGAT;MAPQ=60;MATEID=1979662_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_57330001_57355001_246C;SECONDARY;SPAN=3988;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:98 GQ:13.1 PL:[13.1, 0.0, 224.3] SR:10 DR:2 LR:-13.06 LO:24.39);ALT=G[chr4:57344545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57349437	+	chr4	57350900	+	.	4	8	1979695_1	8.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1979695_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57330001_57355001_209C;SPAN=1463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:117 GQ:8 PL:[8.0, 0.0, 275.3] SR:8 DR:4 LR:-7.914 LO:23.41);ALT=G[chr4:57350900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57514967	+	chr4	57522023	+	.	24	55	1980193_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=1980193_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57501501_57526501_233C;SPAN=7056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:122 GQ:86 PL:[208.1, 0.0, 86.0] SR:55 DR:24 LR:-210.6 LO:210.6);ALT=G[chr4:57522023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57515013	+	chr4	57522465	+	.	36	0	1980194_1	93.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1980194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:57515013(+)-4:57522465(-)__4_57501501_57526501D;SPAN=7452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:93 GQ:93.8 PL:[93.8, 0.0, 130.1] SR:0 DR:36 LR:-93.64 LO:94.0);ALT=A[chr4:57522465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57676351	+	chr4	57687669	+	GTTCTATATTTTGAAAACAGACCAAATTGAGGGATCAGAGAGG	55	32	1980881_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTCTATATTTTGAAAACAGACCAAATTGAGGGATCAGAGAGG;MAPQ=60;MATEID=1980881_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_57673001_57698001_159C;SPAN=11318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:620 GQ:99 PL:[119.3, 0.0, 1387.0] SR:32 DR:55 LR:-119.2 LO:182.4);ALT=C[chr4:57687669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57676353	+	chr4	57677850	+	.	8	82	1980883_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=1980883_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57673001_57698001_164C;SPAN=1497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:502 GQ:99 PL:[158.1, 0.0, 1059.0] SR:82 DR:8 LR:-157.8 LO:196.5);ALT=G[chr4:57677850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57678023	+	chr4	57687778	+	.	105	0	1980896_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1980896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:57678023(+)-4:57687778(-)__4_57673001_57698001D;SPAN=9755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:105 DP:225 GQ:99 PL:[285.8, 0.0, 259.4] SR:0 DR:105 LR:-285.7 LO:285.7);ALT=G[chr4:57687778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57686748	+	chr4	57687774	+	.	5	22	1980941_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=1980941_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_57673001_57698001_209C;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:27 DP:373 GQ:11.6 PL:[0.0, 11.6, 927.5] SR:22 DR:5 LR:11.93 LO:48.39);ALT=G[chr4:57687774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57845170	+	chr4	57852519	+	.	20	11	1981754_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1981754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57844501_57869501_283C;SPAN=7349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:106 GQ:44 PL:[44.0, 0.0, 212.3] SR:11 DR:20 LR:-43.9 LO:50.26);ALT=G[chr4:57852519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57845183	+	chr4	57856909	+	.	21	0	1981755_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1981755_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:57845183(+)-4:57856909(-)__4_57844501_57869501D;SPAN=11726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:110 GQ:39.5 PL:[39.5, 0.0, 227.6] SR:0 DR:21 LR:-39.52 LO:47.12);ALT=T[chr4:57856909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57852592	+	chr4	57856911	+	.	0	19	1981789_1	32.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1981789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57844501_57869501_398C;SPAN=4319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:113 GQ:32.3 PL:[32.3, 0.0, 240.2] SR:19 DR:0 LR:-32.1 LO:41.46);ALT=G[chr4:57856911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57897504	+	chr4	57898590	+	.	5	65	1981984_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=1981984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57893501_57918501_144C;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:133 GQ:99 PL:[191.9, 0.0, 129.2] SR:65 DR:5 LR:-192.3 LO:192.3);ALT=T[chr4:57898590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	57899479	+	chr4	57906988	+	.	6	7	1981995_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=1981995_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_57893501_57918501_199C;SPAN=7509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:122 GQ:3.5 PL:[3.5, 0.0, 290.6] SR:7 DR:6 LR:-3.258 LO:20.81);ALT=T[chr4:57906988[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
