chr8	17859520	-	chr9	105073654	+	.	16	18	5948076_1	92.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5948076_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_105056001_105081001_96C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:32 DP:25 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:18 DR:16 LR:-92.42 LO:92.42);ALT=[chr9:105073654[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	18454620	+	chr8	18455945	+	.	77	53	5407801_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAGGATC;MAPQ=60;MATEID=5407801_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_8_18448501_18473501_238C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:36 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:53 DR:77 LR:-316.9 LO:316.9);ALT=C[chr8:18455945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69675178	+	chr9	105936345	+	.	4	7	5949272_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATAT;MAPQ=60;MATEID=5949272_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_105913501_105938501_10C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:11 DP:5 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:7 DR:4 LR:-29.71 LO:29.71);ALT=]chr15:69675178]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	138479103	+	chr9	138480200	+	.	175	98	6041803_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGC;MAPQ=60;MATEID=6041803_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_9_138474001_138499001_305C;SPAN=1097;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:256 DP:44 GQ:69.1 PL:[759.1, 69.1, 0.0] SR:98 DR:175 LR:-759.2 LO:759.2);ALT=C[chr9:138480200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139054512	+	chr9	139059015	+	.	149	65	6046029_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=GCCTGTAGTCCCAGCTACTCGGGAGGC;MAPQ=38;MATEID=6046029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_139037501_139062501_102C;SPAN=4503;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:197 DP:60 GQ:53.2 PL:[584.2, 53.2, 0.0] SR:65 DR:149 LR:-584.2 LO:584.2);ALT=C[chr9:139059015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139542605	-	chr9	139544318	+	.	8	0	6048374_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6048374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139542605(-)-9:139544318(-)__9_139527501_139552501D;SPAN=1713;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:213 GQ:31 PL:[0.0, 31.0, 577.6] SR:0 DR:8 LR:31.3 LO:12.01);ALT=[chr9:139544318[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	140380858	+	chr9	140382863	+	G	0	8	6052846_1	0	.	EVDNC=ASSMB;INSERTION=G;MAPQ=60;MATEID=6052846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140360501_140385501_46C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:218 GQ:32.5 PL:[0.0, 32.5, 594.1] SR:8 DR:0 LR:32.65 LO:11.93);ALT=A[chr9:140382863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140739167	+	chr17	78375744	+	.	10	0	6056681_1	8.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6056681_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:140739167(+)-17:78375744(-)__9_140728001_140753001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:0 DR:10 LR:-8.898 LO:19.93);ALT=G[chr17:78375744[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr15	67827798	-	chr15	67828941	+	.	8	0	8950677_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=8950677_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:67827798(-)-15:67828941(-)__15_67816001_67841001D;SPAN=1143;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:174 GQ:20.5 PL:[0.0, 20.5, 462.1] SR:0 DR:8 LR:20.73 LO:12.72);ALT=[chr15:67828941[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	68247957	+	chr15	68047969	+	GTTTGAACATGGGTCAGATGGTCTCTCTCCAGGGCCTGACGGTGAGAGGTGCAGCCT	58	85	8953074_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GTTTGAACATGGGTCAGATGGTCTCTCTCCAGGGCCTGACGGTGAGAGGTGCAGCCT;MAPQ=60;MATEID=8953074_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_68232501_68257501_61C;SPAN=199988;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:136 DP:100 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:85 DR:58 LR:-402.7 LO:402.7);ALT=]chr15:68247957]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	68047969	-	chr15	68152479	+	.	21	28	8952275_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;MAPQ=60;MATEID=8952275_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_15_68134501_68159501_194C;SPAN=104510;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:72 GQ:69.8 PL:[102.8, 0.0, 69.8] SR:28 DR:21 LR:-102.9 LO:102.9);ALT=[chr15:68152479[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	68116010	+	chr15	68152570	+	TG	49	17	8952276_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TG;MAPQ=60;MATEID=8952276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_68134501_68159501_286C;SPAN=36560;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:59 DP:104 GQ:84.2 PL:[166.7, 0.0, 84.2] SR:17 DR:49 LR:-168.0 LO:168.0);ALT=C[chr15:68152570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	68152536	+	chr15	68247957	-	.	17	72	8953077_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=8953077_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_68232501_68257501_61C;SPAN=95421;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:78 DP:100 GQ:12.5 PL:[230.3, 0.0, 12.5] SR:72 DR:17 LR:-242.1 LO:242.1);ALT=G]chr15:68247957];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr15	68426020	+	chr15	68428928	+	.	131	89	8954360_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTGAAATTTAGATTTTTA;MAPQ=60;MATEID=8954360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_68404001_68429001_370C;SPAN=2908;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:178 DP:50 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:89 DR:131 LR:-528.1 LO:528.1);ALT=A[chr15:68428928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69257918	+	chr17	78511823	+	GAGAGG	6	19	8958083_1	55.0	.	DISC_MAPQ=11;EVDNC=ASDIS;INSERTION=GAGAGG;MAPQ=19;MATEID=8958083_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_69237001_69262001_210C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:87 GQ:55.7 PL:[55.7, 0.0, 154.7] SR:19 DR:6 LR:-55.65 LO:58.27);ALT=G[chr17:78511823[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr17	77779887	+	chr17	77781124	-	.	8	0	9833278_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9833278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:77779887(+)-17:77781124(+)__17_77763001_77788001D;SPAN=1237;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=G]chr17:77781124];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	77995767	+	chr17	77998937	+	.	18	0	9834782_1	17.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=9834782_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:77995767(+)-17:77998937(-)__17_77983501_78008501D;SPAN=3170;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:157 GQ:17 PL:[17.0, 0.0, 363.5] SR:0 DR:18 LR:-16.88 LO:36.04);ALT=C[chr17:77998937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	78461849	+	chr17	78463568	+	.	10	0	9836885_1	22.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=9836885_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:78461849(+)-17:78463568(-)__17_78449001_78474001D;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:41 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-21.9 LO:23.65);ALT=A[chr17:78463568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
