chr11	122347584	+	chr11	122349281	+	.	170	88	7236565_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAGAAAG;MAPQ=60;MATEID=7236565_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_11_122328501_122353501_410C;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:220 DP:81 GQ:59.5 PL:[653.5, 59.5, 0.0] SR:88 DR:170 LR:-653.6 LO:653.6);ALT=G[chr11:122349281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
