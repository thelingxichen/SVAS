chr3	36433996	-	chr3	36435389	+	.	9	0	1945526_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1945526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:36433996(-)-3:36435389(-)__3_36431501_36456501D;SPAN=1393;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:127 GQ:4.5 PL:[0.0, 4.5, 316.8] SR:0 DR:9 LR:4.698 LO:16.05);ALT=[chr3:36435389[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
