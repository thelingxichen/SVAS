chr7	20764210	-	chr7	20766079	+	.	8	0	4599469_1	0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=4599469_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:20764210(-)-7:20766079(-)__7_20751501_20776501D;SPAN=1869;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:205 GQ:28.9 PL:[0.0, 28.9, 554.5] SR:0 DR:8 LR:29.13 LO:12.14);ALT=[chr7:20766079[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
