chr3	95465768	+	chr3	95470764	+	.	35	42	2179217_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CAAG;MAPQ=60;MATEID=2179217_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_319C;SPAN=4996;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:66 DP:119 GQ:99 PL:[185.6, 0.0, 103.1] SR:42 DR:35 LR:-186.9 LO:186.9);ALT=G[chr3:95470764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	95465790	+	chr3	95468114	+	.	18	0	2179218_1	40.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2179218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:95465790(+)-3:95468114(-)__3_95452001_95477001D;SPAN=2324;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:70 GQ:40.4 PL:[40.4, 0.0, 129.5] SR:0 DR:18 LR:-40.45 LO:43.06);ALT=T[chr3:95468114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	95471000	+	chr3	95468117	+	TGCATAGGG	42	38	2179223_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGCATAGGG;MAPQ=60;MATEID=2179223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_15C;SPAN=2883;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:118 GQ:99 PL:[179.3, 0.0, 106.7] SR:38 DR:42 LR:-180.3 LO:180.3);ALT=]chr3:95471000]A;VARTYPE=BND:DUP-th;JOINTYPE=th
