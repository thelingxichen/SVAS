chr18	29598990	+	chr18	29617079	+	.	21	30	6579445_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6579445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_29596001_29621001_145C;SPAN=18089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:89 GQ:99 PL:[104.6, 0.0, 111.2] SR:30 DR:21 LR:-104.6 LO:104.6);ALT=T[chr18:29617079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	29617234	+	chr18	29622141	+	.	0	7	6579504_1	11.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=6579504_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_29620501_29645501_275C;SPAN=4907;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:44 GQ:11.3 PL:[11.3, 0.0, 93.8] SR:7 DR:0 LR:-11.19 LO:15.09);ALT=T[chr18:29622141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
