chr1	60046769	+	chr1	60050636	+	.	43	0	291937_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=291937_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:60046769(+)-1:60050636(-)__1_60049501_60074501D;SPAN=3867;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:46 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:0 DR:43 LR:-135.3 LO:135.3);ALT=A[chr1:60050636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
