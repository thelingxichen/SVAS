chr1	217793853	+	chr1	217804310	+	.	9	0	549253_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=549253_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:217793853(+)-1:217804310(-)__1_217780501_217805501D;SPAN=10457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:129 GQ:5.1 PL:[0.0, 5.1, 323.4] SR:0 DR:9 LR:5.24 LO:15.98);ALT=A[chr1:217804310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	218182502	+	chr1	218188595	+	.	93	62	550809_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TATTTTGACTTCTT;MAPQ=60;MATEID=550809_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_218172501_218197501_252C;SPAN=6093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:50 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:62 DR:93 LR:-366.4 LO:366.4);ALT=T[chr1:218188595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	218458798	+	chr1	218475634	+	.	0	9	551197_1	14.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=551197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_218442001_218467001_100C;SPAN=16836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:9 DR:0 LR:-14.0 LO:19.3);ALT=G[chr1:218475634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
