chr10	112678389	+	chr10	112457972	+	.	3	2	6523955_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=6523955_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_112675501_112700501_283C;SPAN=220417;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:50 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:2 DR:3 LR:0.3422 LO:7.35);ALT=]chr10:112678389]T;VARTYPE=BND:DUP-th;JOINTYPE=th
