chr5	14404243	+	chr5	14402573	+	.	50	0	2419639_1	99.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2419639_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:14402573(-)-5:14404243(+)__5_14381501_14406501D;SPAN=1670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:80 GQ:50.9 PL:[143.3, 0.0, 50.9] SR:0 DR:50 LR:-145.8 LO:145.8);ALT=]chr5:14404243]T;VARTYPE=BND:DUP-th;JOINTYPE=th
