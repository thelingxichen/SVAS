chr4	46055996	+	chr4	46058203	+	A	24	14	1955762_1	52.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=1955762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_46035501_46060501_3C;SPAN=2207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:161 GQ:52.4 PL:[52.4, 0.0, 336.2] SR:14 DR:24 LR:-52.11 LO:64.25);ALT=T[chr4:46058203[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	46202797	+	chr4	46205027	+	.	35	43	1955738_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=1955738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_46182501_46207501_66C;SPAN=2230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:18 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:43 DR:35 LR:-181.5 LO:181.5);ALT=C[chr4:46205027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
