chr1	83125976	+	chr1	83127570	+	.	58	37	221559_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAAAATGGTTCATGC;MAPQ=60;MATEID=221559_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_1_83104001_83129001_216C;SPAN=1594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:22 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:37 DR:58 LR:-241.0 LO:241.0);ALT=C[chr1:83127570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
