chr7	50343780	+	chr7	50367229	+	.	8	0	3301850_1	21.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3301850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:50343780(+)-7:50367229(-)__7_50323001_50348001D;SPAN=23449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:21.5 PL:[21.5, 0.0, 21.5] SR:0 DR:8 LR:-21.53 LO:21.53);ALT=G[chr7:50367229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	50344407	+	chr7	50358643	+	.	22	0	3301852_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3301852_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:50344407(+)-7:50358643(-)__7_50323001_50348001D;SPAN=14236;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:73 GQ:53 PL:[53.0, 0.0, 122.3] SR:0 DR:22 LR:-52.84 LO:54.44);ALT=T[chr7:50358643[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	50344498	+	chr7	50367229	+	.	12	0	3301853_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3301853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:50344498(+)-7:50367229(-)__7_50323001_50348001D;SPAN=22731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:72 GQ:20.3 PL:[20.3, 0.0, 152.3] SR:0 DR:12 LR:-20.11 LO:26.14);ALT=A[chr7:50367229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
