chr5	101726323	-	chr5	101735627	+	CATTAATGAATGAAACATTAATGACTAACA	39	44	2541862_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CATTAATGAATGAAACATTAATGACTAACA;MAPQ=60;MATEID=2541862_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_5_101724001_101749001_172C;SPAN=9304;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:43 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:44 DR:39 LR:-194.7 LO:194.7);ALT=[chr5:101735627[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	101727275	+	chr5	101730115	-	.	40	0	2541867_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2541867_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:101727275(+)-5:101730115(+)__5_101724001_101749001D;SPAN=2840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:25 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:40 LR:-118.8 LO:118.8);ALT=A]chr5:101730115];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	102456194	+	chr5	102465008	+	.	39	15	2542935_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2542935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_102459001_102484001_6C;SPAN=8814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:25 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:15 DR:39 LR:-135.3 LO:135.3);ALT=T[chr5:102465008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	102487078	+	chr5	102488351	+	.	0	8	2542899_1	13.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=2542899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_102483501_102508501_59C;SPAN=1273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:8 DR:0 LR:-13.13 LO:17.35);ALT=G[chr5:102488351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
