chr4	118579744	+	chr4	118591109	+	.	8	0	2168122_1	14.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2168122_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:118579744(+)-4:118591109(-)__4_118580001_118605001D;SPAN=11365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=T[chr4:118591109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
