chr2	49750842	+	chr2	49649169	+	.	5	7	990606_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=990606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_49735001_49760001_110C;SPAN=101673;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:31 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:7 DR:5 LR:-24.61 LO:25.11);ALT=]chr2:49750842]T;VARTYPE=BND:DUP-th;JOINTYPE=th
