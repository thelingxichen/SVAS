chr6	45872386	+	chr1	47804186	+	.	2	43	4181974_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TCCCT;MAPQ=60;MATEID=4181974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_45864001_45889001_132C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:45 DP:33 GQ:12 PL:[132.0, 12.0, 0.0] SR:43 DR:2 LR:-132.0 LO:132.0);ALT=]chr6:45872386]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	44992731	+	chr6	44946880	+	A	4	7	4178710_1	1.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4178710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44982001_45007001_251C;SPAN=45851;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:79 GQ:1.7 PL:[1.7, 0.0, 189.8] SR:7 DR:4 LR:-1.704 LO:13.19);ALT=]chr6:44992731]T;VARTYPE=BND:DUP-th;JOINTYPE=th
