chr11	132865750	+	chr11	132867628	+	.	0	8	7302572_1	0	.	EVDNC=ASSMB;HOMSEQ=GATTCCAAG;MAPQ=60;MATEID=7302572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_132863501_132888501_442C;SPAN=1878;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:216 GQ:31.9 PL:[0.0, 31.9, 587.5] SR:8 DR:0 LR:32.11 LO:11.96);ALT=G[chr11:132867628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
