chr8	85177892	+	chr10	122156528	+	.	21	48	4705123_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;MAPQ=60;MATEID=4705123_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_122132501_122157501_6C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:40 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:48 DR:21 LR:-158.4 LO:158.4);ALT=T[chr10:122156528[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	85865342	+	chr8	85874154	-	.	11	0	3947744_1	29.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=3947744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:85865342(+)-8:85874154(+)__8_85872501_85897501D;SPAN=8812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=A]chr8:85874154];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	86127280	+	chr8	86132533	+	.	29	0	3948574_1	74.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3948574_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:86127280(+)-8:86132533(-)__8_86117501_86142501D;SPAN=5253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:81 GQ:74 PL:[74.0, 0.0, 120.2] SR:0 DR:29 LR:-73.78 LO:74.45);ALT=A[chr8:86132533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	86129732	+	chr8	86132535	+	.	44	1	3948579_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=C;MAPQ=36;MATEID=3948579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_86117501_86142501_320C;SPAN=2803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:108 GQ:99 PL:[119.3, 0.0, 142.4] SR:1 DR:44 LR:-119.3 LO:119.4);ALT=C[chr8:86132535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	86376321	+	chr8	86377499	+	.	16	0	3949128_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3949128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:86376321(+)-8:86377499(-)__8_86362501_86387501D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:94 GQ:27.5 PL:[27.5, 0.0, 199.1] SR:0 DR:16 LR:-27.35 LO:35.01);ALT=A[chr8:86377499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120095935	+	chr10	120101239	+	.	0	17	4701553_1	48.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4701553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120099001_120124001_33C;SPAN=5304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:28 GQ:18.8 PL:[48.5, 0.0, 18.8] SR:17 DR:0 LR:-49.21 LO:49.21);ALT=T[chr10:120101239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120095963	+	chr10	120101781	+	.	17	0	4701554_1	46.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4701554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120095963(+)-10:120101781(-)__10_120099001_120124001D;SPAN=5818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:35 GQ:36.8 PL:[46.7, 0.0, 36.8] SR:0 DR:17 LR:-46.68 LO:46.68);ALT=T[chr10:120101781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120797954	+	chr10	120801504	+	.	9	11	4702646_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=4702646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120785001_120810001_158C;SPAN=3550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:56 GQ:37.7 PL:[37.7, 0.0, 97.1] SR:11 DR:9 LR:-37.64 LO:39.14);ALT=G[chr10:120801504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120802284	+	chr10	120803565	+	.	4	7	4702653_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4702653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120785001_120810001_166C;SPAN=1281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:64 GQ:19.1 PL:[19.1, 0.0, 134.6] SR:7 DR:4 LR:-18.97 LO:24.12);ALT=C[chr10:120803565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120802329	+	chr10	120809311	+	.	8	0	4702654_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4702654_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120802329(+)-10:120809311(-)__10_120785001_120810001D;SPAN=6982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:0 DR:8 LR:-10.97 LO:16.77);ALT=C[chr10:120809311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120810833	+	chr10	120816252	+	.	0	14	4702805_1	32.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4702805_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120809501_120834501_90C;SPAN=5419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:49 GQ:32.9 PL:[32.9, 0.0, 85.7] SR:14 DR:0 LR:-32.94 LO:34.25);ALT=T[chr10:120816252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120816552	+	chr10	120818724	+	TTCAATATCAATATCTTTGAATGCTTTGGCACCCAGTTCTGTTTTCTTGATCTGCTCCAAACGCTCTCGGACAGTTTTCTTTTTGATTTGTTCATGTTCCTGTAAGATACGCTCCTTCTCTCTCTCCTTTGCTTCCTGGCGCAGCCTCTCTTCCTCAGCCTTCCGCACTTTCTGGAGTTCAGCTTCCCTCTGTTCCAATTCTTCTTTCTCACGCTGAATATTCAGACTCTCAAGGCGCTCTTTTCTCTCCTCAATTGTCTGGCGGCGAGCCAGGATCCGCTGGTGCTCTTTTCGTGAATTTTTAAGGTATGCAGTGACAGCCAACTGATGCTGTTCTTCTTTCTCTTG	0	17	4702822_1	39.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTCAATATCAATATCTTTGAATGCTTTGGCACCCAGTTCTGTTTTCTTGATCTGCTCCAAACGCTCTCGGACAGTTTTCTTTTTGATTTGTTCATGTTCCTGTAAGATACGCTCCTTCTCTCTCTCCTTTGCTTCCTGGCGCAGCCTCTCTTCCTCAGCCTTCCGCACTTTCTGGAGTTCAGCTTCCCTCTGTTCCAATTCTTCTTTCTCACGCTGAATATTCAGACTCTCAAGGCGCTCTTTTCTCTCCTCAATTGTCTGGCGGCGAGCCAGGATCCGCTGGTGCTCTTTTCGTGAATTTTTAAGGTATGCAGTGACAGCCAACTGATGCTGTTCTTCTTTCTCTTG;MAPQ=60;MATEID=4702822_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_120809501_120834501_152C;SPAN=2172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:63 GQ:39.2 PL:[39.2, 0.0, 111.8] SR:17 DR:0 LR:-39.05 LO:41.08);ALT=C[chr10:120818724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120833450	+	chr10	120840140	+	.	22	25	4702855_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4702855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120809501_120834501_45C;SPAN=6690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:26 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:25 DR:22 LR:-105.6 LO:105.6);ALT=C[chr10:120840140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120921926	+	chr10	120923642	+	.	0	19	4703033_1	44.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4703033_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120907501_120932501_137C;SPAN=1716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:69 GQ:44 PL:[44.0, 0.0, 123.2] SR:19 DR:0 LR:-44.03 LO:46.12);ALT=C[chr10:120923642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120921971	+	chr10	120924746	+	.	9	0	4703035_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4703035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120921971(+)-10:120924746(-)__10_120907501_120932501D;SPAN=2775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:60 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.45 LO:19.15);ALT=T[chr10:120924746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120923709	+	chr10	120924714	+	.	0	9	4703041_1	12.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4703041_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120907501_120932501_280C;SPAN=1005;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:63 GQ:12.8 PL:[12.8, 0.0, 138.2] SR:9 DR:0 LR:-12.64 LO:18.94);ALT=C[chr10:120924714[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120923748	+	chr10	120925111	+	.	8	0	4703042_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4703042_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120923748(+)-10:120925111(-)__10_120907501_120932501D;SPAN=1363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:0 DR:8 LR:-9.34 LO:16.4);ALT=A[chr10:120925111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120934104	+	chr10	120936531	+	.	0	79	4703128_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=4703128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_120932001_120957001_287C;SPAN=2427;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:79 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:79 DR:0 LR:-234.4 LO:234.4);ALT=C[chr10:120936531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120934134	+	chr10	120938263	+	.	62	0	4703130_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=4703130_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120934134(+)-10:120938263(-)__10_120932001_120957001D;SPAN=4129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:73 GQ:9.6 PL:[194.7, 9.6, 0.0] SR:0 DR:62 LR:-198.5 LO:198.5);ALT=T[chr10:120938263[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	120936677	+	chr10	120938263	+	.	44	0	4703140_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=4703140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:120936677(+)-10:120938263(-)__10_120932001_120957001D;SPAN=1586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:67 GQ:34.7 PL:[127.1, 0.0, 34.7] SR:0 DR:44 LR:-130.0 LO:130.0);ALT=A[chr10:120938263[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121259773	+	chr10	121275021	+	.	3	13	4703686_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4703686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_121275001_121300001_201C;SPAN=15248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:32 GQ:34.4 PL:[41.0, 0.0, 34.4] SR:13 DR:3 LR:-40.86 LO:40.86);ALT=T[chr10:121275021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121275167	+	chr10	121285544	+	.	0	26	4703688_1	70.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4703688_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_121275001_121300001_228C;SPAN=10377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:57 GQ:67.1 PL:[70.4, 0.0, 67.1] SR:26 DR:0 LR:-70.39 LO:70.39);ALT=G[chr10:121285544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121275223	+	chr10	121302110	+	.	12	0	4703905_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4703905_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:121275223(+)-10:121302110(-)__10_121299501_121324501D;SPAN=26887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:24 GQ:23.3 PL:[33.2, 0.0, 23.3] SR:0 DR:12 LR:-33.17 LO:33.17);ALT=C[chr10:121302110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121285631	+	chr10	121286817	+	.	0	51	4703722_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4703722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_121275001_121300001_284C;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:66 GQ:8.6 PL:[150.5, 0.0, 8.6] SR:51 DR:0 LR:-157.8 LO:157.8);ALT=C[chr10:121286817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121285674	+	chr10	121302106	+	.	34	0	4703906_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4703906_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:121285674(+)-10:121302106(-)__10_121299501_121324501D;SPAN=16432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:20 GQ:9 PL:[99.0, 9.0, 0.0] SR:0 DR:34 LR:-99.02 LO:99.02);ALT=A[chr10:121302106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121286939	+	chr10	121302102	+	.	70	19	4703908_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4703908_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_121299501_121324501_6C;SPAN=15163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:19 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:19 DR:70 LR:-221.2 LO:221.2);ALT=G[chr10:121302102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121342071	+	chr10	121355946	+	CTGTTATCATTTTACAGCTTTTACAGGGTCCAATCTGACTGAACAACTGAAGTATAAGGACTTCTGTCACATCTCTGGAAAGGTTACCTACGTAT	0	15	4703776_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTGTTATCATTTTACAGCTTTTACAGGGTCCAATCTGACTGAACAACTGAAGTATAAGGACTTCTGTCACATCTCTGGAAAGGTTACCTACGTAT;MAPQ=60;MATEID=4703776_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_121324001_121349001_107C;SPAN=13875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:24 GQ:13.4 PL:[43.1, 0.0, 13.4] SR:15 DR:0 LR:-43.74 LO:43.74);ALT=T[chr10:121355946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	121347760	+	chr10	121355946	+	.	0	9	4703795_1	22.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4703795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_121348501_121373501_108C;SPAN=8186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:9 DR:0 LR:-22.39 LO:22.75);ALT=T[chr10:121355946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	122226687	+	chr10	122228789	+	.	42	0	4705478_1	99.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4705478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:122226687(+)-10:122228789(-)__10_122206001_122231001D;SPAN=2102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:19 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=T[chr10:122228789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
