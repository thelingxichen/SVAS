chr4	118096787	-	chr4	118097830	+	.	8	2	2865957_1	0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=TTTGGTTTTCTG;MAPQ=26;MATEID=2865957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_118090001_118115001_50C;SPAN=1043;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:145 GQ:6 PL:[0.0, 6.0, 363.0] SR:2 DR:8 LR:6.274 LO:17.71);ALT=[chr4:118097830[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	118579766	+	chr4	118591109	+	.	9	0	2868369_1	13.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2868369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:118579766(+)-4:118591109(-)__4_118580001_118605001D;SPAN=11343;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:59 GQ:13.7 PL:[13.7, 0.0, 129.2] SR:0 DR:9 LR:-13.72 LO:19.22);ALT=C[chr4:118591109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
