chr17	45175807	+	chr17	44287866	+	ATTAAAGTTTTTTTTT	53	87	9673731_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=ATTAAAGTTTTTTTTT;MAPQ=60;MATEID=9673731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_44271501_44296501_338C;SPAN=887941;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:135 DP:35 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:87 DR:53 LR:-399.4 LO:399.4);ALT=]chr17:45175807]A;VARTYPE=BND:DUP-th;JOINTYPE=th
