chrX	155187867	+	chrX	154871055	+	.	21	0	11435619_1	62.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=11435619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154871055(-)-23:155187867(+)__23_155183001_155208001D;SPAN=316812;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:21 DP:22 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:0 DR:21 LR:-62.72 LO:62.72);ALT=]chrX:155187867]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	154871535	+	chrX	155188331	+	.	9	0	11435620_1	23.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=11435620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:154871535(+)-23:155188331(-)__23_155183001_155208001D;SPAN=316796;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:0 DR:9 LR:-23.21 LO:23.34);ALT=A[chrX:155188331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	155216765	+	chrX	155033311	+	.	48	0	11436071_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=11436071_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:155033311(-)-23:155216765(+)__23_155207501_155232501D;SPAN=183454;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:0 DR:48 LR:-155.1 LO:155.1);ALT=]chrX:155216765]C;VARTYPE=BND:DUP-th;JOINTYPE=th
