chr6	47301087	+	chr6	46988761	+	TATACATACACACACACACAG	0	60	4188833_1	99.0	.	EVDNC=ASSMB;INSERTION=TATACATACACACACACACAG;MAPQ=60;MATEID=4188833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_47285001_47310001_41C;SPAN=312326;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:62 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:60 DR:0 LR:-181.5 LO:181.5);ALT=]chr6:47301087]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	47183544	+	chr6	47185561	-	.	10	0	4187792_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4187792_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:47183544(+)-6:47185561(+)__6_47162501_47187501D;SPAN=2017;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:203 GQ:21.7 PL:[0.0, 21.7, 534.7] SR:0 DR:10 LR:21.99 LO:16.21);ALT=G]chr6:47185561];VARTYPE=BND:INV-hh;JOINTYPE=hh
