chr1	89652020	+	chr1	89598982	+	.	8	0	410113_1	11.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=410113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:89598982(-)-1:89652020(+)__1_89645501_89670501D;SPAN=53038;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:0 DR:8 LR:-10.97 LO:16.77);ALT=]chr1:89652020]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	90354847	-	chr1	90356633	+	.	9	0	413012_1	13.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=413012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:90354847(-)-1:90356633(-)__1_90331501_90356501D;SPAN=1786;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:61 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.18 LO:19.08);ALT=[chr1:90356633[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
