chr9	78919603	+	chr9	78922019	+	.	14	0	4282998_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4282998_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:78919603(+)-9:78922019(-)__9_78914501_78939501D;SPAN=2416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:60 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:0 DR:14 LR:-29.96 LO:32.8);ALT=C[chr9:78922019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	79074231	+	chr9	79115828	+	.	10	0	4283670_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4283670_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:79074231(+)-9:79115828(-)__9_79110501_79135501D;SPAN=41597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=T[chr9:79115828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	79074246	+	chr9	79076213	+	.	12	0	4283630_1	9.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4283630_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:79074246(+)-9:79076213(-)__9_79061501_79086501D;SPAN=1967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:111 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:0 DR:12 LR:-9.539 LO:23.7);ALT=C[chr9:79076213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	79075093	+	chr9	79076214	+	.	0	4	4283632_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4283632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_79061501_79086501_139C;SPAN=1121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:108 GQ:15.9 PL:[0.0, 15.9, 293.7] SR:4 DR:0 LR:16.06 LO:5.98);ALT=G[chr9:79076214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
