chr2	240488047	+	chr2	240486851	+	.	16	0	1259527_1	28.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1259527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:240486851(-)-2:240488047(+)__2_240467501_240492501D;SPAN=1196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:90 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:0 DR:16 LR:-28.43 LO:35.35);ALT=]chr2:240488047]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	240900605	+	chr2	240929491	+	.	0	7	1260478_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1260478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_240908501_240933501_358C;SPAN=28886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:7 DR:0 LR:-10.37 LO:14.87);ALT=T[chr2:240929491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	240960882	+	chr2	240964681	+	.	17	0	1260747_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1260747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:240960882(+)-2:240964681(-)__2_240957501_240982501D;SPAN=3799;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:88 GQ:32.3 PL:[32.3, 0.0, 180.8] SR:0 DR:17 LR:-32.28 LO:38.24);ALT=A[chr2:240964681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	240961758	+	chr2	240964644	+	.	65	9	1260749_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1260749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_240957501_240982501_220C;SPAN=2886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:62 GQ:18 PL:[198.0, 18.0, 0.0] SR:9 DR:65 LR:-198.0 LO:198.0);ALT=C[chr2:240964644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	241070574	+	chr2	241075641	+	.	68	0	1260963_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1260963_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:241070574(+)-2:241075641(-)__2_241055501_241080501D;SPAN=5067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:56 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:0 DR:68 LR:-201.3 LO:201.3);ALT=G[chr2:241075641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	241073424	+	chr2	241075638	+	.	23	22	1260969_1	98.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1260969_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_241055501_241080501_303C;SPAN=2214;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:75 GQ:82.1 PL:[98.6, 0.0, 82.1] SR:22 DR:23 LR:-98.58 LO:98.58);ALT=T[chr2:241075638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	241564979	+	chr2	241569363	+	ATG	7	2	1262141_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATG;MAPQ=60;MATEID=1262141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_241545501_241570501_46C;SPAN=4384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:2 DR:7 LR:-3.059 LO:13.4);ALT=C[chr2:241569363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242039312	+	chr2	242041666	+	.	10	5	1263202_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=1263202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_242035501_242060501_178C;SPAN=2354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:93 GQ:14.6 PL:[14.6, 0.0, 209.3] SR:5 DR:10 LR:-14.42 LO:24.68);ALT=G[chr2:242041666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242089987	+	chr2	242097227	+	.	14	0	1263581_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1263581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242089987(+)-2:242097227(-)__2_242084501_242109501D;SPAN=7240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:0 DR:14 LR:-21.29 LO:29.89);ALT=C[chr2:242097227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242089987	+	chr2	242092889	+	.	17	0	1263580_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1263580_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242089987(+)-2:242092889(-)__2_242084501_242109501D;SPAN=2902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:96 GQ:30.2 PL:[30.2, 0.0, 201.8] SR:0 DR:17 LR:-30.11 LO:37.52);ALT=C[chr2:242092889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242093019	+	chr2	242098626	+	AAGAACATGAGCTGCCTGTGGACATGGAAACCATCAACCTGGACAGAGATGCAGAGGATGTTGATTTGAATCACTATCGCATAGGGAAGATTGAAGGATTTGAGGTACTGAAGAAAGTGA	0	38	1263591_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAGAACATGAGCTGCCTGTGGACATGGAAACCATCAACCTGGACAGAGATGCAGAGGATGTTGATTTGAATCACTATCGCATAGGGAAGATTGAAGGATTTGAGGTACTGAAGAAAGTGA;MAPQ=60;MATEID=1263591_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_242084501_242109501_292C;SPAN=5607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:89 GQ:99 PL:[101.3, 0.0, 114.5] SR:38 DR:0 LR:-101.3 LO:101.4);ALT=G[chr2:242098626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242102816	+	chr2	242105747	+	.	2	18	1263622_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGCAG;MAPQ=60;MATEID=1263622_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_242084501_242109501_65C;SPAN=2931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:87 GQ:39.2 PL:[39.2, 0.0, 171.2] SR:18 DR:2 LR:-39.15 LO:43.89);ALT=G[chr2:242105747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242204022	+	chr2	242207892	+	TTGATTTGTTGCGGAACCAGCCCACTTCGGTGTTCAGCAAAACTCTCTTGGGTCAAAACTGCAACGGAACTCATGGTTGATCTCACACCTACACACAATCCGGGAAAACCA	0	24	1264044_1	70.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTGATTTGTTGCGGAACCAGCCCACTTCGGTGTTCAGCAAAACTCTCTTGGGTCAAAACTGCAACGGAACTCATGGTTGATCTCACACCTACACACAATCCGGGAAAACCA;MAPQ=60;MATEID=1264044_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_2_242182501_242207501_294C;SPAN=3870;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:33 GQ:7.7 PL:[70.4, 0.0, 7.7] SR:24 DR:0 LR:-72.91 LO:72.91);ALT=T[chr2:242207892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242204022	+	chr2	242206209	+	.	0	8	1264151_1	23.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1264151_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_2_242231501_242256501_403C;SPAN=2187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:0 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:8 DR:0 LR:-23.11 LO:23.11);ALT=T[chr2:242206209[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242206354	+	chr2	242254523	+	.	9	0	1264154_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1264154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242206354(+)-2:242254523(-)__2_242231501_242256501D;SPAN=48169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=G[chr2:242254523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242255444	+	chr2	242265404	+	.	10	0	1264218_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1264218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242255444(+)-2:242265404(-)__2_242231501_242256501D;SPAN=9960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:0 DR:10 LR:-19.73 LO:22.76);ALT=C[chr2:242265404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242255444	+	chr2	242274539	+	.	9	0	1264219_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1264219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242255444(+)-2:242274539(-)__2_242231501_242256501D;SPAN=19095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=C[chr2:242274539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242265530	+	chr2	242274540	+	.	0	11	1264099_1	11.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=1264099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_242256001_242281001_86C;SPAN=9010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:11 DR:0 LR:-10.84 LO:22.13);ALT=T[chr2:242274540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242506103	+	chr2	242507335	+	ATT	18	18	1264911_1	91.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=ATT;MAPQ=60;MATEID=1264911_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_242501001_242526001_18C;SPAN=1232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:64 GQ:62 PL:[91.7, 0.0, 62.0] SR:18 DR:18 LR:-91.86 LO:91.86);ALT=A[chr2:242507335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242573496	+	chr2	242576354	+	.	0	9	1265175_1	26.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=1265175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_242574501_242599501_248C;SPAN=2858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:6 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:9 DR:0 LR:-26.41 LO:26.41);ALT=T[chr2:242576354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242618066	+	chr2	242619644	+	.	3	7	1265164_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1265164_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_242599001_242624001_337C;SPAN=1578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:7 DR:3 LR:-9.169 LO:19.98);ALT=T[chr2:242619644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242618113	+	chr2	242626068	+	.	8	0	1265165_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1265165_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242618113(+)-2:242626068(-)__2_242599001_242624001D;SPAN=7955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:0 DR:8 LR:-15.84 LO:18.23);ALT=T[chr2:242626068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242619761	+	chr2	242626078	+	.	10	0	1265643_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1265643_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242619761(+)-2:242626078(-)__2_242623501_242648501D;SPAN=6317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:30 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:0 DR:10 LR:-24.88 LO:25.28);ALT=T[chr2:242626078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242641544	+	chr2	242648628	+	.	9	0	1265711_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1265711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:242641544(+)-2:242648628(-)__2_242623501_242648501D;SPAN=7084;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:6 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=C[chr2:242648628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
