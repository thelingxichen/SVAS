chr10	66398774	+	chr10	66400745	+	.	59	49	6319295_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GATA;MAPQ=60;MATEID=6319295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_66395001_66420001_220C;SPAN=1971;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:78 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:49 DR:59 LR:-260.8 LO:260.8);ALT=A[chr10:66400745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	67306934	+	chr10	67315295	+	.	0	49	6322154_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6322154_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_67301501_67326501_35C;SPAN=8361;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:66 GQ:15.2 PL:[143.9, 0.0, 15.2] SR:49 DR:0 LR:-149.8 LO:149.8);ALT=T[chr10:67315295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
