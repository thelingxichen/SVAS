chr5	172261438	+	chr5	172315700	+	.	6	4	2644850_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2644850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_172308501_172333501_70C;SPAN=54262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:4 DR:6 LR:-17.2 LO:18.78);ALT=T[chr5:172315700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172261466	+	chr5	172324003	+	.	12	0	2644851_1	32.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2644851_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:172261466(+)-5:172324003(-)__5_172308501_172333501D;SPAN=62537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:26 GQ:29.3 PL:[32.6, 0.0, 29.3] SR:0 DR:12 LR:-32.57 LO:32.57);ALT=G[chr5:172324003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172336764	+	chr5	172341717	+	.	0	7	2644914_1	6.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2644914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_172333001_172358001_226C;SPAN=4953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:60 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:7 DR:0 LR:-6.852 LO:14.07);ALT=T[chr5:172341717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172410932	+	chr5	172447240	+	.	73	0	2645216_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2645216_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:172410932(+)-5:172447240(-)__5_172406501_172431501D;SPAN=36308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:65 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:0 DR:73 LR:-214.6 LO:214.6);ALT=G[chr5:172447240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172410967	+	chr5	172461400	+	AGTTATCATTACCATGTTGGTGACCTGTTCAGTTTGCTGCTATCTCTTTTGGCTGATTGCAATTCTGGCCCAACTCAACCCTCTCTTTGGACCGCAATTGAAAAATGAAACCATCTGGTATCTGAAGTATCATTGGCCTTGAGGAAGAAGACATGCTCTACAGTGCTCAGTCTTTG	0	157	2645218_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=AGTTATCATTACCATGTTGGTGACCTGTTCAGTTTGCTGCTATCTCTTTTGGCTGATTGCAATTCTGGCCCAACTCAACCCTCTCTTTGGACCGCAATTGAAAAATGAAACCATCTGGTATCTGAAGTATCATTGGCCTTGAGGAAGAAGACATGCTCTACAGTGCTCAGTCTTTG;MAPQ=60;MATEID=2645218_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_172406501_172431501_324C;SPAN=50433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:157 DP:55 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:157 DR:0 LR:-465.4 LO:465.4);ALT=G[chr5:172461400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172447372	+	chr5	172461400	+	.	0	35	2645260_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=2645260_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_172406501_172431501_324C;SPAN=14028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:0 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:35 DR:0 LR:-102.3 LO:102.3);ALT=T[chr5:172461400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172483491	+	chr5	172507583	+	.	10	0	2645314_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2645314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:172483491(+)-5:172507583(-)__5_172504501_172529501D;SPAN=24092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:24 GQ:26.6 PL:[26.6, 0.0, 29.9] SR:0 DR:10 LR:-26.51 LO:26.53);ALT=C[chr5:172507583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
