chr2	148730398	+	chr2	148733469	+	TTGTATTGTACTTGCACTCCAAATAGGTTACTATGTGGACTCTGACGACAAAATCTTTCACGTAAAATTCTTTGT	0	17	1035850_1	39.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=TTGTATTGTACTTGCACTCCAAATAGGTTACTATGTGGACTCTGACGACAAAATCTTTCACGTAAAATTCTTTGT;MAPQ=60;MATEID=1035850_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_148715001_148740001_204C;SPAN=3071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:61 GQ:39.8 PL:[39.8, 0.0, 105.8] SR:17 DR:0 LR:-39.59 LO:41.37);ALT=T[chr2:148733469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	148731124	+	chr2	148778200	+	.	9	0	1035982_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1035982_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:148731124(+)-2:148778200(-)__2_148764001_148789001D;SPAN=47076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=A[chr2:148778200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
