chr6	142468493	+	chr6	142487364	+	.	8	0	3053959_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3053959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:142468493(+)-6:142487364(-)__6_142467501_142492501D;SPAN=18871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=G[chr6:142487364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	142487459	+	chr6	142490687	+	.	0	9	3054002_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3054002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_142467501_142492501_248C;SPAN=3228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:9 DR:0 LR:-11.83 LO:18.75);ALT=T[chr6:142490687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
