chr20	14962958	+	chr20	15013948	+	.	25	22	6933411_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=60;MATEID=6933411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_14945001_14970001_52C;SPAN=50990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:46 GQ:2.4 PL:[115.5, 2.4, 0.0] SR:22 DR:25 LR:-120.3 LO:120.3);ALT=C[chr20:15013948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	14988825	+	chr20	15108818	+	.	7	3	6933921_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6933921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_15092001_15117001_95C;SPAN=119993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:3 DR:7 LR:-15.03 LO:17.94);ALT=T[chr20:15108818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	15000624	+	chr20	15013842	+	.	25	31	6933271_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=6933271_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_14994001_15019001_138C;SPAN=13218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:58 GQ:23.9 PL:[116.3, 0.0, 23.9] SR:31 DR:25 LR:-119.7 LO:119.7);ALT=T[chr20:15013842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	15301734	+	chr20	15303769	+	.	65	37	6934409_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=6934409_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_15288001_15313001_338C;SPAN=2035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:76 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:37 DR:65 LR:-241.0 LO:241.0);ALT=T[chr20:15303769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
