chr3	83853128	+	chr3	83855350	+	.	107	49	2147295_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TATATGGCCTTTT;MAPQ=60;MATEID=2147295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_83839001_83864001_69C;SPAN=2222;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:127 DP:35 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:49 DR:107 LR:-376.3 LO:376.3);ALT=T[chr3:83855350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	84104942	+	chr3	84107385	+	.	0	61	2148035_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2148035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_84084001_84109001_252C;SPAN=2443;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:61 DP:82 GQ:17.6 PL:[179.3, 0.0, 17.6] SR:61 DR:0 LR:-186.6 LO:186.6);ALT=C[chr3:84107385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
