chr1	214656364	-	chr5	115238579	+	.	11	0	810830_1	4.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=810830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:214656364(-)-5:115238579(-)__1_214644501_214669501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:118 GQ:4.4 PL:[4.4, 0.0, 281.6] SR:0 DR:11 LR:-4.342 LO:20.98);ALT=[chr5:115238579[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	214656709	+	chr5	115177778	-	.	35	0	810835_1	87.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=810835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:214656709(+)-5:115177778(+)__1_214644501_214669501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:105 GQ:87.2 PL:[87.2, 0.0, 166.4] SR:0 DR:35 LR:-87.09 LO:88.49);ALT=A]chr5:115177778];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	215492421	+	chr1	215500995	+	CT	0	56	814247_1	99.0	.	EVDNC=ASSMB;INSERTION=CT;MAPQ=60;MATEID=814247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_215477501_215502501_60C;SPAN=8574;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:92 GQ:61.1 PL:[160.1, 0.0, 61.1] SR:56 DR:0 LR:-162.2 LO:162.2);ALT=A[chr1:215500995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	216185316	+	chr1	230741092	+	.	0	21	817039_1	61.0	.	EVDNC=ASSMB;HOMSEQ=CCTGATCACGCTTGATTT;MAPQ=56;MATEID=817039_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_216163501_216188501_138C;SPAN=14555776;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:29 GQ:8.6 PL:[61.4, 0.0, 8.6] SR:21 DR:0 LR:-63.72 LO:63.72);ALT=T[chr1:230741092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	216689969	-	chr3	68048436	+	.	2	58	2084865_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGTGTGTGTGTGTGTATGTGTGTGT;MAPQ=60;MATEID=2084865_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_68036501_68061501_117C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:48 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:58 DR:2 LR:-171.6 LO:171.6);ALT=[chr3:68048436[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	67493708	+	chr3	67496800	+	.	120	73	2083151_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAATTAGATCTC;MAPQ=60;MATEID=2083151_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_67473001_67498001_32C;SPAN=3092;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:165 DP:31 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:73 DR:120 LR:-488.5 LO:488.5);ALT=C[chr3:67496800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	68634773	+	chr3	68640254	+	.	0	110	2087288_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACT;MAPQ=55;MATEID=2087288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_68624501_68649501_85C;SPAN=5481;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:110 DP:45 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:110 DR:0 LR:-326.8 LO:326.8);ALT=T[chr3:68640254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	68739682	+	chr3	68747864	+	TTAAA	148	45	2087698_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TTAAA;MAPQ=60;MATEID=2087698_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_68747001_68772001_52C;SPAN=8182;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:168 DP:19 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:45 DR:148 LR:-498.4 LO:498.4);ALT=A[chr3:68747864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	114756515	+	chr5	114757890	+	.	63	36	3697881_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTATCTCTTGTTTTCTT;MAPQ=60;MATEID=3697881_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_114733501_114758501_194C;SPAN=1375;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:67 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:36 DR:63 LR:-250.9 LO:250.9);ALT=T[chr5:114757890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115177803	+	chr5	115205713	+	.	9	0	3696745_1	14.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3696745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115177803(+)-5:115205713(-)__5_115174501_115199501D;SPAN=27910;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:0 DR:9 LR:-14.54 LO:19.45);ALT=C[chr5:115205713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115205836	+	chr5	115249055	+	.	15	0	3697039_1	23.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=3697039_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115205836(+)-5:115249055(-)__5_115248001_115273001D;SPAN=43219;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:95 GQ:23.9 PL:[23.9, 0.0, 205.4] SR:0 DR:15 LR:-23.78 LO:32.28);ALT=A[chr5:115249055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115205838	+	chr5	115238578	+	.	9	0	3696933_1	10.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3696933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115205838(+)-5:115238578(-)__5_115223501_115248501D;SPAN=32740;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:70 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:0 DR:9 LR:-10.74 LO:18.5);ALT=T[chr5:115238578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115238690	+	chr5	115249057	+	.	28	55	3697040_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=0;MATEID=3697040_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_115248001_115273001_15C;SPAN=10367;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:72 DP:99 GQ:29.3 PL:[210.8, 0.0, 29.3] SR:55 DR:28 LR:-218.7 LO:218.7);ALT=G[chr5:115249057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
