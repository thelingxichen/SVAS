chr5	85913966	+	chr5	85915167	+	.	44	0	2521751_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2521751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:85913966(+)-5:85915167(-)__5_85897001_85922001D;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:87 GQ:88.7 PL:[121.7, 0.0, 88.7] SR:0 DR:44 LR:-121.9 LO:121.9);ALT=C[chr5:85915167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	86704003	+	chr5	86705106	+	.	0	5	2522785_1	3.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2522785_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_86681001_86706001_99C;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:48 GQ:3.5 PL:[3.5, 0.0, 112.4] SR:5 DR:0 LR:-3.501 LO:9.789);ALT=C[chr5:86705106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	86707166	+	chr5	86708493	+	.	0	28	2522794_1	75.0	.	EVDNC=ASSMB;HOMSEQ=ACCTT;MAPQ=60;MATEID=2522794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_86705501_86730501_189C;SPAN=1327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:63 GQ:75.5 PL:[75.5, 0.0, 75.5] SR:28 DR:0 LR:-75.36 LO:75.36);ALT=T[chr5:86708493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
