chr4	32071051	+	chr4	32065770	+	.	13	27	1934299_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GACT;MAPQ=60;MATEID=1934299_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_4_32070501_32095501_116C;SPAN=5281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:30 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:27 DR:13 LR:-102.3 LO:102.3);ALT=]chr4:32071051]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	32065877	+	chr4	32071042	+	AAATATGTGTCGGTTGTTCAAGAGGGATCCAAAAAATCAGAAATCTTTAGTAACTTCCTCAATGTTATACAGCTGTTATGAAGGACAGGATTT	9	37	1934300_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GACT;INSERTION=AAATATGTGTCGGTTGTTCAAGAGGGATCCAAAAAATCAGAAATCTTTAGTAACTTCCTCAATGTTATACAGCTGTTATGAAGGACAGGATTT;MAPQ=60;MATEID=1934300_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_32070501_32095501_116C;SPAN=5165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:32 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:37 DR:9 LR:-118.8 LO:118.8);ALT=G[chr4:32071042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
