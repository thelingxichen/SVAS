chr20	39906375	+	chr20	39907485	+	.	71	9	10540531_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=TCACTGCAAGCTCCGCCTCCCGGGTTCATGCCATTCTCCTGCCTCAGCCTCCTGAGTAGCTGGGACTACAGG;MAPQ=60;MATEID=10540531_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_20_39886001_39911001_274C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:80 DP:169 GQ:99 PL:[218.3, 0.0, 191.9] SR:9 DR:71 LR:-218.4 LO:218.4);ALT=G[chr20:39907485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	39966366	-	chr20	39967675	+	.	4	2	10540775_1	0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=AGACCAGCCTGGC;MAPQ=60;MATEID=10540775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_39959501_39984501_267C;SPAN=1309;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:196 GQ:36.4 PL:[0.0, 36.4, 547.9] SR:2 DR:4 LR:36.6 LO:6.663);ALT=[chr20:39967675[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
