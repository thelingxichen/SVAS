chr15	62706095	+	chr15	62707793	+	.	0	151	8924288_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ATT;MAPQ=60;MATEID=8924288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_62695501_62720501_246C;SPAN=1698;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:151 DP:54 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:151 DR:0 LR:-445.6 LO:445.6);ALT=T[chr15:62707793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
