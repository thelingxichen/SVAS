chr8	40774633	+	chr8	40779779	+	.	59	50	5452344_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=CTCCTGACCTC;MAPQ=60;MATEID=5452344_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_40768001_40793001_191C;SPAN=5146;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:28 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:50 DR:59 LR:-307.0 LO:307.0);ALT=C[chr8:40779779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
