chr19	40615690	+	chr2	65138905	+	C	50	79	10295986_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=10295986_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_40596501_40621501_63C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:39 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:79 DR:50 LR:-293.8 LO:293.8);ALT=]chr19:40615690]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	111096356	-	chr4	111097434	+	.	8	0	2839070_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2839070_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:111096356(-)-4:111097434(-)__4_111083001_111108001D;SPAN=1078;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.374 LO:14.01);ALT=[chr4:111097434[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	111260224	-	chr19	42476957	+	AGGAAGGGAGGAAGGAAAAGGAAGGAAGGGGAAGGAA	3	77	2839815_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;INSERTION=AGGAAGGGAGGAAGGAAAAGGAAGGAAGGGGAAGGAA;MAPQ=60;MATEID=2839815_2;MATENM=0;NM=8;NUMPARTS=2;SCTG=c_4_111254501_111279501_363C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:54 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:77 DR:3 LR:-227.8 LO:227.8);ALT=[chr19:42476957[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	112091058	-	chrX	64833129	+	.	10	0	11206442_1	12.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=11206442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:112091058(-)-23:64833129(-)__23_64827001_64852001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:77 GQ:12.2 PL:[12.2, 0.0, 173.9] SR:0 DR:10 LR:-12.15 LO:20.6);ALT=[chrX:64833129[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	112816051	+	chr4	112258305	+	.	52	0	2844328_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2844328_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:112258305(-)-4:112816051(+)__4_112234501_112259501D;SPAN=557746;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:84 GQ:53.3 PL:[149.0, 0.0, 53.3] SR:0 DR:52 LR:-151.3 LO:151.3);ALT=]chr4:112816051]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	113088079	+	chr4	113471130	+	.	10	0	2848226_1	11.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2848226_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:113088079(+)-4:113471130(-)__4_113459501_113484501D;SPAN=383051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:79 GQ:11.6 PL:[11.6, 0.0, 179.9] SR:0 DR:10 LR:-11.61 LO:20.48);ALT=G[chr4:113471130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	113397103	+	chr4	113498208	-	TA	0	137	2848914_1	99.0	.	EVDNC=ASSMB;INSERTION=TA;MAPQ=60;MATEID=2848914_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_113484001_113509001_375C;SPAN=101105;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:137 DP:25 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:137 DR:0 LR:-406.0 LO:406.0);ALT=T]chr4:113498208];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	40613104	+	chr19	40615761	+	.	45	44	10296040_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAATTAATAGTTTT;MAPQ=60;MATEID=10296040_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40596501_40621501_360C;SPAN=2657;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:91 GQ:14.4 PL:[247.5, 14.4, 0.0] SR:44 DR:45 LR:-250.7 LO:250.7);ALT=T[chr19:40615761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40623096	+	chr19	40625303	+	.	81	33	10295892_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAAAAAAA;MAPQ=48;MATEID=10295892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40621001_40646001_214C;SPAN=2207;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:98 DP:148 GQ:75.5 PL:[283.4, 0.0, 75.5] SR:33 DR:81 LR:-290.1 LO:290.1);ALT=A[chr19:40625303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41349446	-	chr19	41602066	+	.	10	13	10301608_1	34.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAGAGTAGTAATAATAGCAGCTCTTATTTCCTGA;MAPQ=60;MATEID=10301608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41601001_41626001_152C;SPAN=252620;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:92 GQ:34.7 PL:[34.7, 0.0, 186.5] SR:13 DR:10 LR:-34.49 LO:40.6);ALT=[chr19:41602066[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	41521351	+	chr19	41454002	+	.	12	0	10300726_1	19.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=10300726_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41454002(-)-19:41521351(+)__19_41503001_41528001D;SPAN=67349;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:0 DR:12 LR:-19.29 LO:25.9);ALT=]chr19:41521351]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	41852649	-	chr19	41853692	+	.	10	0	10302916_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=10302916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41852649(-)-19:41853692(-)__19_41846001_41871001D;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:120 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.4991 LO:18.56);ALT=[chr19:41853692[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	43244002	+	chr19	43690010	+	.	3	88	10312203_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=CCTCTTACCAATTC;MAPQ=60;MATEID=10312203_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_19_43683501_43708501_320C;SPAN=446008;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:18 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:88 DR:3 LR:-267.4 LO:267.4);ALT=C[chr19:43690010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	43286563	-	chr19	43541073	+	.	2	8	10311312_1	5.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=ATGTCCTAGTGTTTTATGTGTTACCTCTTTTT;MAPQ=35;MATEID=10311312_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_43536501_43561501_564C;SPAN=254510;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:91 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:8 DR:2 LR:-5.055 LO:17.41);ALT=[chr19:43541073[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	43383213	+	chr19	43690010	+	.	20	26	10310430_1	98.0	.	DISC_MAPQ=8;EVDNC=ASDIS;HOMSEQ=CCTCTTACCAATTCCGGT;MAPQ=33;MATEID=10310430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_43365001_43390001_142C;SPAN=306797;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:86 GQ:98.9 PL:[98.9, 0.0, 108.8] SR:26 DR:20 LR:-98.84 LO:98.87);ALT=T[chr19:43690010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	43690648	+	chr19	43422017	+	.	26	0	10312230_1	74.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=10312230_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:43422017(-)-19:43690648(+)__19_43683501_43708501D;SPAN=268631;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:40 GQ:22.1 PL:[74.9, 0.0, 22.1] SR:0 DR:26 LR:-76.59 LO:76.59);ALT=]chr19:43690648]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	43792337	+	chr19	43730605	+	.	10	0	10312693_1	18.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=10312693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:43730605(-)-19:43792337(+)__19_43781501_43806501D;SPAN=61732;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:0 DR:10 LR:-18.11 LO:22.2);ALT=]chr19:43792337]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	43730752	+	chr19	43792744	+	.	8	0	10312694_1	10.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=10312694_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:43730752(+)-19:43792744(-)__19_43781501_43806501D;SPAN=61992;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=C[chr19:43792744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	149032062	+	chr19	43993142	+	.	22	42	11421780_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=GGGTTTCACCATATTGGCCAGGCTGGTCTCAAATTCCTGACTTCAAGTGATC;MAPQ=44;MATEID=11421780_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_23_149009001_149034001_83C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:6 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:42 DR:22 LR:-184.8 LO:184.8);ALT=]chrX:149032062]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chrX	64607618	-	chrX	67824158	+	.	18	0	11217308_1	43.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=11217308_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:64607618(-)-23:67824158(-)__23_67816001_67841001D;SPAN=3216540;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:61 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:0 DR:18 LR:-42.89 LO:44.34);ALT=[chrX:67824158[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	64607772	+	chrX	67823978	-	.	13	0	11217309_1	28.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=11217309_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:64607772(+)-23:67823978(+)__23_67816001_67841001D;SPAN=3216206;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:0 DR:13 LR:-28.55 LO:30.78);ALT=A]chrX:67823978];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	64641775	+	chrX	64642898	-	.	4	2	11204731_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCTCACTGCAAGCTCC;MAPQ=60;MATEID=11204731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_64631001_64656001_333C;SPAN=1123;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:167 GQ:28.6 PL:[0.0, 28.6, 462.1] SR:2 DR:4 LR:28.74 LO:7.011);ALT=C]chrX:64642898];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	67798572	-	chrX	67825758	+	.	24	0	11217620_1	59.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=11217620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:67798572(-)-23:67825758(-)__23_67791501_67816501D;SPAN=27186;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:73 GQ:59.6 PL:[59.6, 0.0, 115.7] SR:0 DR:24 LR:-59.45 LO:60.5);ALT=[chrX:67825758[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
