chr1	9121445	+	chr14	93713179	-	.	139	55	8686331_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=59;MATEID=8686331_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_93712501_93737501_44C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:167 DP:83 GQ:45.1 PL:[495.1, 45.1, 0.0] SR:55 DR:139 LR:-495.1 LO:495.1);ALT=T]chr14:93713179];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	9121449	-	chr14	93712482	+	.	99	31	8685884_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGGG;MAPQ=60;MATEID=8685884_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_93688001_93713001_419C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:121 DP:122 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:31 DR:99 LR:-359.8 LO:359.8);ALT=[chr14:93712482[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	9595642	+	chr1	9597667	+	.	27	44	49120_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TGCCACTGCACTCCAGCCTGGGTGACAGAG;MAPQ=9;MATEID=49120_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_9579501_9604501_458C;SPAN=2025;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:86 GQ:26.3 PL:[181.4, 0.0, 26.3] SR:44 DR:27 LR:-187.9 LO:187.9);ALT=G[chr1:9597667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111896187	+	chr10	102036213	+	.	17	32	6478712_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6478712_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_102018001_102043001_480C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:45 DP:40 GQ:12 PL:[132.0, 12.0, 0.0] SR:32 DR:17 LR:-132.0 LO:132.0);ALT=C[chr10:102036213[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	112691792	+	chr1	112704704	+	.	73	50	458468_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=458468_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_1_112675501_112700501_26C;SPAN=12912;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:7 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:50 DR:73 LR:-293.8 LO:293.8);ALT=G[chr1:112704704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112835105	+	chr1	112837666	+	.	34	45	458862_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=AAAAGAGGACACAAACAA;MAPQ=60;MATEID=458862_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_112822501_112847501_253C;SPAN=2561;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:21 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:45 DR:34 LR:-221.2 LO:221.2);ALT=A[chr1:112837666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113716653	+	chr1	113507412	+	.	0	56	461272_1	99.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=461272_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_113704501_113729501_289C;SPAN=209241;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:56 DP:46 GQ:15 PL:[165.0, 15.0, 0.0] SR:56 DR:0 LR:-165.0 LO:165.0);ALT=]chr1:113716653]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	113611339	+	chr1	113613778	+	.	132	71	461020_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAACACATATTTGCG;MAPQ=60;MATEID=461020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_113606501_113631501_224C;SPAN=2439;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:178 DP:39 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:71 DR:132 LR:-528.1 LO:528.1);ALT=G[chr1:113613778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102074838	+	chr2	2824194	+	.	10	0	897129_1	27.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=897129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:2824194(-)-10:102074838(+)__2_2817501_2842501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:19 GQ:17.9 PL:[27.8, 0.0, 17.9] SR:0 DR:10 LR:-27.97 LO:27.97);ALT=]chr10:102074838]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	97320864	+	chr12	130794392	+	.	18	0	1186982_1	42.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1186982_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97320864(+)-12:130794392(-)__2_97314001_97339001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:63 GQ:42.5 PL:[42.5, 0.0, 108.5] SR:0 DR:18 LR:-42.35 LO:44.03);ALT=A[chr12:130794392[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	97854268	+	chr2	97856173	+	.	8	0	1190946_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1190946_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97854268(+)-2:97856173(-)__2_97853001_97878001D;SPAN=1905;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:115 GQ:4.5 PL:[0.0, 4.5, 287.1] SR:0 DR:8 LR:4.748 LO:14.2);ALT=A[chr2:97856173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	98559528	-	chr5	176585252	+	.	12	0	1194533_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1194533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:98559528(-)-5:176585252(-)__2_98539001_98564001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=[chr5:176585252[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	98664284	+	chrX	35566369	-	.	6	32	11070347_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=AGGAAAGGAAAGGAAAGGAAAGGAAAGGAAAGGAAAGG;MAPQ=59;MATEID=11070347_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_23_35549501_35574501_167C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:53 GQ:18.8 PL:[107.9, 0.0, 18.8] SR:32 DR:6 LR:-111.1 LO:111.1);ALT=T]chrX:35566369];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	99113005	-	chr2	99114182	+	.	11	3	1196761_1	7.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGCTTCTGCACAGCAAAG;MAPQ=60;MATEID=1196761_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_99102501_99127501_170C;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:130 GQ:7.7 PL:[7.7, 0.0, 308.0] SR:3 DR:11 LR:-7.693 LO:25.21);ALT=[chr2:99114182[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	132850328	+	chr21	14480725	+	.	2	4	1351428_1	17.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=ATAAATATATTATACCAATATTTA;MAPQ=60;MATEID=1351428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_132839001_132864001_359C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:6 DP:8 GQ:1.1 PL:[17.6, 0.0, 1.1] SR:4 DR:2 LR:-18.4 LO:18.4);ALT=A[chr21:14480725[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	133429898	+	chr2	133431213	+	.	0	44	1354352_1	99.0	.	EVDNC=ASSMB;HOMSEQ=T;MAPQ=60;MATEID=1354352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_133427001_133452001_173C;SPAN=1315;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:70 GQ:43.7 PL:[126.2, 0.0, 43.7] SR:44 DR:0 LR:-128.5 LO:128.5);ALT=T[chr2:133431213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	133690699	+	chr2	133863715	-	.	9	30	1356529_1	99.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=TTTTTGTATTTTTAGTAGAGATGGGGTTTCACC;MAPQ=60;MATEID=1356529_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_133843501_133868501_127C;SPAN=173016;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:46 GQ:5.7 PL:[122.1, 5.7, 0.0] SR:30 DR:9 LR:-124.8 LO:124.8);ALT=C]chr2:133863715];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	133717772	+	chr17	1547322	-	.	30	38	9466527_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=9466527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_1543501_1568501_120C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:55 DP:31 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:38 DR:30 LR:-161.7 LO:161.7);ALT=T]chr17:1547322];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	133776695	-	chrX	35939541	+	.	51	36	11071725_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=11071725_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_35917001_35942001_206C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:67 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:36 DR:51 LR:-224.5 LO:224.5);ALT=[chrX:35939541[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	133784339	-	chrX	36143221	+	.	6	3	11072845_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=11072845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_36137501_36162501_357C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:81 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:3 DR:6 LR:-4.463 LO:15.47);ALT=[chrX:36143221[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	134568710	+	chr2	134566522	+	.	14	0	1358530_1	11.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1358530_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:134566522(-)-2:134568710(+)__2_134554001_134579001D;SPAN=2188;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:127 GQ:11.9 PL:[11.9, 0.0, 295.7] SR:0 DR:14 LR:-11.81 LO:27.77);ALT=]chr2:134568710]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	134966717	+	chr2	134970131	+	.	108	45	1360402_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAACTGGCTTATTTTT;MAPQ=60;MATEID=1360402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_134946001_134971001_341C;SPAN=3414;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:150 DP:687 GQ:99 PL:[309.2, 0.0, 1359.0] SR:45 DR:108 LR:-309.0 LO:346.4);ALT=T[chr2:134970131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	72285074	+	chr7	39209628	-	.	8	0	2102779_1	7.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2102779_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:72285074(+)-7:39209628(+)__3_72275001_72300001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:0 DR:8 LR:-6.901 LO:15.9);ALT=A]chr7:39209628];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	118073384	+	chr5	176753871	-	.	8	21	3955893_1	63.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TCTTTCTTTCTTTCTTTCTTTCTTTCTTTCTTTC;MAPQ=60;MATEID=3955893_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_5_176743001_176768001_337C;SPAN=58680487;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:47 GQ:50 PL:[63.2, 0.0, 50.0] SR:21 DR:8 LR:-63.26 LO:63.26);ALT=C]chr5:176753871];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	118459444	-	chr7	38582435	+	.	4	18	4719064_1	38.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=40;MATEID=4719064_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_38563001_38588001_131C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:102 GQ:38.6 PL:[38.6, 0.0, 206.9] SR:18 DR:4 LR:-38.39 LO:45.13);ALT=[chr7:38582435[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	119380146	+	chr5	119382681	+	GAG	137	84	3713139_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GAG;MAPQ=60;MATEID=3713139_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_5_119364001_119389001_81C;SPAN=2535;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:183 DP:36 GQ:49.3 PL:[541.3, 49.3, 0.0] SR:84 DR:137 LR:-541.3 LO:541.3);ALT=T[chr5:119382681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9873710	+	chr5	119855963	+	.	20	15	3715050_1	93.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GCCTGTAATCCCAGCTGCTCAAGAGGCTGAGGCAGGAGAATC;MAPQ=11;MATEID=3715050_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_5_119854001_119879001_376C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:68 GQ:70.7 PL:[93.8, 0.0, 70.7] SR:15 DR:20 LR:-93.97 LO:93.97);ALT=]chr18:9873710]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	175720563	+	chr5	175721733	-	.	8	0	3950772_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=3950772_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:175720563(+)-5:175721733(+)__5_175714001_175739001D;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:167 GQ:18.7 PL:[0.0, 18.7, 442.3] SR:0 DR:8 LR:18.84 LO:12.87);ALT=A]chr5:175721733];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	175733390	+	chr18	55381820	-	.	19	38	3950848_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3950848_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_175714001_175739001_179C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:49 DP:44 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:38 DR:19 LR:-145.2 LO:145.2);ALT=C]chr18:55381820];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	176387587	+	chr5	176390181	+	.	62	32	3953761_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAAAA;MAPQ=60;MATEID=3953761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176375501_176400501_241C;SPAN=2594;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:77 DP:246 GQ:99 PL:[187.6, 0.0, 408.8] SR:32 DR:62 LR:-187.5 LO:192.1);ALT=A[chr5:176390181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38297779	+	chr7	38317403	+	.	18	0	4717771_1	12.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4717771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:38297779(+)-7:38317403(-)__7_38293501_38318501D;SPAN=19624;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:173 GQ:12.7 PL:[12.7, 0.0, 405.5] SR:0 DR:18 LR:-12.55 LO:35.23);ALT=A[chr7:38317403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	40124984	+	chr7	40485684	+	.	77	26	4730310_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AGGAA;MAPQ=60;MATEID=4730310_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_40106501_40131501_239C;SPAN=360700;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:51 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:26 DR:77 LR:-274.0 LO:274.0);ALT=A[chr7:40485684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	40782042	+	chr7	41038527	+	.	65	36	4734455_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=4734455_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_41037501_41062501_63C;SPAN=256485;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:67 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:36 DR:65 LR:-250.9 LO:250.9);ALT=A[chr7:41038527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	40879376	-	chr7	40880470	+	.	115	94	4733800_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4733800_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_7_40866001_40891001_122C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:185 DP:80 GQ:49.9 PL:[547.9, 49.9, 0.0] SR:94 DR:115 LR:-547.9 LO:547.9);ALT=[chr7:40880470[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	41856778	+	chr7	41876279	+	.	18	0	4739015_1	52.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4739015_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:41856778(+)-7:41876279(-)__7_41870501_41895501D;SPAN=19501;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:18 DP:14 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=C[chr7:41876279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11098997	-	chr18	22222390	+	.	19	33	5391187_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=ACTACTGATAA;MAPQ=60;MATEID=5391187_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_11098501_11123501_2C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:46 DP:8 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:33 DR:19 LR:-135.3 LO:135.3);ALT=[chr18:22222390[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	11893345	+	chr8	11788240	+	.	32	0	5392857_1	92.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=5392857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:11788240(-)-8:11893345(+)__8_11784501_11809501D;SPAN=105105;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:32 DP:8 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=]chr8:11893345]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	12233486	+	chr8	12236124	+	.	47	12	5394903_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=TGTGTGTGTGTGTGTGTGT;MAPQ=52;MATEID=5394903_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_12225501_12250501_50C;SPAN=2638;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:109 GQ:99 PL:[145.4, 0.0, 119.0] SR:12 DR:47 LR:-145.6 LO:145.6);ALT=T[chr8:12236124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	101384912	+	chr18	24804845	+	AGTGTTACAGC	24	79	6474935_1	99.0	.	DISC_MAPQ=43;EVDNC=TSI_L;INSERTION=AGTGTTACAGC;MAPQ=60;MATEID=6474935_2;MATENM=2;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_10_101381001_101406001_214C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:97 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:79 DR:24 LR:-300.4 LO:300.4);ALT=G[chr18:24804845[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	131144870	+	chr10	102686149	+	TGCTGACATAAAACATCGGGGAGACCTCCAGGAAGCAAGAACACCGCCCATAGCTCTTGGGTTTGGTAAGTGGAATGTAAATATGCCGGAAGGCTGGGCTCAGTGGCTCATGCCTTTAATCCCAACACTTTGGGAGGCCAAGGCCAGTGGATCACTGGAGG	3	76	7915017_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=TGCTGACATAAAACATCGGGGAGACCTCCAGGAAGCAAGAACACCGCCCATAGCTCTTGGGTTTGGTAAGTGGAATGTAAATATGCCGGAAGGCTGGGCTCAGTGGCTCATGCCTTTAATCCCAACACTTTGGGAGGCCAAGGCCAGTGGATCACTGGAGG;MAPQ=60;MATEID=7915017_2;MATENM=6;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_12_131124001_131149001_142C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:49 GQ:21 PL:[231.0, 21.0, 0.0] SR:76 DR:3 LR:-231.1 LO:231.1);ALT=]chr12:131144870]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	103513175	-	chr10	103514547	+	.	3	4	6485153_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=6485153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_103512501_103537501_250C;SPAN=1372;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:114 GQ:10.8 PL:[0.0, 10.8, 297.0] SR:4 DR:3 LR:11.08 LO:9.9);ALT=[chr10:103514547[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	94081927	+	chr10	103623538	+	AATATGGTGAAACCCTGTCTCTACTAAAAATACAAAAATTAGCTGGGTGTGGTGCCATGTGCCTGTAGT	0	18	6486312_1	34.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCCAGCTA;INSERTION=AATATGGTGAAACCCTGTCTCTACTAAAAATACAAAAATTAGCTGGGTGTGGTGCCATGTGCCTGTAGT;MAPQ=60;MATEID=6486312_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_103610501_103635501_234C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:93 GQ:34.4 PL:[34.4, 0.0, 189.5] SR:18 DR:0 LR:-34.22 LO:40.51);ALT=]chr14:94081927]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr18	21903372	+	chr10	104027094	+	.	5	26	6488145_1	67.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=TCTACTAAAAATACAAAAATTAGC;MAPQ=13;MATEID=6488145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_104027001_104052001_468C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:81 GQ:67.4 PL:[67.4, 0.0, 126.8] SR:26 DR:5 LR:-67.18 LO:68.26);ALT=]chr18:21903372]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	131917518	+	chr12	131918759	+	.	18	0	7918237_1	28.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7918237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:131917518(+)-12:131918759(-)__12_131908001_131933001D;SPAN=1241;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:116 GQ:28.1 PL:[28.1, 0.0, 252.5] SR:0 DR:18 LR:-27.99 LO:38.59);ALT=T[chr12:131918759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	723817	+	chr17	724921	+	.	99	0	9463955_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=9463955_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:723817(+)-17:724921(-)__17_710501_735501D;SPAN=1104;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:36 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:0 DR:99 LR:-293.8 LO:293.8);ALT=A[chr17:724921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1625043	-	chr17	1626115	+	.	8	0	9466610_1	11.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=9466610_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1625043(-)-17:1626115(-)__17_1617001_1642001D;SPAN=1072;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=[chr17:1626115[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	10222280	+	chr18	10223605	+	.	0	127	9894043_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AA;MAPQ=60;MATEID=9894043_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_10216501_10241501_97C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:127 DP:43 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:127 DR:0 LR:-376.3 LO:376.3);ALT=A[chr18:10223605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21903372	+	chr18	21904594	+	.	62	49	9936440_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAAATTAGC;MAPQ=60;MATEID=9936440_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21903001_21928001_293C;SPAN=1222;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:115 GQ:21 PL:[320.1, 21.0, 0.0] SR:49 DR:62 LR:-323.4 LO:323.4);ALT=C[chr18:21904594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	14816896	+	chr21	14818166	+	.	58	0	10708023_1	99.0	.	DISC_MAPQ=7;EVDNC=DSCRD;IMPRECISE;MAPQ=7;MATEID=10708023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:14816896(+)-21:14818166(-)__21_14798001_14823001D;SPAN=1270;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:20 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=A[chr21:14818166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	15460416	+	chr21	15461865	+	TTATAAATGATATATAAATCAATAATATATCATTAATAATATATCATATATAATAATTAATATAATTAATAATATAATTAAAATATAATATATAATTATAAATATAATATATAATTATAATTATATTTTTATGTATTTTTAATAATTCATATA	5	36	10710062_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;INSERTION=TTATAAATGATATATAAATCAATAATATATCATTAATAATATATCATATATAATAATTAATATAATTAATAATATAATTAAAATATAATATATAATTATAAATATAATATATAATTATAATTATATTTTTATGTATTTTTAATAATTCATATA;MAPQ=60;MATEID=10710062_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_15459501_15484501_27C;SPAN=1449;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:40 DP:12 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:36 DR:5 LR:-118.8 LO:118.8);ALT=A[chr21:15461865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	15460780	+	chr21	15461865	+	AATAATTCATATA	7	11	10710063_1	38.0	.	DISC_MAPQ=30;EVDNC=TSI_L;INSERTION=AATAATTCATATA;MAPQ=60;MATEID=10710063_2;MATENM=0;NM=5;NUMPARTS=3;REPSEQ=TTTTT;SCTG=c_21_15459501_15484501_27C;SPAN=1085;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:10 GQ:3.9 PL:[38.9, 3.9, 0.0] SR:11 DR:7 LR:-38.99 LO:38.99);ALT=T[chr21:15461865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
