chr3	85396173	+	chr3	85397188	-	.	2	3	2152725_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAGGAGTTCAAG;MAPQ=60;MATEID=2152725_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_85382501_85407501_102C;SPAN=1015;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:141 GQ:24.6 PL:[0.0, 24.6, 389.4] SR:3 DR:2 LR:25.0 LO:5.515);ALT=G]chr3:85397188];VARTYPE=BND:INV-hh;JOINTYPE=hh
