chr10	28214513	-	chr10	28215800	+	.	3	2	6161755_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGCCAG;MAPQ=0;MATEID=6161755_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_10_28199501_28224501_289C;SECONDARY;SPAN=1287;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:142 GQ:24.9 PL:[0.0, 24.9, 392.7] SR:2 DR:3 LR:25.27 LO:5.502);ALT=[chr10:28215800[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
