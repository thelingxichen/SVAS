chr15	22373079	+	chr15	22383653	+	.	59	44	5894402_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=5894402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_22368501_22393501_393C;SPAN=10574;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:80 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:44 DR:59 LR:-250.9 LO:250.9);ALT=T[chr15:22383653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
