chr1	25158703	+	chr1	25161510	+	.	83	65	132183_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTGATTTTTTATTTTT;MAPQ=60;MATEID=132183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25161501_25186501_315C;SPAN=2807;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:12 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:65 DR:83 LR:-333.4 LO:333.4);ALT=T[chr1:25161510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25186264	-	chr2	22740187	+	.	3	30	933980_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATTTATTTATTTATTTATTTATTTATTTAT;MAPQ=60;MATEID=933980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_22736001_22761001_241C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:33 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:30 DR:3 LR:-102.3 LO:102.3);ALT=[chr2:22740187[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
