chr7	57471578	+	chr7	57496109	+	.	46	50	3328533_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=3328533_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_57477001_57502001_167C;SPAN=24531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:38 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:50 DR:46 LR:-214.6 LO:214.6);ALT=C[chr7:57496109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	57957731	+	chr7	57959391	+	.	95	23	3331055_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGACAGAAGAATTCTGAGAAACTTCTTTGTGAT;MAPQ=60;MATEID=3331055_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_7_57942501_57967501_322C;SPAN=1660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:19 GQ:30 PL:[330.0, 30.0, 0.0] SR:23 DR:95 LR:-330.1 LO:330.1);ALT=T[chr7:57959391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	58008342	+	chr7	58006979	+	.	4	1	3331254_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=A;MAPQ=49;MATEID=3331254_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_57991501_58016501_186C;SPAN=1363;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:89 GQ:10.8 PL:[0.0, 10.8, 237.6] SR:1 DR:4 LR:10.91 LO:6.32);ALT=]chr7:58008342]A;VARTYPE=BND:DUP-th;JOINTYPE=th
