chr5	77947061	-	chr5	77948740	+	.	12	0	3554445_1	1.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=3554445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:77947061(-)-5:77948740(-)__5_77934501_77959501D;SPAN=1679;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:140 GQ:1.7 PL:[1.7, 0.0, 338.3] SR:0 DR:12 LR:-1.683 LO:22.43);ALT=[chr5:77948740[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	78426619	+	chr16	67746178	+	.	21	0	3557691_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3557691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:78426619(+)-16:67746178(-)__5_78424501_78449501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:51 GQ:55.7 PL:[55.7, 0.0, 65.6] SR:0 DR:21 LR:-55.5 LO:55.58);ALT=T[chr16:67746178[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	79074616	+	chr8	92534313	-	.	19	0	5542526_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5542526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:79074616(+)-8:92534313(+)__8_92512001_92537001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:41 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:0 DR:19 LR:-51.62 LO:51.62);ALT=C]chr8:92534313];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	79176062	-	chr5	79178207	+	.	9	0	3560201_1	0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=3560201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:79176062(-)-5:79178207(-)__5_79159501_79184501D;SPAN=2145;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:141 GQ:8.1 PL:[0.0, 8.1, 356.4] SR:0 DR:9 LR:8.491 LO:15.62);ALT=[chr5:79178207[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	66925768	+	chr16	66926920	-	.	9	0	9377995_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9377995_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:66925768(+)-16:66926920(+)__16_66909501_66934501D;SPAN=1152;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:142 GQ:8.4 PL:[0.0, 8.4, 359.7] SR:0 DR:9 LR:8.762 LO:15.59);ALT=C]chr16:66926920];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	68543287	-	chr16	68544574	+	.	12	0	9385537_1	10.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=9385537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:68543287(-)-16:68544574(-)__16_68526501_68551501D;SPAN=1287;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:109 GQ:10.1 PL:[10.1, 0.0, 254.3] SR:0 DR:12 LR:-10.08 LO:23.8);ALT=[chr16:68544574[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
