chr8	93190431	-	chr8	93195305	+	TGTATGTATGTAGAAAAAATCTGTA	10	26	3970858_1	76.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGA;INSERTION=TGTATGTATGTAGAAAAAATCTGTA;MAPQ=60;MATEID=3970858_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_93173501_93198501_230C;SPAN=4874;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:72 GQ:76.4 PL:[76.4, 0.0, 96.2] SR:26 DR:10 LR:-76.22 LO:76.38);ALT=[chr8:93195305[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	93190489	+	chr8	93195166	-	TGTATGTATGTAGAAAAAATCTGTA	5	29	3970859_1	86.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=TGTATGTATGTAGAAAAAATCTGTA;MAPQ=60;MATEID=3970859_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_93173501_93198501_230C;SPAN=4677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:69 GQ:80.3 PL:[86.9, 0.0, 80.3] SR:29 DR:5 LR:-86.95 LO:86.95);ALT=A]chr8:93195166];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	93966816	+	chr8	93978261	+	.	11	0	3972685_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3972685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:93966816(+)-8:93978261(-)__8_93957501_93982501D;SPAN=11445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:0 DR:11 LR:-10.84 LO:22.13);ALT=A[chr8:93978261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
