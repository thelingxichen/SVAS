chr5	56205572	+	chr5	56208836	+	.	7	4	2476980_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=2476980_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_56203001_56228001_218C;SPAN=3264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:4 DR:7 LR:-18.11 LO:22.2);ALT=T[chr5:56208836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	56205572	+	chr5	56209698	+	ACAGTATATCAGAAGTATGAGCCGATCTTTTTCCAGTCCATTGGAAATCCGTTTATTTTTAGATGCCTGGATGGGGTACTCATTGATGGGAATGACAAAGGGATATCAAAAGTTGTGTA	0	10	2476981_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=ACAGTATATCAGAAGTATGAGCCGATCTTTTTCCAGTCCATTGGAAATCCGTTTATTTTTAGATGCCTGGATGGGGTACTCATTGATGGGAATGACAAAGGGATATCAAAAGTTGTGTA;MAPQ=60;MATEID=2476981_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_5_56203001_56228001_218C;SPAN=4126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:10 DR:0 LR:-17.84 LO:22.11);ALT=T[chr5:56209698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	56470040	+	chr5	56471273	+	.	47	13	2477435_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2477435_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_56448001_56473001_206C;SPAN=1233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:44 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:13 DR:47 LR:-151.8 LO:151.8);ALT=T[chr5:56471273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57323478	+	chr5	57333779	+	.	54	43	2478738_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=2478738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_57330001_57355001_95C;SPAN=10301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:11 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:43 DR:54 LR:-241.0 LO:241.0);ALT=C[chr5:57333779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57680001	+	chr5	57686102	+	.	48	21	2479414_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAACAC;MAPQ=60;MATEID=2479414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_57673001_57698001_181C;SPAN=6101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:24 GQ:15 PL:[165.0, 15.0, 0.0] SR:21 DR:48 LR:-165.0 LO:165.0);ALT=C[chr5:57686102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57778087	+	chr5	57776911	+	.	14	0	2479318_1	28.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2479318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:57776911(-)-5:57778087(+)__5_57771001_57796001D;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:66 GQ:28.4 PL:[28.4, 0.0, 130.7] SR:0 DR:14 LR:-28.33 LO:32.13);ALT=]chr5:57778087]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	57787413	+	chr5	57789455	+	.	10	0	2479335_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2479335_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:57787413(+)-5:57789455(-)__5_57771001_57796001D;SPAN=2042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:0 DR:10 LR:-17.03 LO:21.86);ALT=T[chr5:57789455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57787413	+	chr5	57792546	+	.	12	0	2479336_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2479336_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:57787413(+)-5:57792546(-)__5_57771001_57796001D;SPAN=5133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:0 DR:12 LR:-24.71 LO:27.71);ALT=T[chr5:57792546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	57787419	+	chr5	57789971	+	.	18	0	2479337_1	46.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2479337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:57787419(+)-5:57789971(-)__5_57771001_57796001D;SPAN=2552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:47 GQ:46.7 PL:[46.7, 0.0, 66.5] SR:0 DR:18 LR:-46.68 LO:46.89);ALT=A[chr5:57789971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
