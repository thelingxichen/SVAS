chr6	84207449	+	chr6	84610825	-	.	35	0	4308545_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=4308545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:84207449(+)-6:84610825(+)__6_84182001_84207001D;SPAN=403376;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:0 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:35 LR:-102.3 LO:102.3);ALT=T]chr6:84610825];VARTYPE=BND:INV-hh;JOINTYPE=hh
