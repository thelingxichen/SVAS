chr3	41680987	+	chr1	7846059	+	.	31	32	1968874_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=GTAATCCCAGCACTTTGGGAGGCCGAG;MAPQ=20;MATEID=1968874_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_41674501_41699501_353C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:62 GQ:9.9 PL:[168.3, 9.9, 0.0] SR:32 DR:31 LR:-170.1 LO:170.1);ALT=]chr3:41680987]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	7846227	+	chr3	41681110	+	.	25	36	1968876_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;HOMSEQ=TCGGGAGGCTGAGACAGGAGAA;MAPQ=60;MATEID=1968876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_41674501_41699501_1C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:56 DP:52 GQ:15 PL:[165.0, 15.0, 0.0] SR:36 DR:25 LR:-165.0 LO:165.0);ALT=A[chr3:41681110[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
