chr1	725394	+	chr1	724145	+	.	10	0	7818_1	0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=7818_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:724145(-)-1:725394(+)__1_710501_735501D;SPAN=1249;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:224 GQ:27.4 PL:[0.0, 27.4, 597.4] SR:0 DR:10 LR:27.68 LO:15.77);ALT=]chr1:725394]T;VARTYPE=BND:DUP-th;JOINTYPE=th
