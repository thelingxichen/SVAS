chr4	120219935	+	chr4	120221491	+	.	0	95	2173114_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2173114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_120197001_120222001_119C;SPAN=1556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:95 DP:145 GQ:76.4 PL:[274.4, 0.0, 76.4] SR:95 DR:0 LR:-280.4 LO:280.4);ALT=C[chr4:120221491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
