chr5	125498520	+	chr5	125496391	+	.	35	0	2573710_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2573710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:125496391(-)-5:125498520(+)__5_125489001_125514001D;SPAN=2129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:49 GQ:16.4 PL:[102.2, 0.0, 16.4] SR:0 DR:35 LR:-105.8 LO:105.8);ALT=]chr5:125498520]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	125496664	+	chr5	125498727	+	.	20	0	2573711_1	51.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2573711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:125496664(+)-5:125498727(-)__5_125489001_125514001D;SPAN=2063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:53 GQ:51.8 PL:[51.8, 0.0, 74.9] SR:0 DR:20 LR:-51.66 LO:51.93);ALT=T[chr5:125498727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	126065136	+	chr14	20777471	+	G	13	37	5665081_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=5665081_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_14_20776001_20801001_223C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:31 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:37 DR:13 LR:-112.2 LO:112.2);ALT=C[chr14:20777471[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	126146042	+	chr5	126147465	+	.	3	2	2574716_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2574716_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_126126001_126151001_280C;SPAN=1423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:2 DR:3 LR:-1.062 LO:9.396);ALT=A[chr5:126147465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	126156828	+	chr5	126158471	+	.	3	4	2574788_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2574788_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_126150501_126175501_174C;SPAN=1643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:55 GQ:5 PL:[5.0, 0.0, 127.1] SR:4 DR:3 LR:-4.905 LO:11.87);ALT=G[chr5:126158471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	126853449	+	chr5	126859149	+	.	9	0	2575808_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2575808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:126853449(+)-5:126859149(-)__5_126836501_126861501D;SPAN=5700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:60 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.45 LO:19.15);ALT=G[chr5:126859149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	127407443	+	chr5	127410917	+	.	42	21	2576543_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=0;MATEID=2576543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_127400001_127425001_182C;SPAN=3474;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:19 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:21 DR:42 LR:-151.8 LO:151.8);ALT=G[chr5:127410917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	14954406	+	chr12	14956342	+	.	11	0	5104324_1	11.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=5104324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:14954406(+)-12:14956342(-)__12_14945001_14970001D;SPAN=1936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:0 DR:11 LR:-10.84 LO:22.13);ALT=T[chr12:14956342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15095657	+	chr12	15097710	+	.	14	29	5105333_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5105333_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_12_15092001_15117001_201C;SPAN=2053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:107 GQ:99 PL:[109.7, 0.0, 149.3] SR:29 DR:14 LR:-109.7 LO:110.0);ALT=T[chr12:15097710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15095657	+	chr12	15114471	+	TTCACCCCAGTCCTGTAGGTGTGCTGAACGTATTTCAGGCCTGACACAATATCCCTGTTCACTTTGAAGTGAATTTTGACTCTATATTCAGAACCTTCCTTTAACACAATGGTTTCCTTTTTGAGGGCTTCCAGATCTCCAGTAAGGTCCATGGTGATTGGTCCCGGGGCACTCTCACAAACCAGGGTGAGCCGGGTGACAACGACATTGGGGGCTTTCGGATCTGTCACCACAGGACCATCTCCCAGCAGCGTTTTCTTGTACTTAATTAGACTCTCATCATCTTTGTCCATTTCCTGCAGCTCTTTCAGGGACTTCTGTGGTGGAGGCTTATAATTGAGCTTGCTGTCCAGCTCATCATCGTCATCCTCCTCCACATGTGGCTCTGGGGCTTTTTCAGTCATTCTGATCTATTT	9	45	5105334_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TTCACCCCAGTCCTGTAGGTGTGCTGAACGTATTTCAGGCCTGACACAATATCCCTGTTCACTTTGAAGTGAATTTTGACTCTATATTCAGAACCTTCCTTTAACACAATGGTTTCCTTTTTGAGGGCTTCCAGATCTCCAGTAAGGTCCATGGTGATTGGTCCCGGGGCACTCTCACAAACCAGGGTGAGCCGGGTGACAACGACATTGGGGGCTTTCGGATCTGTCACCACAGGACCATCTCCCAGCAGCGTTTTCTTGTACTTAATTAGACTCTCATCATCTTTGTCCATTTCCTGCAGCTCTTTCAGGGACTTCTGTGGTGGAGGCTTATAATTGAGCTTGCTGTCCAGCTCATCATCGTCATCCTCCTCCACATGTGGCTCTGGGGCTTTTTCAGTCATTCTGATCTATTT;MAPQ=60;MATEID=5105334_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_12_15092001_15117001_201C;SPAN=18814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:226 GQ:99 PL:[110.5, 0.0, 437.3] SR:45 DR:9 LR:-110.4 LO:121.5);ALT=T[chr12:15114471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15095673	+	chr12	15102734	+	.	8	0	5105335_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5105335_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15095673(+)-12:15102734(-)__12_15092001_15117001D;SPAN=7061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:0 DR:8 LR:3.123 LO:14.39);ALT=T[chr12:15102734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15095683	+	chr12	15100804	+	.	14	0	5105336_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5105336_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15095683(+)-12:15100804(-)__12_15092001_15117001D;SPAN=5121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:89 GQ:22.1 PL:[22.1, 0.0, 193.7] SR:0 DR:14 LR:-22.1 LO:30.11);ALT=T[chr12:15100804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15097817	+	chr12	15103472	+	.	12	0	5105354_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5105354_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15097817(+)-12:15103472(-)__12_15092001_15117001D;SPAN=5655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:219 GQ:19.6 PL:[0.0, 19.6, 571.0] SR:0 DR:12 LR:19.72 LO:20.01);ALT=T[chr12:15103472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15100884	+	chr12	15102735	+	.	3	96	5105360_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=5105360_2;MATENM=0;NM=0;NUMPARTS=6;REPSEQ=CC;SCTG=c_12_15092001_15117001_201C;SPAN=1851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:98 DP:136 GQ:42.5 PL:[286.7, 0.0, 42.5] SR:96 DR:3 LR:-296.9 LO:296.9);ALT=C[chr12:15102735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15100931	+	chr12	15103464	+	.	28	0	5105361_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5105361_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15100931(+)-12:15103464(-)__12_15092001_15117001D;SPAN=2533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:150 GQ:51.8 PL:[51.8, 0.0, 312.5] SR:0 DR:28 LR:-51.79 LO:62.52);ALT=A[chr12:15103464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15100932	+	chr12	15114469	+	.	29	0	5105362_1	46.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5105362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15100932(+)-12:15114469(-)__12_15092001_15117001D;SPAN=13537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:184 GQ:46 PL:[46.0, 0.0, 399.2] SR:0 DR:29 LR:-45.88 LO:62.39);ALT=A[chr12:15114469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15102871	+	chr12	15114469	+	.	109	0	5105367_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5105367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:15102871(+)-12:15114469(-)__12_15092001_15117001D;SPAN=11598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:109 DP:186 GQ:99 PL:[309.5, 0.0, 141.2] SR:0 DR:109 LR:-312.8 LO:312.8);ALT=G[chr12:15114469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	15103658	+	chr12	15114471	+	.	129	13	5105371_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5105371_2;MATENM=0;NM=1;NUMPARTS=6;REPSEQ=TTT;SCTG=c_12_15092001_15117001_201C;SPAN=10813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:134 DP:253 GQ:99 PL:[374.0, 0.0, 238.6] SR:13 DR:129 LR:-375.3 LO:375.3);ALT=T[chr12:15114471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16018671	+	chr12	16021662	+	.	30	22	5106892_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TAAA;MAPQ=60;MATEID=5106892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_15998501_16023501_183C;SPAN=2991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:58 GQ:17.3 PL:[122.9, 0.0, 17.3] SR:22 DR:30 LR:-127.4 LO:127.4);ALT=A[chr12:16021662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16064398	+	chr12	16111118	+	.	22	0	5107207_1	59.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5107207_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:16064398(+)-12:16111118(-)__12_16096501_16121501D;SPAN=46720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:49 GQ:59.3 PL:[59.3, 0.0, 59.3] SR:0 DR:22 LR:-59.35 LO:59.35);ALT=G[chr12:16111118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16109968	+	chr12	16111119	+	.	0	10	5107241_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=5107241_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_12_16096501_16121501_144C;SPAN=1151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:10 DR:0 LR:-7.814 LO:19.72);ALT=G[chr12:16111119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16109968	+	chr12	16112761	+	CTGCTTGGCTCCTGAAAGCTGTTACCTTTATAGATCTTACTACACTTTCAGGTGATGATACATCTTCCAACATTCAAAGGCTCTGTTATAAAGCCAAATACCCAATCCGGGAAGATCTCTTAAAAGCTTTAAATATGCATGATAA	0	23	5107242_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTGCTTGGCTCCTGAAAGCTGTTACCTTTATAGATCTTACTACACTTTCAGGTGATGATACATCTTCCAACATTCAAAGGCTCTGTTATAAAGCCAAATACCCAATCCGGGAAGATCTCTTAAAAGCTTTAAATATGCATGATAA;MAPQ=60;MATEID=5107242_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_16096501_16121501_144C;SPAN=2793;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:73 GQ:56.3 PL:[56.3, 0.0, 119.0] SR:23 DR:0 LR:-56.15 LO:57.45);ALT=G[chr12:16112761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16420123	+	chr12	16421291	+	TGTGCTTA	40	38	5107951_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TGTGCTTA;MAPQ=60;MATEID=5107951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_16415001_16440001_122C;SPAN=1168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:48 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:38 DR:40 LR:-178.2 LO:178.2);ALT=T[chr12:16421291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16500741	+	chr12	16510533	+	.	80	0	5108242_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5108242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:16500741(+)-12:16510533(-)__12_16488501_16513501D;SPAN=9792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:80 DP:113 GQ:38.9 PL:[233.6, 0.0, 38.9] SR:0 DR:80 LR:-241.2 LO:241.2);ALT=C[chr12:16510533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16500832	+	chr12	16507164	+	.	76	4	5108243_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5108243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_16488501_16513501_187C;SPAN=6332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:93 GQ:11.7 PL:[247.5, 11.7, 0.0] SR:4 DR:76 LR:-252.9 LO:252.9);ALT=G[chr12:16507164[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16507312	+	chr12	16516727	+	.	11	16	5108341_1	70.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5108341_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_16513001_16538001_20C;SPAN=9415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:68 GQ:70.7 PL:[70.7, 0.0, 93.8] SR:16 DR:11 LR:-70.7 LO:70.89);ALT=G[chr12:16516727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16507314	+	chr12	16510537	+	.	10	78	5108260_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5108260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_16488501_16513501_72C;SPAN=3223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:167 GQ:99 PL:[238.7, 0.0, 166.1] SR:78 DR:10 LR:-239.3 LO:239.3);ALT=T[chr12:16510537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16510633	+	chr12	16516726	+	.	10	99	5108342_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=5108342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_16513001_16538001_119C;SPAN=6093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:65 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:99 DR:10 LR:-323.5 LO:323.5);ALT=G[chr12:16516726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	16555269	+	chr14	21852097	+	.	10	0	5667937_1	19.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=5667937_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:16555269(+)-14:21852097(-)__14_21829501_21854501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:0 DR:10 LR:-19.73 LO:22.76);ALT=G[chr14:21852097[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	17444827	+	chr12	17445938	+	.	57	50	5110035_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=5110035_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_17419501_17444501_23C;SPAN=1111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:0 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:50 DR:57 LR:-247.6 LO:247.6);ALT=C[chr12:17445938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20770122	+	chr14	20774044	+	.	8	0	5664758_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5664758_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:20770122(+)-14:20774044(-)__14_20751501_20776501D;SPAN=3922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:0 DR:8 LR:-3.109 LO:15.25);ALT=T[chr14:20774044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20779914	+	chr14	20781623	+	.	6	9	5665099_1	21.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TTACCTA;MAPQ=60;MATEID=5665099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_20776001_20801001_337C;SPAN=1709;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:80 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:9 DR:6 LR:-21.24 LO:28.16);ALT=A[chr14:20781623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20797477	+	chr14	20801410	+	.	13	0	5665146_1	29.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5665146_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:20797477(+)-14:20801410(-)__14_20776001_20801001D;SPAN=3933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:48 GQ:29.9 PL:[29.9, 0.0, 86.0] SR:0 DR:13 LR:-29.91 LO:31.44);ALT=T[chr14:20801410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20920609	+	chr14	20922727	+	.	27	30	5665280_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=5665280_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_20898501_20923501_283C;SPAN=2118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:107 GQ:99 PL:[116.3, 0.0, 142.7] SR:30 DR:27 LR:-116.3 LO:116.4);ALT=T[chr14:20922727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20937694	+	chr14	20940466	+	.	28	10	5665535_1	83.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5665535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_20923001_20948001_178C;SPAN=2772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:95 GQ:83.3 PL:[83.3, 0.0, 146.0] SR:10 DR:28 LR:-83.2 LO:84.17);ALT=G[chr14:20940466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	20940636	+	chr14	20942626	+	.	0	13	5665547_1	19.0	.	EVDNC=ASSMB;HOMSEQ=TACAG;MAPQ=60;MATEID=5665547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_20923001_20948001_244C;SPAN=1990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:86 GQ:19.7 PL:[19.7, 0.0, 188.0] SR:13 DR:0 LR:-19.61 LO:27.71);ALT=G[chr14:20942626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21490685	+	chr14	21493186	+	.	8	0	5666739_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5666739_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:21490685(+)-14:21493186(-)__14_21486501_21511501D;SPAN=2501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=G[chr14:21493186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21702388	+	chr14	21737457	+	TGTAGCTGAAGATCAAAAAAATCTCA	0	26	5667764_1	72.0	.	EVDNC=ASSMB;INSERTION=TGTAGCTGAAGATCAAAAAAATCTCA;MAPQ=52;MATEID=5667764_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21731501_21756501_268C;SPAN=35069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:48 GQ:43.1 PL:[72.8, 0.0, 43.1] SR:26 DR:0 LR:-73.21 LO:73.21);ALT=A[chr14:21737457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21731989	+	chr14	21737456	+	.	90	26	5667770_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5667770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21731501_21756501_115C;SPAN=5467;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:109 GQ:16.2 PL:[297.0, 16.2, 0.0] SR:26 DR:90 LR:-302.9 LO:302.9);ALT=C[chr14:21737456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21840205	+	chr14	21841497	+	.	0	25	5667968_1	57.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=39;MATEID=5667968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21829501_21854501_43C;SPAN=1292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:92 GQ:57.8 PL:[57.8, 0.0, 163.4] SR:25 DR:0 LR:-57.6 LO:60.51);ALT=T[chr14:21841497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21945487	+	chr14	21955606	+	.	37	0	5668366_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5668366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:21945487(+)-14:21955606(-)__14_21952001_21977001D;SPAN=10119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:37 LR:-118.8 LO:118.8);ALT=G[chr14:21955606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21945723	+	chr14	21955608	+	.	0	16	5668259_1	39.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5668259_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21927501_21952501_132C;SPAN=9885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:48 GQ:39.8 PL:[39.8, 0.0, 76.1] SR:16 DR:0 LR:-39.81 LO:40.45);ALT=G[chr14:21955608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	21952624	+	chr14	21954663	+	T	59	61	5668368_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=5668368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21952001_21977001_104C;SPAN=2039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:24 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:61 DR:59 LR:-274.0 LO:274.0);ALT=C[chr14:21954663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	22887925	+	chr14	22896680	+	.	0	9	5670799_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5670799_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_22883001_22908001_180C;SPAN=8755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:9 DR:0 LR:-5.597 LO:17.5);ALT=C[chr14:22896680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	22887927	+	chr14	22901657	+	.	65	6	5670800_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5670800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_22883001_22908001_354C;SPAN=13730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:92 GQ:24.8 PL:[196.4, 0.0, 24.8] SR:6 DR:65 LR:-203.6 LO:203.6);ALT=T[chr14:22901657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	22896837	+	chr14	22901664	+	.	16	0	5670826_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5670826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:22896837(+)-14:22901664(-)__14_22883001_22908001D;SPAN=4827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:105 GQ:24.5 PL:[24.5, 0.0, 229.1] SR:0 DR:16 LR:-24.37 LO:34.16);ALT=C[chr14:22901664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23044134	+	chr14	23057853	+	.	65	39	5671056_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5671056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23030001_23055001_142C;SPAN=13719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:60 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:39 DR:65 LR:-194.7 LO:194.7);ALT=C[chr14:23057853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23105129	+	chr14	23107949	+	.	23	40	5671237_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AAATTAAGACACTAGC;MAPQ=60;MATEID=5671237_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_14_23103501_23128501_73C;SPAN=2820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:32 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:40 DR:23 LR:-151.8 LO:151.8);ALT=C[chr14:23107949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23105129	+	chr14	23110702	+	AAGATACCATTTTATACCCACTATATTGTCAAGAAGCAAAAATATGACAATAACAAGTGTTGACGAGGATGTGGAGACTTAAAAAATTTACACTGCTAGTGGGAGCGTAAATTTATATAATTGCTTTGGAAAATAATTTGTCATGACCTTGTAAAGATGAACATTCACATACTCTGTGACCCAATAATTCTACTCCTAGGTAGAGAAACTTGCACATATGCCCCAGGAGACAAACAAGAATATGTATAGGGAAGGGGGAGAGGGGGAGGGAGGGAAAAGAGAGAGGGAGGGAGGGAGGGAC	6	70	5671238_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AAAAAATTTACACTGCTAG;INSERTION=AAGATACCATTTTATACCCACTATATTGTCAAGAAGCAAAAATATGACAATAACAAGTGTTGACGAGGATGTGGAGACTTAAAAAATTTACACTGCTAGTGGGAGCGTAAATTTATATAATTGCTTTGGAAAATAATTTGTCATGACCTTGTAAAGATGAACATTCACATACTCTGTGACCCAATAATTCTACTCCTAGGTAGAGAAACTTGCACATATGCCCCAGGAGACAAACAAGAATATGTATAGGGAAGGGGGAGAGGGGGAGGGAGGGAAAAGAGAGAGGGAGGGAGGGAGGGAC;MAPQ=60;MATEID=5671238_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_14_23103501_23128501_73C;SPAN=5573;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:25 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:70 DR:6 LR:-217.9 LO:217.9);ALT=C[chr14:23110702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23105156	+	chr14	23109270	+	.	25	0	5671239_1	79.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5671239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:23105156(+)-14:23109270(-)__14_23103501_23128501D;SPAN=4114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:29 GQ:4.5 PL:[79.2, 4.5, 0.0] SR:0 DR:25 LR:-80.54 LO:80.54);ALT=C[chr14:23109270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23108063	+	chr14	23109271	+	.	10	41	5671243_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AAAAAATTTACACTGCTAG;MAPQ=60;MATEID=5671243_2;MATENM=2;NM=0;NUMPARTS=4;REPSEQ=GGG;SCTG=c_14_23103501_23128501_73C;SPAN=1208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:25 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:41 DR:10 LR:-141.9 LO:141.9);ALT=G[chr14:23109271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23108113	+	chr14	23110701	+	.	10	0	5671244_1	28.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5671244_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:23108113(+)-14:23110701(-)__14_23103501_23128501D;SPAN=2588;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:16 GQ:8.9 PL:[28.7, 0.0, 8.9] SR:0 DR:10 LR:-29.16 LO:29.16);ALT=T[chr14:23110701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23109490	+	chr14	23110702	+	C	33	15	5671245_1	49.0	.	DISC_MAPQ=52;EVDNC=TSI_L;HOMSEQ=AAAAAATTTACACTGCTAG;INSERTION=C;MAPQ=60;MATEID=5671245_2;MATENM=0;NM=2;NUMPARTS=4;REPSEQ=AGGGAGGGAGGGAGGG;SCTG=c_14_23103501_23128501_73C;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:16 GQ:10.1 PL:[49.6, 10.1, 0.0] SR:15 DR:33 LR:-49.7 LO:49.7);ALT=A[chr14:23110702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23235975	+	chr14	23237164	+	CCACAGCGTCGCAGGGCCCTCGCAATGGCTTGGGAAACCGCTGACCACACGGCTCCTATTCCCAGTAGCCCCGTGCTGCTGTCGCCCACACTACCTCTTCCTTGCGGCTTCCGGCCCCCGCAGCCTCAGTACCTCTGCTATCTCTTTTGCAGAAGTC	32	82	5671528_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CAGGT;INSERTION=CCACAGCGTCGCAGGGCCCTCGCAATGGCTTGGGAAACCGCTGACCACACGGCTCCTATTCCCAGTAGCCCCGTGCTGCTGTCGCCCACACTACCTCTTCCTTGCGGCTTCCGGCCCCCGCAGCCTCAGTACCTCTGCTATCTCTTTTGCAGAAGTC;MAPQ=60;MATEID=5671528_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_23226001_23251001_366C;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:111 GQ:19.8 PL:[306.9, 19.8, 0.0] SR:82 DR:32 LR:-309.7 LO:309.7);ALT=T[chr14:23237164[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23282627	+	chr14	23284580	+	.	8	0	5671971_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5671971_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:23282627(+)-14:23284580(-)__14_23275001_23300001D;SPAN=1953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=T[chr14:23284580[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23299196	+	chr14	23302624	+	.	38	0	5672037_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5672037_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:23299196(+)-14:23302624(-)__14_23275001_23300001D;SPAN=3428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:56 GQ:24.5 PL:[110.3, 0.0, 24.5] SR:0 DR:38 LR:-113.2 LO:113.2);ALT=A[chr14:23302624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23299463	+	chr14	23302626	+	.	0	92	5672040_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5672040_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23275001_23300001_177C;SPAN=3163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:64 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:92 DR:0 LR:-270.7 LO:270.7);ALT=G[chr14:23302626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23299463	+	chr14	23303380	+	.	22	4	5672041_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5672041_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23275001_23300001_38C;SPAN=3917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:64 GQ:62 PL:[62.0, 0.0, 91.7] SR:4 DR:22 LR:-61.89 LO:62.24);ALT=G[chr14:23303380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23421895	+	chr14	23424309	+	.	0	19	5672290_1	51.0	.	EVDNC=ASSMB;HOMSEQ=CTT;MAPQ=60;MATEID=5672290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23422001_23447001_68C;SPAN=2414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:40 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:19 DR:0 LR:-51.91 LO:51.91);ALT=T[chr14:23424309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23421939	+	chr14	23426172	+	.	11	0	5673056_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5673056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:23421939(+)-14:23426172(-)__14_23397501_23422501D;SPAN=4233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:0 DR:11 LR:-25.75 LO:26.84);ALT=A[chr14:23426172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23424386	+	chr14	23426133	+	.	22	15	5672299_1	73.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5672299_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23422001_23447001_177C;SPAN=1747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:83 GQ:73.4 PL:[73.4, 0.0, 126.2] SR:15 DR:22 LR:-73.24 LO:74.06);ALT=C[chr14:23426133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23502885	+	chr14	23503893	+	.	0	30	5672469_1	68.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5672469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23495501_23520501_251C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:113 GQ:68.6 PL:[68.6, 0.0, 203.9] SR:30 DR:0 LR:-68.42 LO:72.25);ALT=T[chr14:23503893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23559845	+	chr14	23564183	+	GGAATTTGGCTGGAATGCAGCATGGGGTGTTGAGTGTTTCTGTAAATTTTCTAGCATTAGAG	0	17	5672578_1	35.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GGAATTTGGCTGGAATGCAGCATGGGGTGTTGAGTGTTTCTGTAAATTTTCTAGCATTAGAG;MAPQ=60;MATEID=5672578_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_23544501_23569501_127C;SPAN=4338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:78 GQ:35 PL:[35.0, 0.0, 153.8] SR:17 DR:0 LR:-34.99 LO:39.25);ALT=G[chr14:23564183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	23564829	+	chr14	23566865	+	.	10	2	5672603_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5672603_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_23544501_23569501_375C;SPAN=2036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:2 DR:10 LR:-9.219 LO:21.81);ALT=G[chr14:23566865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24098401	+	chr14	97971487	-	.	6	30	5674476_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATTTTATATGACAACCAGCAATGACCA;MAPQ=60;MATEID=5674476_2;MATENM=0;NM=17;NUMPARTS=2;SCTG=c_14_24083501_24108501_274C;SPAN=73873086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:12 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:30 DR:6 LR:-89.12 LO:89.12);ALT=A]chr14:97971487];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	24423126	+	chr14	24424243	+	.	82	72	5675227_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=29;MATEID=5675227_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24402001_24427001_377C;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:113 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:72 DR:82 LR:-389.5 LO:389.5);ALT=G[chr14:24424243[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24458285	+	chr14	24459390	+	.	33	35	5675564_1	99.0	.	DISC_MAPQ=29;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5675564_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24451001_24476001_239C;SPAN=1105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:116 GQ:99 PL:[150.2, 0.0, 130.4] SR:35 DR:33 LR:-150.2 LO:150.2);ALT=G[chr14:24459390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24563644	+	chr14	24566100	+	.	17	6	5675642_1	45.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5675642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24549001_24574001_177C;SPAN=2456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:76 GQ:45.5 PL:[45.5, 0.0, 137.9] SR:6 DR:17 LR:-45.43 LO:48.08);ALT=G[chr14:24566100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24681036	+	chr14	24682614	+	.	69	5	5676125_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5676125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24671501_24696501_263C;SPAN=1578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:100 GQ:38.9 PL:[203.9, 0.0, 38.9] SR:5 DR:69 LR:-210.4 LO:210.4);ALT=C[chr14:24682614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24687424	+	chr14	24701456	+	ACGCTGACCGGAAAGGAGATTGAGATTGACATTGAACCTACAGAC	55	114	5676272_1	99.0	.	DISC_MAPQ=26;EVDNC=TSI_G;HOMSEQ=AAGGTG;INSERTION=ACGCTGACCGGAAAGGAGATTGAGATTGACATTGAACCTACAGAC;MAPQ=60;MATEID=5676272_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_24696001_24721001_381C;SPAN=14032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:34 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:114 DR:55 LR:-435.7 LO:435.7);ALT=T[chr14:24701456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24702804	+	chr14	24704941	+	.	0	9	5676295_1	8.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5676295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24696001_24721001_145C;SPAN=2137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-8.035 LO:17.94);ALT=G[chr14:24704941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24740516	+	chr14	24767818	+	.	7	4	5676183_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5676183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24745001_24770001_335C;SPAN=27302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:4 DR:7 LR:-23.21 LO:23.34);ALT=G[chr14:24767818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24761806	+	chr14	24767818	+	.	0	8	5676231_1	8.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5676231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_24745001_24770001_246C;SPAN=6012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:8 DR:0 LR:-8.256 LO:16.17);ALT=G[chr14:24767818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	24910134	+	chr14	24911384	+	ACACCTGTGACTAAGACCCAGGCCTTGGGGGGTTGTGGGGCTTTGGTGATGGCTTTAGCCAGCAATTGGGTGGTCTCTAGGCGGCTGCCGAGAACCTCTTTTTGGAAGGTTTCATTCCAT	0	27	5676868_1	69.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ACACCTGTGACTAAGACCCAGGCCTTGGGGGGTTGTGGGGCTTTGGTGATGGCTTTAGCCAGCAATTGGGTGGTCTCTAGGCGGCTGCCGAGAACCTCTTTTTGGAAGGTTTCATTCCAT;MAPQ=60;MATEID=5676868_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_24892001_24917001_354C;SPAN=1250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:73 GQ:69.5 PL:[69.5, 0.0, 105.8] SR:27 DR:0 LR:-69.35 LO:69.81);ALT=T[chr14:24911384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	25043757	+	chr14	25045381	+	.	9	0	5677095_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5677095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:25043757(+)-14:25045381(-)__14_25039001_25064001D;SPAN=1624;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:0 DR:9 LR:-4.784 LO:17.36);ALT=T[chr14:25045381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	25044071	+	chr14	25045376	+	.	77	0	5677098_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5677098_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:25044071(+)-14:25045376(-)__14_25039001_25064001D;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:94 GQ:2.1 PL:[231.0, 2.1, 0.0] SR:0 DR:77 LR:-243.1 LO:243.1);ALT=C[chr14:25045376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	96968937	+	chr14	96986392	+	.	0	66	5856503_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5856503_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_96946501_96971501_183C;SPAN=17455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:138 GQ:99 PL:[180.5, 0.0, 154.1] SR:66 DR:0 LR:-180.6 LO:180.6);ALT=T[chr14:96986392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	96969237	+	chr14	96986390	+	.	71	0	5856512_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5856512_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:96969237(+)-14:96986390(-)__14_96946501_96971501D;SPAN=17153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:53 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=C[chr14:96986390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	96991730	+	chr14	96993765	+	.	2	3	5856321_1	0	.	DISC_MAPQ=40;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=5856321_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_96971001_96996001_157C;SPAN=2035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:3 DR:2 LR:6.574 LO:6.671);ALT=T[chr14:96993765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	97027049	+	chr14	97029154	+	.	2	4	5856172_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5856172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_97020001_97045001_241C;SPAN=2105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:67 GQ:1.7 PL:[1.7, 0.0, 160.1] SR:4 DR:2 LR:-1.654 LO:11.33);ALT=G[chr14:97029154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	97263828	+	chr14	97299802	+	.	11	0	5857201_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5857201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:97263828(+)-14:97299802(-)__14_97289501_97314501D;SPAN=35974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:0 DR:11 LR:-25.75 LO:26.84);ALT=A[chr14:97299802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	97322925	+	chr14	97326892	+	.	3	6	5857328_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5857328_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_97314001_97339001_173C;SPAN=3967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:6 DR:3 LR:-6.631 LO:15.85);ALT=T[chr14:97326892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	97342459	+	chr14	97347514	+	.	2	4	5857374_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=5857374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_97338501_97363501_150C;SPAN=5055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:77 GQ:4.2 PL:[0.0, 4.2, 194.7] SR:4 DR:2 LR:4.356 LO:8.718);ALT=T[chr14:97347514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	98784003	+	chr14	98785088	+	.	51	34	5860915_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATTATGAATTGAAAGATTTTTTT;MAPQ=60;MATEID=5860915_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_98784001_98809001_258C;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:275 GQ:99 PL:[143.5, 0.0, 523.1] SR:34 DR:51 LR:-143.4 LO:155.6);ALT=T[chr14:98785088[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
