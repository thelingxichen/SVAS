chr10	89619592	+	chr18	20574391	+	TGGCGGGCA	0	50	9929260_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GTCAGGAGATCGAGACCATCCTG;INSERTION=TGGCGGGCA;MAPQ=60;MATEID=9929260_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_20555501_20580501_30C;SECONDARY;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:17 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:50 DR:0 LR:-148.5 LO:148.5);ALT=G[chr18:20574391[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr18	20101032	+	chr18	20096522	+	TTTGCAGTA	9	6	9927557_1	1.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TTTGCAGTA;MAPQ=60;MATEID=9927557_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_20090001_20115001_369C;SPAN=4510;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:143 GQ:1.1 PL:[1.1, 0.0, 344.3] SR:6 DR:9 LR:-0.8698 LO:22.31);ALT=]chr18:20101032]T;VARTYPE=BND:DUP-th;JOINTYPE=th
