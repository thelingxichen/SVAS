chr22	20950623	+	chr22	20953840	+	.	54	39	10844014_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=10844014_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_20947501_20972501_214C;SPAN=3217;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:12 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:39 DR:54 LR:-237.7 LO:237.7);ALT=C[chr22:20953840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
