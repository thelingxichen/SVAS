chr4	170190508	+	chr4	170192038	+	.	19	0	2329695_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2329695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:170190508(+)-4:170192038(-)__4_170177001_170202001D;SPAN=1530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:74 GQ:42.8 PL:[42.8, 0.0, 135.2] SR:0 DR:19 LR:-42.67 LO:45.43);ALT=A[chr4:170192038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	170671877	+	chr4	170674827	+	.	0	9	2331565_1	7.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2331565_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_170667001_170692001_282C;SPAN=2950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:9 DR:0 LR:-6.951 LO:17.74);ALT=C[chr4:170674827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	170671906	+	chr4	170678979	+	.	11	0	2331566_1	8.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2331566_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:170671906(+)-4:170678979(-)__4_170667001_170692001D;SPAN=7073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:0 DR:11 LR:-8.677 LO:21.71);ALT=T[chr4:170678979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	170674989	+	chr4	170678981	+	.	14	3	2331578_1	16.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2331578_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_170667001_170692001_60C;SPAN=3992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:109 GQ:16.7 PL:[16.7, 0.0, 247.7] SR:3 DR:14 LR:-16.68 LO:28.77);ALT=G[chr4:170678981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
