chr9	23362801	+	chr9	23377686	+	GA	0	33	5800729_1	95.0	.	EVDNC=ASSMB;INSERTION=GA;MAPQ=60;MATEID=5800729_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_23373001_23398001_110C;SPAN=14885;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:33 DP:7 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:33 DR:0 LR:-95.72 LO:95.72);ALT=A[chr9:23377686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
