chr17	5143547	+	chr17	5144658	+	.	8	0	9485330_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=9485330_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5143547(+)-17:5144658(-)__17_5120501_5145501D;SPAN=1111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:151 GQ:14.2 PL:[0.0, 14.2, 392.7] SR:0 DR:8 LR:14.5 LO:13.22);ALT=C[chr17:5144658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5902766	+	chr17	5903795	-	.	9	0	9488999_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=9488999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5902766(+)-17:5903795(+)__17_5880001_5905001D;SPAN=1029;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:141 GQ:8.1 PL:[0.0, 8.1, 356.4] SR:0 DR:9 LR:8.491 LO:15.62);ALT=A]chr17:5903795];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	6057534	-	chr17	6059384	+	.	11	0	9490004_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=9490004_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:6057534(-)-17:6059384(-)__17_6051501_6076501D;SPAN=1850;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:137 GQ:0.6 PL:[0.0, 0.6, 333.3] SR:0 DR:11 LR:0.8057 LO:20.23);ALT=[chr17:6059384[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
