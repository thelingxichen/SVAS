chr8	68311601	+	chr8	68761635	+	GG	52	55	5496681_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=GG;MAPQ=60;MATEID=5496681_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_8_68747001_68772001_0C;SPAN=450034;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:10 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:55 DR:52 LR:-267.4 LO:267.4);ALT=A[chr8:68761635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
