chr8	71354477	+	chr8	71353380	+	.	12	0	5501304_1	25.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5501304_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:71353380(-)-8:71354477(+)__8_71344001_71369001D;SPAN=1097;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=]chr8:71354477]A;VARTYPE=BND:DUP-th;JOINTYPE=th
