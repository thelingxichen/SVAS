chr1	153434943	+	chr1	153386986	+	.	0	11	551641_1	11.0	.	EVDNC=ASSMB;HOMSEQ=TGCTCCACATC;MAPQ=60;MATEID=551641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_153419001_153444001_28C;SPAN=47957;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:93 GQ:11.3 PL:[11.3, 0.0, 212.6] SR:11 DR:0 LR:-11.12 LO:22.18);ALT=]chr1:153434943]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	153842762	-	chr1	153843790	+	.	8	0	553431_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=553431_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153842762(-)-1:153843790(-)__1_153835501_153860501D;SPAN=1028;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:150 GQ:14.2 PL:[0.0, 14.2, 392.7] SR:0 DR:8 LR:14.23 LO:13.25);ALT=[chr1:153843790[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
