chr11	8839663	+	chr4	109329904	+	.	19	44	6636338_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;MAPQ=38;MATEID=6636338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_8820001_8845001_288C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:55 DP:37 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:44 DR:19 LR:-161.7 LO:161.7);ALT=]chr11:8839663]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	109721097	+	chr4	109722216	+	.	73	32	2833904_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TGGGGTTTCACCATGTTGGCCAGGCTGGTCTTGAACTCCTGACCT;MAPQ=60;MATEID=2833904_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_4_109711001_109736001_449C;SPAN=1119;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:80 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:32 DR:73 LR:-290.5 LO:290.5);ALT=T[chr4:109722216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	9104550	+	chr11	83028918	-	G	29	54	6979513_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=6979513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_83006001_83031001_252C;SPAN=73924368;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:70 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:54 DR:29 LR:-208.0 LO:208.0);ALT=T]chr11:83028918];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	82835551	+	chr11	82860295	+	.	7	3	6978512_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6978512_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_82859001_82884001_222C;SPAN=24744;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:3 DR:7 LR:-8.798 LO:16.28);ALT=T[chr11:82860295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
