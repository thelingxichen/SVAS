chr2	60773428	+	chr2	60778002	+	.	9	0	812999_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=812999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:60773428(+)-2:60778002(-)__2_60760001_60785001D;SPAN=4574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:101 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.346 LO:16.98);ALT=A[chr2:60778002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	60773435	+	chr2	60780351	+	.	0	42	813000_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=813000_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_60760001_60785001_247C;SPAN=6916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:99 GQ:99 PL:[111.8, 0.0, 128.3] SR:42 DR:0 LR:-111.8 LO:111.9);ALT=G[chr2:60780351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	61108988	+	chr2	61118817	+	.	0	11	813904_1	7.0	.	EVDNC=ASSMB;HOMSEQ=GGTG;MAPQ=60;MATEID=813904_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_61103001_61128001_245C;SPAN=9829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:11 DR:0 LR:-7.051 LO:21.42);ALT=G[chr2:61118817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	61118960	+	chr2	61121529	+	.	4	3	813938_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=813938_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_61103001_61128001_200C;SPAN=2569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:3 DR:4 LR:0.4634 LO:12.88);ALT=G[chr2:61121529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	61244986	+	chr2	61258554	+	.	6	2	814392_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=814392_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_61250001_61275001_104C;SPAN=13568;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:52 GQ:9.2 PL:[9.2, 0.0, 114.8] SR:2 DR:6 LR:-9.019 LO:14.54);ALT=A[chr2:61258554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	61293162	+	chr2	61295982	+	.	10	1	814507_1	14.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=814507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_61274501_61299501_26C;SPAN=2820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:1 DR:10 LR:-13.82 LO:22.76);ALT=G[chr2:61295982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	61700753	+	chr2	61703458	-	.	25	31	815792_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=ATT;MAPQ=60;MATEID=815792_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_61691001_61716001_292C;SPAN=2705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:52 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:31 DR:25 LR:-151.8 LO:151.8);ALT=T]chr2:61703458];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	61700774	-	chr2	61703160	+	.	54	25	815793_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCTCAGCCTCCCCAGTAGCTGGGA;MAPQ=60;MATEID=815793_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_61691001_61716001_29C;SPAN=2386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:25 DR:54 LR:-208.0 LO:208.0);ALT=[chr2:61703160[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	62095843	+	chr2	62099213	+	.	5	5	817424_1	10.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=TTACCT;MAPQ=60;MATEID=817424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62083001_62108001_325C;SPAN=3370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:5 DR:5 LR:-10.52 LO:20.25);ALT=T[chr2:62099213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62096690	+	chr2	62099216	+	.	9	8	817428_1	32.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=817428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62083001_62108001_82C;SPAN=2526;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:75 GQ:32.6 PL:[32.6, 0.0, 148.1] SR:8 DR:9 LR:-32.5 LO:36.77);ALT=T[chr2:62099216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62100430	+	chr2	62103230	+	.	4	3	817444_1	2.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=817444_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62083001_62108001_177C;SPAN=2800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:3 DR:4 LR:-2.788 LO:13.35);ALT=T[chr2:62103230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62104651	+	chr2	62106001	+	.	4	6	817461_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=817461_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62083001_62108001_299C;SPAN=1350;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:84 GQ:10.4 PL:[10.4, 0.0, 191.9] SR:6 DR:4 LR:-10.25 LO:20.2);ALT=T[chr2:62106001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62110729	+	chr2	62115515	+	.	12	0	817499_1	17.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=817499_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:62110729(+)-2:62115515(-)__2_62107501_62132501D;SPAN=4786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:0 DR:12 LR:-17.4 LO:25.39);ALT=A[chr2:62115515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62112255	+	chr2	62115687	+	.	16	0	817515_1	27.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=817515_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:62112255(+)-2:62115687(-)__2_62107501_62132501D;SPAN=3432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:95 GQ:27.2 PL:[27.2, 0.0, 202.1] SR:0 DR:16 LR:-27.08 LO:34.93);ALT=T[chr2:62115687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62132993	+	chr2	62227834	+	.	40	27	817700_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=817700_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62205501_62230501_203C;SPAN=94841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:45 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:27 DR:40 LR:-148.5 LO:148.5);ALT=G[chr2:62227834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	62423490	+	chr2	62449345	+	.	0	13	818244_1	28.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=818244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_62401501_62426501_346C;SPAN=25855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:54 GQ:28.4 PL:[28.4, 0.0, 101.0] SR:13 DR:0 LR:-28.28 LO:30.66);ALT=G[chr2:62449345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
