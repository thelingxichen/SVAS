chr13	99853223	+	chr13	99896083	+	.	12	0	5617659_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5617659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:99853223(+)-13:99896083(-)__13_99886501_99911501D;SPAN=42860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:0 DR:12 LR:-30.4 LO:30.71);ALT=C[chr13:99896083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	99853223	+	chr13	99890677	+	.	19	0	5617658_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5617658_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:99853223(+)-13:99890677(-)__13_99886501_99911501D;SPAN=37454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:44 GQ:50.9 PL:[50.9, 0.0, 54.2] SR:0 DR:19 LR:-50.8 LO:50.81);ALT=C[chr13:99890677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	99890808	+	chr13	99896769	+	ATTTGGAGGTTGATATGTGGAAGAATAATTTGCCTTGATTTGAAAGATACTTTCTGCAGTAGTCTGCTTATTTATAATTTTAGGATATTTGAAAGAAGATATGGAAGCAGAAAATTTGCA	2	20	5617673_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATTTGGAGGTTGATATGTGGAAGAATAATTTGCCTTGATTTGAAAGATACTTTCTGCAGTAGTCTGCTTATTTATAATTTTAGGATATTTGAAAGAAGATATGGAAGCAGAAAATTTGCA;MAPQ=60;MATEID=5617673_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_99886501_99911501_124C;SPAN=5961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:87 GQ:45.8 PL:[45.8, 0.0, 164.6] SR:20 DR:2 LR:-45.75 LO:49.56);ALT=G[chr13:99896769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	99948417	+	chr13	99959594	+	.	41	6	5617468_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5617468_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_99935501_99960501_50C;SPAN=11177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:105 GQ:99 PL:[110.3, 0.0, 143.3] SR:6 DR:41 LR:-110.2 LO:110.5);ALT=T[chr13:99959594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	100189036	+	chr13	100190067	+	.	9	0	5618498_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5618498_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:100189036(+)-13:100190067(-)__13_100180501_100205501D;SPAN=1031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:0 DR:9 LR:-9.119 LO:18.15);ALT=T[chr13:100190067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	100193922	+	chr13	100196116	+	.	2	4	5618513_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5618513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_100180501_100205501_255C;SPAN=2194;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:83 GQ:5.7 PL:[0.0, 5.7, 211.2] SR:4 DR:2 LR:5.982 LO:8.55);ALT=G[chr13:100196116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	100207902	+	chr13	100211615	+	.	5	3	5618551_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5618551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_100205001_100230001_356C;SPAN=3713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:80 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:3 DR:5 LR:-1.433 LO:13.15);ALT=G[chr13:100211615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	100211789	+	chr13	100214943	+	.	8	9	5618561_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5618561_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_100205001_100230001_220C;SPAN=3154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:75 GQ:32.6 PL:[32.6, 0.0, 148.1] SR:9 DR:8 LR:-32.5 LO:36.77);ALT=G[chr13:100214943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
