chr4	69373760	+	chr4	69491085	+	.	13	0	2743943_1	37.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2743943_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:69373760(+)-4:69491085(-)__4_69359501_69384501D;SPAN=117325;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:20 GQ:11 PL:[37.4, 0.0, 11.0] SR:0 DR:13 LR:-38.29 LO:38.29);ALT=T[chr4:69491085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	70039757	+	chr4	70180417	-	.	8	0	2745066_1	17.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2745066_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70039757(+)-4:70180417(+)__4_70021001_70046001D;SPAN=140660;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:0 DR:8 LR:-17.2 LO:18.78);ALT=A]chr4:70180417];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	70088022	+	chr4	70135840	-	.	19	0	2745190_1	56.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2745190_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70088022(+)-4:70135840(+)__4_70119001_70144001D;SPAN=47818;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:19 DP:8 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:0 DR:19 LR:-56.11 LO:56.11);ALT=G]chr4:70135840];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	70107391	-	chr4	70174159	+	.	9	0	2745302_1	18.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2745302_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70107391(-)-4:70174159(-)__4_70168001_70193001D;SPAN=66768;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:43 GQ:18.2 PL:[18.2, 0.0, 84.2] SR:0 DR:9 LR:-18.06 LO:20.6);ALT=[chr4:70174159[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	70107422	-	chr4	70173806	+	.	16	0	2745303_1	46.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2745303_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70107422(-)-4:70173806(-)__4_70168001_70193001D;SPAN=66384;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:16 DP:15 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:0 DR:16 LR:-46.21 LO:46.21);ALT=[chr4:70173806[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	70108182	+	chr4	70173131	-	.	12	0	2745305_1	33.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=2745305_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70108182(+)-4:70173131(+)__4_70168001_70193001D;SPAN=64949;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:12 DP:3 GQ:3 PL:[33.0, 3.0, 0.0] SR:0 DR:12 LR:-33.01 LO:33.01);ALT=T]chr4:70173131];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	70780008	+	chr4	70435023	+	.	59	49	2747119_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=2747119_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_70756001_70781001_3C;SPAN=344985;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:41 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:49 DR:59 LR:-244.3 LO:244.3);ALT=]chr4:70780008]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	70459360	+	chr4	70504417	+	GCATAAAATGCTATCCAT	38	50	2745867_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GCATAAAATGCTATCCAT;MAPQ=60;MATEID=2745867_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_70437501_70462501_256C;SPAN=45057;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:36 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:50 DR:38 LR:-208.0 LO:208.0);ALT=A[chr4:70504417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
