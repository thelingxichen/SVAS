chr6	37479956	+	chr6	46297896	+	.	0	22	6205266_1	58.0	.	BX=TCAATCTAGCGATATA-1_1,CGCTATCCAGACTATC-1_1,GCGCTAGCACCATGAT-1_1,GATGGTTTCAAACCGT-1_1,GGTGGCTAGTCCCGGT-1_1,TTAGGACCACGTCCGA-1_1,ACGATCATCACGGTAT-1_1,TAACTCTAGTCGGTCC-1_1,GTGCAGCAGTCCTCCT-1_1,CGGAGCTGTAAGTAAC-1_1,CTACCCATCTGTGCAA-1_1,ACCGTAAAGACTAGAT-1_1,ACCACGGGTAGTTGGG-1_1,GATGGTTGTGACGCCT-1_1,TGGCATAAGCGGTGAT-1_1,TAGAGCTTCGCATGAT-1_1,GTCGACGTCGGTGGCT-1_1,CCTAGTCCACATGCGC-1_1,GGGCCATGTACGAGGT-1_1;EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6205266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_46280501_46305501_83C;SPAN=8817940;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:46 GQ:12.6 PL:[0.0, 12.6, 138.6] SR:0 DR:0 LR:12.92 LO:0.0),OC001T.bam(GT:0/1 AD:22 DP:50 GQ:58.7 PL:[58.7, 0.0, 65.3] SR:22 DR:0 LR:-58.57 LO:58.61);ALT=g[chr6:46297896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht	.
chr6	37479956	+	chr6	46297896	+	.	0	22	6205266_1	58.0	.	BX=TCAATCTAGCGATATA-1_1,CGCTATCCAGACTATC-1_1,GCGCTAGCACCATGAT-1_1,GATGGTTTCAAACCGT-1_1,GGTGGCTAGTCCCGGT-1_1,TTAGGACCACGTCCGA-1_1,ACGATCATCACGGTAT-1_1,TAACTCTAGTCGGTCC-1_1,GTGCAGCAGTCCTCCT-1_1,CGGAGCTGTAAGTAAC-1_1,CTACCCATCTGTGCAA-1_1,ACCGTAAAGACTAGAT-1_1,ACCACGGGTAGTTGGG-1_1,GATGGTTGTGACGCCT-1_1,TGGCATAAGCGGTGAT-1_1,TAGAGCTTCGCATGAT-1_1,GTCGACGTCGGTGGCT-1_1,CCTAGTCCACATGCGC-1_1,GGGCCATGTACGAGGT-1_1;EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6205266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_46280501_46305501_83C;SPAN=8817940;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:46 GQ:12.6 PL:[0.0, 12.6, 138.6] SR:0 DR:0 LR:12.92 LO:0.0),OC001T.bam(GT:0/1 AD:22 DP:50 GQ:58.7 PL:[58.7, 0.0, 65.3] SR:22 DR:0 LR:-58.57 LO:58.61);ALT=g[chr6:46297896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht	.
