chr1	43694063	+	chr1	43695544	+	.	62	38	218436_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=218436_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_43683501_43708501_309C;SPAN=1481;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:77 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:38 DR:62 LR:-257.5 LO:257.5);ALT=G[chr1:43695544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
