chr3	6815013	+	chr5	68513729	-	.	19	0	2494161_1	53.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2494161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:6815013(+)-5:68513729(+)__5_68502001_68527001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:34 GQ:27.2 PL:[53.6, 0.0, 27.2] SR:0 DR:19 LR:-53.9 LO:53.9);ALT=C]chr5:68513729];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	67511783	+	chr5	67522115	+	.	39	25	2492499_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAGGT;MAPQ=60;MATEID=2492499_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_67522001_67547001_90C;SPAN=10332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:35 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:25 DR:39 LR:-161.7 LO:161.7);ALT=T[chr5:67522115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	68513733	+	chr5	68524025	+	.	67	0	2494191_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2494191_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:68513733(+)-5:68524025(-)__5_68502001_68527001D;SPAN=10292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:66 GQ:18 PL:[198.0, 18.0, 0.0] SR:0 DR:67 LR:-198.0 LO:198.0);ALT=G[chr5:68524025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	68661581	+	chr12	34402512	-	.	15	0	5152472_1	40.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5152472_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:68661581(+)-12:34402512(+)__12_34398001_34423001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:33 GQ:37.4 PL:[40.7, 0.0, 37.4] SR:0 DR:15 LR:-40.58 LO:40.58);ALT=A]chr12:34402512];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	68661634	+	chr5	68665286	+	.	43	0	2494428_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2494428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:68661634(+)-5:68665286(-)__5_68649001_68674001D;SPAN=3652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:63 GQ:26 PL:[125.0, 0.0, 26.0] SR:0 DR:43 LR:-128.3 LO:128.3);ALT=T[chr5:68665286[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	32832399	+	chr12	32854346	+	.	0	16	5148769_1	31.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=5148769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_32830001_32855001_235C;SPAN=21947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:79 GQ:31.4 PL:[31.4, 0.0, 160.1] SR:16 DR:0 LR:-31.41 LO:36.36);ALT=G[chr12:32854346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	33296559	+	chr12	33307367	+	.	40	43	5149898_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=CCTGAG;MAPQ=60;MATEID=5149898_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_33295501_33320501_72C;SPAN=10808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:36 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:43 DR:40 LR:-194.7 LO:194.7);ALT=G[chr12:33307367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	33715123	+	chr12	33716966	+	.	38	27	5150885_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AACAA;MAPQ=60;MATEID=5150885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_33712001_33737001_297C;SPAN=1843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:74 GQ:26.3 PL:[151.7, 0.0, 26.3] SR:27 DR:38 LR:-156.4 LO:156.4);ALT=A[chr12:33716966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	34845064	+	chr12	34849138	+	.	69	28	5153403_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CTTTGTGATGTGTGCATTCAACTCACAGAGTTTAACCTT;MAPQ=60;MATEID=5153403_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_34839001_34864001_134C;SPAN=4074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:21 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:28 DR:69 LR:-270.7 LO:270.7);ALT=T[chr12:34849138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
