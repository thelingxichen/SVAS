chr1	214656755	+	chr5	115177749	-	.	62	0	2559812_1	99.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2559812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:214656755(+)-5:115177749(+)__5_115174501_115199501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:32 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:0 DR:62 LR:-181.5 LO:181.5);ALT=G]chr5:115177749];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	214776664	+	chr1	214787055	+	.	11	4	540341_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=540341_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_214767001_214792001_105C;SPAN=10391;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:99 GQ:12.8 PL:[12.8, 0.0, 227.3] SR:4 DR:11 LR:-12.79 LO:24.33);ALT=G[chr1:214787055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115173466	+	chr5	115177020	+	.	11	0	2559815_1	28.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=2559815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115173466(+)-5:115177020(-)__5_115174501_115199501D;SPAN=3554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:28 GQ:28.7 PL:[28.7, 0.0, 38.6] SR:0 DR:11 LR:-28.73 LO:28.81);ALT=A[chr5:115177020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	71064319	+	chr5	115177196	+	.	15	0	6490193_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6490193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115177196(-)-17:71064319(+)__17_71050001_71075001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:45 GQ:37.4 PL:[37.4, 0.0, 70.4] SR:0 DR:15 LR:-37.32 LO:37.92);ALT=]chr17:71064319]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	115177773	+	chr5	115205712	+	.	13	0	2559822_1	34.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2559822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115177773(+)-5:115205712(-)__5_115174501_115199501D;SPAN=27939;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:30 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:0 DR:13 LR:-34.79 LO:34.79);ALT=G[chr5:115205712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115420829	+	chr5	115426772	+	.	10	0	2560102_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2560102_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:115420829(+)-5:115426772(-)__5_115419501_115444501D;SPAN=5943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=G[chr5:115426772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	115426887	+	chr5	115428240	+	.	0	4	2560113_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2560113_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_5_115419501_115444501_180C;SPAN=1353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:49 GQ:0 PL:[0.0, 0.0, 118.8] SR:4 DR:0 LR:0.0713 LO:7.387);ALT=G[chr5:115428240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	70301136	+	chr17	70300006	+	.	50	0	6488034_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6488034_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:70300006(-)-17:70301136(+)__17_70290501_70315501D;SPAN=1130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:133 GQ:99 PL:[129.2, 0.0, 191.9] SR:0 DR:50 LR:-129.0 LO:129.7);ALT=]chr17:70301136]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	71027854	+	chr17	71084796	+	CCTGCAGCAAAGCCAAGACTTCCATCTAAGATCCGCCT	0	10	6490279_1	20.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CCTGCAGCAAAGCCAAGACTTCCATCTAAGATCCGCCT;MAPQ=60;MATEID=6490279_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_71074501_71099501_61C;SPAN=56942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:10 DR:0 LR:-20.82 LO:23.18);ALT=C[chr17:71084796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	71223406	+	chr17	71228224	+	.	0	7	6490775_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=6490775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_71221501_71246501_368C;SPAN=4818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:76 GQ:2.6 PL:[2.6, 0.0, 180.8] SR:7 DR:0 LR:-2.517 LO:13.31);ALT=G[chr17:71228224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
