chr6	15452408	+	chr6	15468771	+	.	5	3	2715497_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2715497_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_15459501_15484501_283C;SPAN=16363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:3 DR:5 LR:-3.059 LO:13.4);ALT=T[chr6:15468771[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	16145548	+	chr6	16146890	+	.	0	12	2717855_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=2717855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_16145501_16170501_296C;SPAN=1342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:129 GQ:4.7 PL:[4.7, 0.0, 308.3] SR:12 DR:0 LR:-4.663 LO:22.87);ALT=G[chr6:16146890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	16884968	+	chr6	16886094	+	.	52	48	2720775_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGA;MAPQ=60;MATEID=2720775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_16880501_16905501_63C;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:70 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:48 DR:52 LR:-234.4 LO:234.4);ALT=A[chr6:16886094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	17376781	+	chr6	17381279	+	.	46	31	2722352_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCTCACGCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=60;MATEID=2722352_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_17370501_17395501_235C;SECONDARY;SPAN=4498;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:31 DR:46 LR:-208.0 LO:208.0);ALT=C[chr6:17381279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18160214	+	chr6	18161556	+	.	0	5	2725756_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2725756_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_18154501_18179501_181C;SPAN=1342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:104 GQ:11.4 PL:[0.0, 11.4, 273.9] SR:5 DR:0 LR:11.67 LO:8.049);ALT=G[chr6:18161556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18225963	+	chr6	18236681	+	CTTTTACAGTTGTTTTTATGAAATCTTTTCTTTCAGTTAAATCATAAGTAGGATAATTTTCATAG	6	14	2725963_1	34.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=CTTTTACAGTTGTTTTTATGAAATCTTTTCTTTCAGTTAAATCATAAGTAGGATAATTTTCATAG;MAPQ=60;MATEID=2725963_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_18228001_18253001_115C;SPAN=10718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:44 GQ:34.4 PL:[34.4, 0.0, 70.7] SR:14 DR:6 LR:-34.29 LO:35.04);ALT=T[chr6:18236681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18237749	+	chr6	18249882	+	.	12	10	2725998_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2725998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_18228001_18253001_215C;SPAN=12133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:98 GQ:39.5 PL:[39.5, 0.0, 197.9] SR:10 DR:12 LR:-39.47 LO:45.53);ALT=T[chr6:18249882[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18250070	+	chr6	18258182	+	TTTGCCAGAAGGCTTTGGATGCATTAAGAAATTCAAGATCCTCTTCACTAGTTCACTATTTACACCTGATCTCTCCAAATCAAGAACCTCACAGATGCTCTTTAACATGGCATTTCTAAATTTTTTCAACATTTCTTCCTTCTTTTTATATTGGACACTTCCTTTTTCAAATGGAAAGCCACTGAACTGACCCACATTCTTCTTTAATGAGGAC	2	48	2726052_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=TTTGCCAGAAGGCTTTGGATGCATTAAGAAATTCAAGATCCTCTTCACTAGTTCACTATTTACACCTGATCTCTCCAAATCAAGAACCTCACAGATGCTCTTTAACATGGCATTTCTAAATTTTTTCAACATTTCTTCCTTCTTTTTATATTGGACACTTCCTTTTTCAAATGGAAAGCCACTGAACTGACCCACATTCTTCTTTAATGAGGAC;MAPQ=60;MATEID=2726052_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_18252501_18277501_230C;SPAN=8112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:51 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:48 DR:2 LR:-148.5 LO:148.5);ALT=G[chr6:18258182[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18256724	+	chr6	18258244	+	.	8	0	2726073_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2726073_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:18256724(+)-6:18258244(-)__6_18252501_18277501D;SPAN=1520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=C[chr6:18258244[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18258638	+	chr6	18264614	+	TTTTCCTCCTCCTCCTCCTCCTCGTCGTCCTCGTCCTCTTCCTCCTCGCTCTCCTCTCTGGGACCGGGCATTTCGGGTTCTTTCTCGGACGCGGGCTGGGTGGGGGTTCCCTCCCCCTCCGCAGCAGGGGCCGAGGCGGACATGCTGTGA	13	70	2726081_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TTTTCCTCCTCCTCCTCCTCCTCGTCGTCCTCGTCCTCTTCCTCCTCGCTCTCCTCTCTGGGACCGGGCATTTCGGGTTCTTTCTCGGACGCGGGCTGGGTGGGGGTTCCCTCCCCCTCCGCAGCAGGGGCCGAGGCGGACATGCTGTGA;MAPQ=60;MATEID=2726081_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_18252501_18277501_40C;SPAN=5976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:87 GQ:3.6 PL:[217.8, 3.6, 0.0] SR:70 DR:13 LR:-228.1 LO:228.1);ALT=T[chr6:18264614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	18258638	+	chr6	18264082	+	TTT	2	19	2726080_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTT;MAPQ=60;MATEID=2726080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_18252501_18277501_121C;SPAN=5444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:113 GQ:38.9 PL:[38.9, 0.0, 233.6] SR:19 DR:2 LR:-38.71 LO:46.84);ALT=T[chr6:18264082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
