chr11	38760424	+	chr11	38761807	-	.	5	2	4830382_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCCTTTGGGTATA;MAPQ=60;MATEID=4830382_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_38759001_38784001_50C;SPAN=1383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:72 GQ:0.5 PL:[0.5, 0.0, 172.1] SR:2 DR:5 LR:-0.2994 LO:11.14);ALT=A]chr11:38761807];VARTYPE=BND:INV-hh;JOINTYPE=hh
