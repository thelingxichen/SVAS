chrY	21729368	+	chrY	21749095	+	.	21	2	7565353_1	66.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7565353_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_24_21707001_21732001_0C;SPAN=19727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:3 GQ:6 PL:[66.0, 6.0, 0.0] SR:2 DR:21 LR:-66.02 LO:66.02);ALT=G[chrY:21749095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	22737776	+	chrY	22741492	+	.	24	13	7565395_1	65.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGGTA;MAPQ=60;MATEID=7565395_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AGGAGG;SCTG=c_24_22736001_22761001_4C;SPAN=3716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:8 GQ:7.4 PL:[65.0, 7.4, 0.0] SR:13 DR:24 LR:-65.02 LO:65.02);ALT=A[chrY:22741492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	22737795	+	chrY	22744473	+	.	29	0	7565397_1	85.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7565397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=24:22737795(+)-24:22744473(-)__24_22736001_22761001D;SPAN=6678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:9 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=A[chrY:22744473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	22751461	+	chrY	22754227	+	.	0	11	7565402_1	29.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7565402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_24_22736001_22761001_5C;SPAN=2766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:5 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:11 DR:0 LR:-29.71 LO:29.71);ALT=T[chrY:22754227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
