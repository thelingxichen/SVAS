chrY	2709729	+	chrY	2712117	+	.	18	0	7562658_1	52.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7562658_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=24:2709729(+)-24:2712117(-)__24_2695001_2720001D;SPAN=2388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:12 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=T[chrY:2712117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	2710288	+	chrY	2712116	+	.	78	0	7562661_1	99.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=7562661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=24:2710288(+)-24:2712116(-)__24_2695001_2720001D;SPAN=1828;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:12 GQ:21 PL:[231.0, 21.0, 0.0] SR:0 DR:78 LR:-231.1 LO:231.1);ALT=G[chrY:2712116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	2710291	+	chrY	2713685	+	.	15	0	7562662_1	41.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=7562662_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=24:2710291(+)-24:2713685(-)__24_2695001_2720001D;SPAN=3394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:31 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:0 DR:15 LR:-41.15 LO:41.15);ALT=T[chrY:2713685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	2713784	+	chrY	2722639	+	.	5	17	7562667_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=7562667_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_24_2695001_2720001_2C;SPAN=8855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:10 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:17 DR:5 LR:-62.72 LO:62.72);ALT=G[chrY:2722639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	2722813	+	chrY	2733127	+	.	9	31	7562758_1	99.0	.	DISC_MAPQ=52;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=7562758_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_24_2719501_2744501_0C;SPAN=10314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:26 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:31 DR:9 LR:-118.8 LO:118.8);ALT=G[chrY:2733127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrY	2722813	+	chrY	2734834	+	CAATTTGTGTATGGTGATTGGTGGAGCCAACCTCGGTCGTGTTGGTGTGATCACCAACAGGGAAAGACATCCTGGTTCTTTTGATGTGGTGCATGTGAAGGATGCCAATGGCAACAGCTTTGCCACGAGGCTTTCCAACATTTTTGTCATTGGCAAT	0	143	7562759_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CAATTTGTGTATGGTGATTGGTGGAGCCAACCTCGGTCGTGTTGGTGTGATCACCAACAGGGAAAGACATCCTGGTTCTTTTGATGTGGTGCATGTGAAGGATGCCAATGGCAACAGCTTTGCCACGAGGCTTTCCAACATTTTTGTCATTGGCAAT;MAPQ=60;MATEID=7562759_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_24_2719501_2744501_0C;SPAN=12021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:56 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:143 DR:0 LR:-422.5 LO:422.5);ALT=G[chrY:2734834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
