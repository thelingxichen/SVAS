chr10	49893046	+	chr10	49917758	+	.	2	2	4593017_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4593017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_49906501_49931501_354C;SPAN=24712;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:21 GQ:7.7 PL:[7.7, 0.0, 40.7] SR:2 DR:2 LR:-7.515 LO:8.97);ALT=G[chr10:49917758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	50375074	+	chr10	50396338	+	.	10	0	4593451_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4593451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:50375074(+)-10:50396338(-)__10_50372001_50397001D;SPAN=21264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=T[chr10:50396338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
