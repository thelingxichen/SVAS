chr1	184814743	+	chr1	184820785	+	.	56	27	688584_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAATTTTAAAAAG;MAPQ=60;MATEID=688584_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_184803501_184828501_237C;SPAN=6042;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:72 DP:112 GQ:62.3 PL:[207.5, 0.0, 62.3] SR:27 DR:56 LR:-211.5 LO:211.5);ALT=G[chr1:184820785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	185025687	-	chr19	45828385	+	CACAAAAAATAAAAAAAACTACAAAAATTATCTGGGCGTAGTGGAGTGCATCTGTGGTCCCAGCTACTC	20	115	10324330_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=CACAAAAAATAAAAAAAACTACAAAAATTATCTGGGCGTAGTGGAGTGCATCTGTGGTCCCAGCTACTC;MAPQ=60;MATEID=10324330_2;MATENM=0;NM=6;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_19_45815001_45840001_480C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:129 DP:67 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:115 DR:20 LR:-382.9 LO:382.9);ALT=[chr19:45828385[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	185025805	+	chr19	45828412	-	GCTCAGGAGTTCAAGACCACCCTGGCCAACGCGGTGAAACCCTGTCTCTACTAAAAATACAAAAATTAGCCGGACATGGTGGGACACACCTATAGTCTCAGCTACTCAGGAGGCCGAGATGGGAGGATCACTTGAGCCTGGGGAGGTGAGGCTGCGGTGAGCTGTGATCGCACTGCTGCACTCCAGCCTTGGTGACAGAGCGAGACTGTGTCTAAAAAAAAAACAAAAAACAAAAAACAATTGAACTGAGGGAGACAGAGCAGAAGGATGGACTCCAGAGCCTGAGAAGGGTA	6	144	10324331_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=GCTCAGGAGTTCAAGACCACCCTGGCCAACGCGGTGAAACCCTGTCTCTACTAAAAATACAAAAATTAGCCGGACATGGTGGGACACACCTATAGTCTCAGCTACTCAGGAGGCCGAGATGGGAGGATCACTTGAGCCTGGGGAGGTGAGGCTGCGGTGAGCTGTGATCGCACTGCTGCACTCCAGCCTTGGTGACAGAGCGAGACTGTGTCTAAAAAAAAAACAAAAAACAAAAAACAATTGAACTGAGGGAGACAGAGCAGAAGGATGGACTCCAGAGCCTGAGAAGGGTA;MAPQ=60;MATEID=10324331_2;MATENM=0;NM=6;NUMPARTS=3;SCTG=c_19_45815001_45840001_480C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:147 DP:76 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:144 DR:6 LR:-435.7 LO:435.7);ALT=T]chr19:45828412];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	185698571	-	chr1	185699887	+	.	13	0	691720_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=691720_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:185698571(-)-1:185699887(-)__1_185685501_185710501D;SPAN=1316;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:136 GQ:6.2 PL:[6.2, 0.0, 323.0] SR:0 DR:13 LR:-6.067 LO:24.94);ALT=[chr1:185699887[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	186606581	+	chr1	189443822	-	.	23	0	708036_1	58.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=708036_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:186606581(+)-1:189443822(+)__1_189434001_189459001D;SPAN=2837241;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:64 GQ:58.7 PL:[58.7, 0.0, 95.0] SR:0 DR:23 LR:-58.58 LO:59.1);ALT=G]chr1:189443822];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	186606693	-	chr1	189443700	+	.	8	0	708037_1	2.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=708037_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:186606693(-)-1:189443700(-)__1_189434001_189459001D;SPAN=2837007;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-2.025 LO:15.08);ALT=[chr1:189443700[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	187464828	+	chr1	187466730	+	AATATGCTTTCTGTTTTTGGGTGTCACTCTCAATTTTTTTGAAACAATACATTTTTCCGTCTTACTTTAATTCATCCCTTGTCATCCATTTCTCATCCATTACATTCTAGCATTCATATCTATCCCTTCCCCACTGAAATCGATCTCACTAAGTCACTGATGTTCCCAAGTTTTTAACACAAGTTTCTGTCTTTGGTTTTCAGCCTAATTTTTTAGATATTACTACCAATAGAATGGTCTCCTGGATTT	22	174	698815_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=AATATGCTTTCTGTTTTTGGGTGTCACTCTCAATTTTTTTGAAACAATACATTTTTCCGTCTTACTTTAATTCATCCCTTGTCATCCATTTCTCATCCATTACATTCTAGCATTCATATCTATCCCTTCCCCACTGAAATCGATCTCACTAAGTCACTGATGTTCCCAAGTTTTTAACACAAGTTTCTGTCTTTGGTTTTCAGCCTAATTTTTTAGATATTACTACCAATAGAATGGTCTCCTGGATTT;MAPQ=60;MATEID=698815_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_187449501_187474501_273C;SPAN=1902;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:184 DP:48 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:174 DR:22 LR:-544.6 LO:544.6);ALT=T[chr1:187466730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	188198933	+	chr1	187721213	+	.	53	31	702508_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAA;MAPQ=60;MATEID=702508_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_188184501_188209501_229C;SPAN=477720;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:51 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:31 DR:53 LR:-201.3 LO:201.3);ALT=]chr1:188198933]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	188342935	-	chr11	40727082	+	.	8	23	702999_1	83.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=GAACTCATTCTTTTTTATGCCTGCATAGTATTCC;MAPQ=10;MATEID=702999_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_1_188331501_188356501_1C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:69 GQ:83.6 PL:[83.6, 0.0, 83.6] SR:23 DR:8 LR:-83.64 LO:83.64);ALT=[chr11:40727082[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	188806259	+	chr1	188807274	-	.	9	0	704338_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=704338_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:188806259(+)-1:188807274(+)__1_188797001_188822001D;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:134 GQ:6.3 PL:[0.0, 6.3, 336.6] SR:0 DR:9 LR:6.595 LO:15.83);ALT=C]chr1:188807274];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	40650725	+	chr11	40647110	+	CAC	4	3	6761143_1	0	.	DISC_MAPQ=47;EVDNC=ASDIS;INSERTION=CAC;MAPQ=46;MATEID=6761143_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_40645501_40670501_141C;SPAN=3615;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:126 GQ:17.4 PL:[0.0, 17.4, 339.9] SR:3 DR:4 LR:17.63 LO:7.626);ALT=]chr11:40650725]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	40734100	+	chr11	40682825	+	A	51	39	6761865_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=6761865_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_40719001_40744001_339C;SPAN=51275;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:55 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:39 DR:51 LR:-217.9 LO:217.9);ALT=]chr11:40734100]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	45067393	+	chr19	56442260	-	.	2	16	10382264_1	47.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATATA;MAPQ=37;MATEID=10382264_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_56423501_56448501_513C;SPAN=11374867;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:20 GQ:1.1 PL:[47.3, 0.0, 1.1] SR:16 DR:2 LR:-50.09 LO:50.09);ALT=T]chr19:56442260];VARTYPE=BND:INV-hh;JOINTYPE=hh
