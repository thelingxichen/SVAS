chr6	114223945	+	chr6	114225040	+	TTTTT	0	63	4362125_1	99.0	.	EVDNC=ASSMB;INSERTION=TTTTT;MAPQ=60;MATEID=4362125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_114219001_114244001_25C;SPAN=1095;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:24 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:63 DR:0 LR:-184.8 LO:184.8);ALT=A[chr6:114225040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	114953133	+	chr6	115295453	+	.	19	0	4364339_1	56.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=4364339_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:114953133(+)-6:115295453(-)__6_115272501_115297501D;SPAN=342320;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:19 DP:16 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:0 DR:19 LR:-56.11 LO:56.11);ALT=T[chr6:115295453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
