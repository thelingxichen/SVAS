chr1	196745109	+	chr1	196735808	+	.	40	0	733797_1	99.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=733797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:196735808(-)-1:196745109(+)__1_196735001_196760001D;SPAN=9301;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:108 GQ:99 PL:[102.8, 0.0, 158.9] SR:0 DR:40 LR:-102.8 LO:103.4);ALT=]chr1:196745109]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	196736078	+	chr1	196745437	+	.	10	0	733800_1	0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=733800_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:196736078(+)-1:196745437(-)__1_196735001_196760001D;SPAN=9359;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:120 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.4991 LO:18.56);ALT=A[chr1:196745437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	196936321	+	chr1	196937484	+	.	65	49	734062_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AACTT;MAPQ=60;MATEID=734062_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_196931001_196956001_197C;SPAN=1163;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:84 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:49 DR:65 LR:-260.8 LO:260.8);ALT=T[chr1:196937484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	197500520	+	chr1	197503272	+	.	139	99	737158_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AACAAATCTTTT;MAPQ=60;MATEID=737158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_197494501_197519501_99C;SPAN=2752;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:187 DP:59 GQ:50.5 PL:[554.5, 50.5, 0.0] SR:99 DR:139 LR:-554.5 LO:554.5);ALT=T[chr1:197503272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
