chr10	19986839	-	chr10	19987957	+	.	8	0	6126458_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6126458_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:19986839(-)-10:19987957(-)__10_19967501_19992501D;SPAN=1118;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:129 GQ:8.4 PL:[0.0, 8.4, 330.0] SR:0 DR:8 LR:8.541 LO:13.78);ALT=[chr10:19987957[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
