chr4	164415956	+	chr4	164428184	+	.	7	10	2311592_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2311592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_164395001_164420001_212C;SPAN=12228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:63 GQ:32.6 PL:[32.6, 0.0, 118.4] SR:10 DR:7 LR:-32.45 LO:35.29);ALT=G[chr4:164428184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	164507088	+	chr4	164534466	+	.	13	9	2311694_1	40.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTGCAGA;MAPQ=60;MATEID=2311694_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_164517501_164542501_389C;SPAN=27378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:45 GQ:40.7 PL:[40.7, 0.0, 67.1] SR:9 DR:13 LR:-40.62 LO:41.02);ALT=A[chr4:164534466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
