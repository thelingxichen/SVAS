chrX	30578475	+	chrX	30594869	+	.	0	9	7392049_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7392049_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_30576001_30601001_96C;SPAN=16394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:9 DR:0 LR:-14.27 LO:19.37);ALT=T[chrX:30594869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	30578515	+	chrX	30595769	+	.	11	0	7392050_1	17.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7392050_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:30578515(+)-23:30595769(-)__23_30576001_30601001D;SPAN=17254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=C[chrX:30595769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	30820351	+	chrX	30819339	+	.	15	0	7392877_1	24.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=7392877_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:30819339(-)-23:30820351(+)__23_30796501_30821501D;SPAN=1012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:94 GQ:24.2 PL:[24.2, 0.0, 202.4] SR:0 DR:15 LR:-24.05 LO:32.36);ALT=]chrX:30820351]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	31196943	+	chrX	31216211	+	ATGTAGTG	22	18	7393158_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATGTAGTG;MAPQ=60;MATEID=7393158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_31213001_31238001_3C;SPAN=19268;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:23 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:18 DR:22 LR:-95.72 LO:95.72);ALT=A[chrX:31216211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	31301203	+	chrX	32038750	+	TATTCATTATTATAA	0	11	7393554_1	31.0	.	EVDNC=ASSMB;INSERTION=TATTCATTATTATAA;MAPQ=60;MATEID=7393554_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_32021501_32046501_8C;SPAN=737547;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:17 GQ:8.6 PL:[31.7, 0.0, 8.6] SR:11 DR:0 LR:-32.36 LO:32.36);ALT=T[chrX:32038750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	32077855	+	chrX	32293097	+	GGC	27	14	7393730_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GGC;MAPQ=60;MATEID=7393730_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_32291001_32316001_251C;SPAN=215242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:18 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:14 DR:27 LR:-102.3 LO:102.3);ALT=G[chrX:32293097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	32098533	+	chrX	32201251	+	.	26	10	7393663_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=7393663_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_32193001_32218001_67C;SPAN=102718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:6 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:10 DR:26 LR:-85.82 LO:85.82);ALT=A[chrX:32201251[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
