chr3	167438062	+	chr3	167452594	+	.	30	3	1774070_1	71.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1774070_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_167433001_167458001_250C;SPAN=14532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:101 GQ:71.9 PL:[71.9, 0.0, 170.9] SR:3 DR:30 LR:-71.67 LO:74.0);ALT=C[chr3:167452594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	167565014	-	chr3	167566215	+	.	8	0	1774457_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1774457_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:167565014(-)-3:167566215(-)__3_167555501_167580501D;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr3:167566215[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
