chr3	109103303	+	chr3	109104947	+	.	64	59	2232375_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCT;MAPQ=60;MATEID=2232375_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_109098501_109123501_294C;SPAN=1644;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:94 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:59 DR:64 LR:-310.3 LO:310.3);ALT=T[chr3:109104947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
