chr16	14741501	-	chr16	14742739	+	.	8	0	9164682_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=9164682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:14741501(-)-16:14742739(-)__16_14724501_14749501D;SPAN=1238;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.374 LO:14.01);ALT=[chr16:14742739[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	14905998	+	chr21	42239025	+	.	0	35	10795665_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGAGAGAGAGAGAGAGA;MAPQ=60;MATEID=10795665_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_42238001_42263001_77C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:14 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:35 DR:0 LR:-102.3 LO:102.3);ALT=A[chr21:42239025[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
