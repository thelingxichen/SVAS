chr5	7917050	+	chr5	7920555	+	.	102	83	3187966_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAC;MAPQ=60;MATEID=3187966_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_7913501_7938501_260C;SPAN=3505;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:157 DP:90 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:83 DR:102 LR:-465.4 LO:465.4);ALT=C[chr5:7920555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
