chr9	17945740	+	chr9	17925734	+	.	14	0	5793379_1	37.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=5793379_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:17925734(-)-9:17945740(+)__9_17909501_17934501D;SPAN=20006;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:33 GQ:37.4 PL:[37.4, 0.0, 40.7] SR:0 DR:14 LR:-37.27 LO:37.3);ALT=]chr9:17945740]G;VARTYPE=BND:DUP-th;JOINTYPE=th
