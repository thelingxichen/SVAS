chr8	107681249	+	chr8	107581244	+	.	11	0	5605510_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5605510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:107581244(-)-8:107681249(+)__8_107579501_107604501D;SPAN=100005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=]chr8:107681249]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	108491567	+	chr8	108472574	+	.	56	49	5608735_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=5608735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_108486001_108511001_57C;SPAN=18993;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:79 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:49 DR:56 LR:-250.9 LO:250.9);ALT=]chr8:108491567]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	108504819	+	chr8	108506364	+	.	65	62	5608812_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5608812_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_108486001_108511001_358C;SPAN=1545;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:109 GQ:22.8 PL:[310.2, 22.8, 0.0] SR:62 DR:65 LR:-312.5 LO:312.5);ALT=C[chr8:108506364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
