chr16	72127950	+	chr16	72130036	+	.	14	4	6246081_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6246081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_72128001_72153001_124C;SPAN=2086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:37 GQ:36.2 PL:[36.2, 0.0, 52.7] SR:4 DR:14 LR:-36.19 LO:36.38);ALT=G[chr16:72130036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
