chr6	35626434	+	chr6	35629745	+	.	126	97	4134755_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4134755_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35623001_35648001_349C;SPAN=3311;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:184 DP:36 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:97 DR:126 LR:-544.6 LO:544.6);ALT=G[chr6:35629745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35917093	-	chr6	35918108	+	.	8	0	4136987_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4136987_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:35917093(-)-6:35918108(-)__6_35917001_35942001D;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:125 GQ:7.2 PL:[0.0, 7.2, 316.8] SR:0 DR:8 LR:7.458 LO:13.9);ALT=[chr6:35918108[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
