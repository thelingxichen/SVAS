chr2	55711875	-	chr2	55712985	+	.	8	1	1011437_1	14.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=30;MATEID=1011437_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_55713001_55738001_317C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:1 DR:8 LR:-14.54 LO:19.45);ALT=[chr2:55712985[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	56009777	+	chr2	56011055	-	.	10	0	1013951_1	0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=1013951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:56009777(+)-2:56011055(+)__2_56007001_56032001D;SPAN=1278;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:130 GQ:2.1 PL:[0.0, 2.1, 320.1] SR:0 DR:10 LR:2.21 LO:18.2);ALT=A]chr2:56011055];VARTYPE=BND:INV-hh;JOINTYPE=hh
