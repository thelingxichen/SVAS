chr7	110290537	+	chr7	110273899	+	.	2	3	3522312_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGAA;MAPQ=60;MATEID=3522312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_110274501_110299501_422C;SPAN=16638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:40 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:3 DR:2 LR:-5.668 LO:10.21);ALT=]chr7:110290537]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	110393332	+	chr7	110394461	+	.	27	22	3522596_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3522596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_110372501_110397501_32C;SPAN=1129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:71 GQ:53.6 PL:[116.3, 0.0, 53.6] SR:22 DR:27 LR:-117.2 LO:117.2);ALT=T[chr7:110394461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	111127442	+	chr7	111201933	+	.	11	0	3524733_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3524733_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:111127442(+)-7:111201933(-)__7_111181001_111206001D;SPAN=74491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:69 GQ:17.6 PL:[17.6, 0.0, 149.6] SR:0 DR:11 LR:-17.62 LO:23.72);ALT=C[chr7:111201933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	111161527	+	chr7	111201930	+	.	16	0	3524735_1	34.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3524735_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:111161527(+)-7:111201930(-)__7_111181001_111206001D;SPAN=40403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:67 GQ:34.7 PL:[34.7, 0.0, 127.1] SR:0 DR:16 LR:-34.66 LO:37.67);ALT=C[chr7:111201930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	111846862	+	chr7	111926927	+	.	21	4	3527430_1	60.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3527430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_111916001_111941001_259C;SPAN=80065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:56 GQ:60.8 PL:[60.8, 0.0, 74.0] SR:4 DR:21 LR:-60.75 LO:60.84);ALT=G[chr7:111926927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	112090839	+	chr7	112095816	+	.	0	7	3527965_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=3527965_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_112087501_112112501_289C;SPAN=4977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:100 GQ:3.9 PL:[0.0, 3.9, 250.8] SR:7 DR:0 LR:3.985 LO:12.44);ALT=T[chr7:112095816[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
