chr4	111792671	+	chr4	112242413	+	.	12	50	2148880_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=27;MATEID=2148880_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_112234501_112259501_180C;SPAN=449742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:37 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:50 DR:12 LR:-158.4 LO:158.4);ALT=C[chr4:112242413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	112237555	+	chr4	112242412	+	.	13	0	2148889_1	25.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2148889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:112237555(+)-4:112242412(-)__4_112234501_112259501D;SPAN=4857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:64 GQ:25.7 PL:[25.7, 0.0, 128.0] SR:0 DR:13 LR:-25.57 LO:29.56);ALT=T[chr4:112242412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	112816036	+	chr4	112258296	+	.	45	0	2148948_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2148948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:112258296(-)-4:112816036(+)__4_112234501_112259501D;SPAN=557740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:55 GQ:1.5 PL:[135.3, 1.5, 0.0] SR:0 DR:45 LR:-142.0 LO:142.0);ALT=]chr4:112816036]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	113088071	+	chr4	113471139	+	.	9	0	2151559_1	16.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2151559_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:113088071(+)-4:113471139(-)__4_113067501_113092501D;SPAN=383068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=C[chr4:113471139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	113471279	+	chr4	113088203	+	.	10	0	2151561_1	13.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=2151561_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:113088203(-)-4:113471279(+)__4_113067501_113092501D;SPAN=383076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:0 DR:10 LR:-12.96 LO:20.79);ALT=]chr4:113471279]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	113129342	+	chr10	17058115	-	.	13	0	4528177_1	34.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=4528177_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:113129342(+)-10:17058115(+)__10_17052001_17077001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:33 GQ:34.1 PL:[34.1, 0.0, 44.0] SR:0 DR:13 LR:-33.97 LO:34.07);ALT=C]chr10:17058115];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	113199593	+	chr4	113206794	+	.	0	12	2151609_1	7.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=2151609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_113190001_113215001_25C;SPAN=7201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:118 GQ:7.7 PL:[7.7, 0.0, 278.3] SR:12 DR:0 LR:-7.643 LO:23.36);ALT=G[chr4:113206794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	113558786	+	chr4	113565832	+	.	9	0	2152952_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2152952_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:113558786(+)-4:113565832(-)__4_113557501_113582501D;SPAN=7046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=A[chr4:113565832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	113566027	+	chr4	113567507	+	.	4	8	2152978_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2152978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_113557501_113582501_308C;SPAN=1480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:8 DR:4 LR:-9.44 LO:20.03);ALT=T[chr4:113567507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	113571739	+	chr4	113574232	+	.	3	2	2153004_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2153004_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_113557501_113582501_183C;SPAN=2493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:94 GQ:8.7 PL:[0.0, 8.7, 244.2] SR:2 DR:3 LR:8.962 LO:8.273);ALT=G[chr4:113574232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	16454895	+	chrX	5708272	+	.	14	0	7356933_1	39.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=7356933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:16454895(+)-23:5708272(-)__23_5708501_5733501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:0 GQ:3.6 PL:[39.6, 3.6, 0.0] SR:0 DR:14 LR:-39.61 LO:39.61);ALT=A[chrX:5708272[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	16796989	+	chr10	16806389	+	.	0	10	4527620_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4527620_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_10_16856001_16881001_84C;SPAN=9400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:0 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:10 DR:0 LR:-29.71 LO:29.71);ALT=C[chr10:16806389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	16806550	+	chr10	16859338	+	.	19	0	4527623_1	46.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4527623_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:16806550(+)-10:16859338(-)__10_16856001_16881001D;SPAN=52788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:59 GQ:46.7 PL:[46.7, 0.0, 96.2] SR:0 DR:19 LR:-46.73 LO:47.68);ALT=A[chr10:16859338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	16824132	+	chr10	16859339	+	.	9	0	4527519_1	19.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=4527519_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:16824132(+)-10:16859339(-)__10_16807001_16832001D;SPAN=35207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:0 DR:9 LR:-19.68 LO:21.27);ALT=T[chr10:16859339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17216661	+	chr10	17243570	+	.	8	4	4528603_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4528603_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_17199001_17224001_203C;SPAN=26909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:29 GQ:25.1 PL:[25.1, 0.0, 44.9] SR:4 DR:8 LR:-25.15 LO:25.47);ALT=T[chr10:17243570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17271984	+	chr10	17275584	+	ATTGCAGGAGGAGATGCTTCAGAGAGAGGAAGCCGAAAACACCCTGCAATCTTTCAGAC	47	83	4529011_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTGCAGGAGGAGATGCTTCAGAGAGAGGAAGCCGAAAACACCCTGCAATCTTTCAGAC;MAPQ=60;MATEID=4529011_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_17272501_17297501_71C;SPAN=3600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:63 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:83 DR:47 LR:-323.5 LO:323.5);ALT=A[chr10:17275584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17272759	+	chr10	17275766	+	.	21	0	4529017_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4529017_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:17272759(+)-10:17275766(-)__10_17272501_17297501D;SPAN=3007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:108 GQ:40.1 PL:[40.1, 0.0, 221.6] SR:0 DR:21 LR:-40.06 LO:47.3);ALT=A[chr10:17275766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17275930	+	chr10	17277168	+	TTTGCTGACCTCTCTGAGGCTGCCAACCGGAACAATGACGCCCTGCGCCAGGCAAAGCAGGAGTCCACTGAGTACCGGAGACAGGTGCAGTCCCTCACCTGTGAAGTGGATGCCCTTAAAGGAACC	0	103	4529034_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTTGCTGACCTCTCTGAGGCTGCCAACCGGAACAATGACGCCCTGCGCCAGGCAAAGCAGGAGTCCACTGAGTACCGGAGACAGGTGCAGTCCCTCACCTGTGAAGTGGATGCCCTTAAAGGAACC;MAPQ=60;MATEID=4529034_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_17272501_17297501_271C;SPAN=1238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:103 DP:179 GQ:99 PL:[291.5, 0.0, 143.0] SR:103 DR:0 LR:-294.3 LO:294.3);ALT=G[chr10:17277168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17277430	+	chr10	17279224	+	.	14	0	4529045_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4529045_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:17277430(+)-10:17279224(-)__10_17272501_17297501D;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:14 DP:211 GQ:10.6 PL:[0.0, 10.6, 531.4] SR:0 DR:14 LR:10.95 LO:24.55);ALT=T[chr10:17279224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17582925	+	chr10	17627107	+	.	12	0	4529753_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4529753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:17582925(+)-10:17627107(-)__10_17615501_17640501D;SPAN=44182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=G[chr10:17627107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17595895	+	chr10	17627103	+	.	4	2	4529756_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4529756_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_17615501_17640501_3C;SPAN=31208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:37 GQ:3.2 PL:[3.2, 0.0, 85.7] SR:2 DR:4 LR:-3.18 LO:7.9);ALT=T[chr10:17627103[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	17604764	+	chr10	17627112	+	.	8	0	4529757_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4529757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:17604764(+)-10:17627112(-)__10_17615501_17640501D;SPAN=22348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=A[chr10:17627112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	5729125	-	chrX	5730607	+	.	32	37	7356970_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTGGA;MAPQ=60;MATEID=7356970_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_5708501_5733501_80C;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:61 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:37 DR:32 LR:-184.8 LO:184.8);ALT=[chrX:5730607[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	5729126	+	chrX	5730792	-	.	22	42	7356971_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=7356971_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_5708501_5733501_122C;SPAN=1666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:61 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:42 DR:22 LR:-178.2 LO:178.2);ALT=T]chrX:5730792];VARTYPE=BND:INV-hh;JOINTYPE=hh
