chr22	27168076	+	chr22	27169793	+	.	62	49	10860934_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTAACCTCT;MAPQ=60;MATEID=10860934_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_22_27146001_27171001_65C;SPAN=1717;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:17 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:49 DR:62 LR:-244.3 LO:244.3);ALT=T[chr22:27169793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
