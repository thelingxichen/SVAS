chr16	58007178	-	chr16	58008400	+	.	8	0	9342349_1	0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=9342349_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:58007178(-)-16:58008400(-)__16_57991501_58016501D;SPAN=1222;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:163 GQ:17.5 PL:[0.0, 17.5, 429.1] SR:0 DR:8 LR:17.75 LO:12.95);ALT=[chr16:58008400[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
