chr6	151485910	+	chr6	151486940	+	.	28	0	3075447_1	76.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3075447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:151485910(+)-6:151486940(-)__6_151483501_151508501D;SPAN=1030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:59 GQ:66.5 PL:[76.4, 0.0, 66.5] SR:0 DR:28 LR:-76.48 LO:76.48);ALT=T[chr6:151486940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
