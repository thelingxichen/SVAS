chr7	151010035	-	chr7	151012106	+	.	32	48	5327745_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=5327745_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_150993501_151018501_252C;SPAN=2071;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:77 DP:259 GQ:99 PL:[184.0, 0.0, 444.8] SR:48 DR:32 LR:-184.0 LO:190.0);ALT=[chr7:151012106[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
