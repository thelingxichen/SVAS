chr1	84517939	+	chr1	84524630	+	.	63	44	389401_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGATTTGTTTTTCT;MAPQ=60;MATEID=389401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84525001_84550001_26C;SPAN=6691;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:0 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:44 DR:63 LR:-257.5 LO:257.5);ALT=T[chr1:84524630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84712005	+	chr1	84715875	+	GTGCACAAT	0	52	390533_1	99.0	.	EVDNC=ASSMB;INSERTION=GTGCACAAT;MAPQ=60;MATEID=390533_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84696501_84721501_41C;SPAN=3870;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:85 GQ:56.3 PL:[148.7, 0.0, 56.3] SR:52 DR:0 LR:-150.8 LO:150.8);ALT=T[chr1:84715875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84756829	-	chr1	84758982	+	.	10	0	389960_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=389960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:84756829(-)-1:84758982(-)__1_84745501_84770501D;SPAN=2153;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:176 GQ:14.5 PL:[0.0, 14.5, 455.5] SR:0 DR:10 LR:14.67 LO:16.84);ALT=[chr1:84758982[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
