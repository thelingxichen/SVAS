chr2	91751062	+	chr2	91759767	+	.	94	28	894272_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=19;MATEID=894272_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_91728001_91753001_466C;SPAN=8705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:100 GQ:30 PL:[330.0, 30.0, 0.0] SR:28 DR:94 LR:-330.1 LO:330.1);ALT=T[chr2:91759767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	92276743	+	chr2	92280093	+	.	22	0	899882_1	45.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=899882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:92276743(+)-2:92280093(-)__2_92267001_92292001D;SPAN=3350;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:101 GQ:45.5 PL:[45.5, 0.0, 197.3] SR:0 DR:22 LR:-45.26 LO:50.79);ALT=A[chr2:92280093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	92285674	+	chr2	92289070	+	.	12	0	899927_1	20.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=899927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:92285674(+)-2:92289070(-)__2_92267001_92292001D;SPAN=3396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:70 GQ:20.6 PL:[20.6, 0.0, 149.3] SR:0 DR:12 LR:-20.65 LO:26.3);ALT=A[chr2:92289070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
