chr2	8967273	+	chr2	8977667	+	.	9	0	681202_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=681202_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:8967273(+)-2:8977667(-)__2_8967001_8992001D;SPAN=10394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:0 DR:9 LR:-6.139 LO:17.59);ALT=C[chr2:8977667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9552538	+	chr2	9558755	+	GCTTTTGGTGGAATCTGTGTCGAGGCTGGCCACAGTGCTGGATCGTGAAAGACCCCCAAGGCTAGAATCCACAGA	0	34	682768_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GCTTTTGGTGGAATCTGTGTCGAGGCTGGCCACAGTGCTGGATCGTGAAAGACCCCCAAGGCTAGAATCCACAGA;MAPQ=60;MATEID=682768_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_9555001_9580001_234C;SPAN=6217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:34 DR:0 LR:-110.1 LO:110.1);ALT=A[chr2:9558755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9552538	+	chr2	9554306	+	.	0	8	682746_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCTGA;MAPQ=60;MATEID=682746_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_9530501_9555501_202C;SPAN=1768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-2.025 LO:15.08);ALT=A[chr2:9554306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9552573	+	chr2	9563500	+	.	9	0	682769_1	21.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=682769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:9552573(+)-2:9563500(-)__2_9555001_9580001D;SPAN=10927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.31 LO:22.09);ALT=T[chr2:9563500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9554430	+	chr2	9563500	+	.	13	0	682771_1	34.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=682771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:9554430(+)-2:9563500(-)__2_9555001_9580001D;SPAN=9070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:31 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:0 DR:13 LR:-34.51 LO:34.54);ALT=C[chr2:9563500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9558863	+	chr2	9563501	+	.	25	18	682786_1	84.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=682786_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9555001_9580001_207C;SPAN=4638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:67 GQ:77.6 PL:[84.2, 0.0, 77.6] SR:18 DR:25 LR:-84.19 LO:84.19);ALT=T[chr2:9563501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9568957	+	chr2	9570051	+	.	0	4	682817_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=682817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9555001_9580001_84C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:4 DR:0 LR:6.844 LO:6.647);ALT=G[chr2:9570051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9607906	+	chr2	9611472	+	.	2	7	682867_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=682867_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9604001_9629001_97C;SPAN=3566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:7 DR:2 LR:-0.6203 LO:13.03);ALT=G[chr2:9611472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9611568	+	chr2	9613044	+	.	0	9	682877_1	5.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=682877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9604001_9629001_87C;SPAN=1476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:9 DR:0 LR:-5.868 LO:17.54);ALT=G[chr2:9613044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9614774	+	chr2	9621411	+	.	13	0	682886_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=682886_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:9614774(+)-2:9621411(-)__2_9604001_9629001D;SPAN=6637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:70 GQ:23.9 PL:[23.9, 0.0, 146.0] SR:0 DR:13 LR:-23.95 LO:28.99);ALT=C[chr2:9621411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9614776	+	chr2	9616112	+	.	6	6	682887_1	11.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=CCAG;MAPQ=60;MATEID=682887_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_2_9604001_9629001_200C;SPAN=1336;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:6 DR:6 LR:-10.97 LO:16.77);ALT=G[chr2:9616112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9614776	+	chr2	9618348	+	.	74	4	682889_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=682889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9604001_9629001_117C;SPAN=3572;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:63 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:4 DR:74 LR:-221.2 LO:221.2);ALT=G[chr2:9618348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9618499	+	chr2	9621413	+	.	0	36	682899_1	95.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=682899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9604001_9629001_103C;SPAN=2914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:86 GQ:95.6 PL:[95.6, 0.0, 112.1] SR:36 DR:0 LR:-95.54 LO:95.62);ALT=G[chr2:9621413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9624680	+	chr2	9628274	+	.	3	4	682906_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=682906_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9604001_9629001_64C;SPAN=3594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:4 DR:3 LR:-3.059 LO:13.4);ALT=G[chr2:9628274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9728457	+	chr2	9731521	+	.	4	3	683413_1	0	.	DISC_MAPQ=54;EVDNC=ASDIS;MAPQ=60;MATEID=683413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9726501_9751501_131C;SPAN=3064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:81 GQ:1.8 PL:[0.0, 1.8, 198.0] SR:3 DR:4 LR:2.139 LO:10.82);ALT=T[chr2:9731521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	9731645	+	chr2	9770287	+	.	5	11	683418_1	38.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=683418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_9726501_9751501_193C;SPAN=38642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:30 GQ:34.7 PL:[38.0, 0.0, 34.7] SR:11 DR:5 LR:-38.09 LO:38.09);ALT=C[chr2:9770287[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10443193	+	chr2	10536957	+	.	12	0	685809_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=685809_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:10443193(+)-2:10536957(-)__2_10535001_10560001D;SPAN=93764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=C[chr2:10536957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10585392	+	chr2	10588247	+	.	27	20	685894_1	94.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=685894_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_10584001_10609001_3C;SPAN=2855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:77 GQ:91.4 PL:[94.7, 0.0, 91.4] SR:20 DR:27 LR:-94.68 LO:94.68);ALT=T[chr2:10588247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10925158	+	chr2	10927406	+	.	6	4	687286_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=687286_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_10927001_10952001_335C;SPAN=2248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:40 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:4 DR:6 LR:-22.17 LO:23.78);ALT=T[chr2:10927406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10927566	+	chr2	10928821	+	.	3	9	687288_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=687288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_10927001_10952001_35C;SPAN=1255;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:95 GQ:14 PL:[14.0, 0.0, 215.3] SR:9 DR:3 LR:-13.87 LO:24.56);ALT=C[chr2:10928821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10930016	+	chr2	10931921	+	CCGTATCGGGAGGCCAGAACCTGATTGACTGTAGCATCCACAGCTGCCAGTTTCACTTTTCCTTTCGTCTGCTCTTTTACTTCTGAAGCTGCGGCAGCCCACTCTGGCTCTAGG	0	13	687310_1	18.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCGTATCGGGAGGCCAGAACCTGATTGACTGTAGCATCCACAGCTGCCAGTTTCACTTTTCCTTTCGTCTGCTCTTTTACTTCTGAAGCTGCGGCAGCCCACTCTGGCTCTAGG;MAPQ=60;MATEID=687310_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_10927001_10952001_86C;SPAN=1905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:13 DR:0 LR:-18.53 LO:27.43);ALT=C[chr2:10931921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10932051	+	chr2	10933221	+	.	3	6	687321_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=687321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_10927001_10952001_77C;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:90 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:6 DR:3 LR:1.276 LO:12.77);ALT=C[chr2:10933221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10933330	+	chr2	10952802	+	TGGTAATCTTCTGGTCTGTTTTTGTTGGATCCAAAAATCTTAATGGTAGGAAATCCCTGAACACCATACTGACCTCCTAGGGAATGATGCTTATCTGCATCAACTGCACCAACTTTGACAACATCTTTTAATGCAGTTGCTGCTTTCTTCCATTCTGGTGTTAATCTTTGACAGTGACCACACCATGGAGCATAGAATTCTACAAGCCACAAACTATCACTCTGAATAACTTCTCGGTTGAAATTCGATGGAGTTAATTCGATCACATCATCACTAGAGGAATACAGACCATTCACTGCCAGAAAGAAGGTACAGCTCACCAG	0	34	687325_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TGGTAATCTTCTGGTCTGTTTTTGTTGGATCCAAAAATCTTAATGGTAGGAAATCCCTGAACACCATACTGACCTCCTAGGGAATGATGCTTATCTGCATCAACTGCACCAACTTTGACAACATCTTTTAATGCAGTTGCTGCTTTCTTCCATTCTGGTGTTAATCTTTGACAGTGACCACACCATGGAGCATAGAATTCTACAAGCCACAAACTATCACTCTGAATAACTTCTCGGTTGAAATTCGATGGAGTTAATTCGATCACATCATCACTAGAGGAATACAGACCATTCACTGCCAGAAAGAAGGTACAGCTCACCAG;MAPQ=60;MATEID=687325_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_2_10927001_10952001_132C;SPAN=19472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:30 GQ:9 PL:[99.0, 9.0, 0.0] SR:34 DR:0 LR:-99.02 LO:99.02);ALT=T[chr2:10952802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10933330	+	chr2	10937205	+	.	4	5	687324_1	8.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=687324_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GG;SCTG=c_2_10927001_10952001_132C;SPAN=3875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:5 DR:4 LR:-8.798 LO:16.28);ALT=T[chr2:10937205[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10937884	+	chr2	10942623	+	.	5	64	687336_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=687336_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=CC;SCTG=c_2_10927001_10952001_132C;SPAN=4739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:97 GQ:36.5 PL:[198.2, 0.0, 36.5] SR:64 DR:5 LR:-204.4 LO:204.4);ALT=C[chr2:10942623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10937931	+	chr2	10952801	+	.	47	0	687337_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=687337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:10937931(+)-2:10952801(-)__2_10927001_10952001D;SPAN=14870;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:35 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=C[chr2:10952801[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	10942767	+	chr2	10952802	+	.	88	24	687370_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=687370_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=CC;SCTG=c_2_10927001_10952001_132C;SPAN=10035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:41 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:24 DR:88 LR:-283.9 LO:283.9);ALT=C[chr2:10952802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	11295815	+	chr2	11300591	+	.	41	26	688250_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=688250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_11294501_11319501_32C;SPAN=4776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:85 GQ:53 PL:[152.0, 0.0, 53.0] SR:26 DR:41 LR:-154.5 LO:154.5);ALT=G[chr2:11300591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	11886849	+	chr2	11905692	+	.	15	0	689906_1	28.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=689906_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:11886849(+)-2:11905692(-)__2_11882501_11907501D;SPAN=18843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:77 GQ:28.7 PL:[28.7, 0.0, 157.4] SR:0 DR:15 LR:-28.65 LO:33.8);ALT=C[chr2:11905692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	11905861	+	chr2	11907888	+	.	0	13	689963_1	29.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=689963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_11882501_11907501_346C;SPAN=2027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:48 GQ:29.9 PL:[29.9, 0.0, 86.0] SR:13 DR:0 LR:-29.91 LO:31.44);ALT=T[chr2:11907888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	11922633	+	chr2	11923953	+	.	3	3	690148_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=690148_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_11907001_11932001_349C;SPAN=1320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:69 GQ:5.4 PL:[0.0, 5.4, 178.2] SR:3 DR:3 LR:5.49 LO:6.772);ALT=G[chr2:11923953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	11929912	-	chr4	162053660	+	.	20	0	2304400_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2304400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:11929912(-)-4:162053660(-)__4_162043001_162068001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:16 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:20 LR:-59.41 LO:59.41);ALT=[chr4:162053660[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	11930018	+	chr4	162053250	-	ATAAAT	12	25	2304401_1	95.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=ATAAAT;MAPQ=60;MATEID=2304401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_162043001_162068001_361C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:31 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:25 DR:12 LR:-95.72 LO:95.72);ALT=G]chr4:162053250];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	162054302	+	chr4	162063311	+	ATT	66	53	2304428_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=ATT;MAPQ=60;MATEID=2304428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_162043001_162068001_54C;SPAN=9009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:69 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:53 DR:66 LR:-310.3 LO:310.3);ALT=A[chr4:162063311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	162449277	+	chr4	162451667	+	.	39	49	2305723_1	99.0	.	DISC_MAPQ=14;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=56;MATEID=2305723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_162435001_162460001_320C;SPAN=2390;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:25 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:49 DR:39 LR:-221.2 LO:221.2);ALT=T[chr4:162451667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
