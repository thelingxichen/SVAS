chr4	35146799	+	chr4	35152239	+	.	41	19	1938212_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=1938212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_35133001_35158001_65C;SPAN=5440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:41 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:19 DR:41 LR:-151.8 LO:151.8);ALT=G[chr4:35152239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
