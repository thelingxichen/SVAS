chr6	170104186	+	chr6	170105227	+	.	0	4	3122664_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3122664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_170103501_170128501_222C;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:84 GQ:9.3 PL:[0.0, 9.3, 221.1] SR:4 DR:0 LR:9.554 LO:6.423);ALT=T[chr6:170105227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170484770	+	chr6	170483704	+	.	37	0	3124018_1	95.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=3124018_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:170483704(-)-6:170484770(+)__6_170471001_170496001D;SPAN=1066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:98 GQ:95.6 PL:[95.6, 0.0, 141.8] SR:0 DR:37 LR:-95.59 LO:96.09);ALT=]chr6:170484770]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	170485162	+	chr6	170486284	+	.	0	5	3124046_1	0	.	EVDNC=ASSMB;HOMSEQ=CTGTTCGGGGTTGTTCC;MAPQ=60;MATEID=3124046_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_170471001_170496001_293C;SPAN=1122;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:196 GQ:36.4 PL:[0.0, 36.4, 547.9] SR:5 DR:0 LR:36.6 LO:6.663);ALT=C[chr6:170486284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170844498	+	chr6	170846320	+	.	5	36	3124876_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTGGT;MAPQ=60;MATEID=3124876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_170838501_170863501_123C;SPAN=1822;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:101 GQ:99 PL:[104.9, 0.0, 137.9] SR:36 DR:5 LR:-104.7 LO:105.0);ALT=T[chr6:170846320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170846431	+	chr6	170852688	+	.	0	10	3124882_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CCTT;MAPQ=60;MATEID=3124882_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_170838501_170863501_334C;SPAN=6257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:10 DR:0 LR:-10.52 LO:20.25);ALT=T[chr6:170852688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170852820	+	chr6	170855191	+	.	6	34	3124895_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3124895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_170838501_170863501_204C;SPAN=2371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:100 GQ:99 PL:[101.6, 0.0, 141.2] SR:34 DR:6 LR:-101.6 LO:102.0);ALT=T[chr6:170855191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170852859	+	chr6	170862273	+	.	11	0	3124897_1	1.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3124897_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:170852859(+)-6:170862273(-)__6_170838501_170863501D;SPAN=9414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:131 GQ:1.1 PL:[1.1, 0.0, 314.6] SR:0 DR:11 LR:-0.8199 LO:20.45);ALT=G[chr6:170862273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170855272	+	chr6	170862218	+	AATTTGTAACATTTGGGGCTATCCCGCGTATGAATTGAAAACCCTTCACTCAATCGAGTATCAGAAGCAACAATTGCAAAATCTTCTCCAGCAATTGCCAGTATAGTA	53	159	3124903_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AATTTGTAACATTTGGGGCTATCCCGCGTATGAATTGAAAACCCTTCACTCAATCGAGTATCAGAAGCAACAATTGCAAAATCTTCTCCAGCAATTGCCAGTATAGTA;MAPQ=60;MATEID=3124903_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_170838501_170863501_79C;SPAN=6946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:178 DP:127 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:159 DR:53 LR:-528.1 LO:528.1);ALT=T[chr6:170862218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170858202	+	chr6	170862218	+	.	104	86	3124913_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3124913_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_170838501_170863501_79C;SPAN=4016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:149 DP:128 GQ:40.3 PL:[442.3, 40.3, 0.0] SR:86 DR:104 LR:-442.3 LO:442.3);ALT=C[chr6:170862218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	170886808	+	chr6	170887943	+	.	0	5	3124789_1	5.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=3124789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_170887501_170912501_298C;SPAN=1135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:41 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:5 DR:0 LR:-5.397 LO:10.15);ALT=G[chr6:170887943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
