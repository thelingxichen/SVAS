chr2	91679897	+	chr2	91685489	+	TGTAGAAAGCCCAGG	49	110	1168374_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;INSERTION=TGTAGAAAGCCCAGG;MAPQ=26;MATEID=1168374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_91679001_91704001_309C;SPAN=5592;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:139 DP:277 GQ:99 PL:[383.9, 0.0, 288.1] SR:110 DR:49 LR:-384.5 LO:384.5);ALT=C[chr2:91685489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	92115622	-	chr2	92119864	+	.	10	0	1175051_1	0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=1175051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:92115622(-)-2:92119864(-)__2_92095501_92120501D;SPAN=4242;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:122 GQ:0.2 PL:[0.2, 0.0, 293.9] SR:0 DR:10 LR:0.04279 LO:18.48);ALT=[chr2:92119864[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	92120521	+	chr2	92126609	-	.	53	0	1175087_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=1175087_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:92120521(+)-2:92126609(+)__2_92095501_92120501D;SPAN=6088;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:34 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:0 DR:53 LR:-155.1 LO:155.1);ALT=T]chr2:92126609];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	92120521	-	chr2	92135983	+	.	28	42	1174353_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=1174353_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_2_92120001_92145001_198C;SECONDARY;SPAN=15462;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:88 GQ:29 PL:[184.1, 0.0, 29.0] SR:42 DR:28 LR:-190.5 LO:190.5);ALT=[chr2:92135983[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
