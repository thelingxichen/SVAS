chr17	39790038	+	chr17	39788816	+	.	10	0	9647706_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=9647706_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:39788816(-)-17:39790038(+)__17_39788001_39813001D;SPAN=1222;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:307 GQ:50 PL:[0.0, 50.0, 845.0] SR:0 DR:10 LR:50.16 LO:14.39);ALT=]chr17:39790038]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	39959032	+	chr17	39960688	-	.	15	3	9648345_1	47.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CCAGGCTGGTCTTGAACTCCTG;MAPQ=60;MATEID=9648345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_39959501_39984501_1C;SPAN=1656;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:44 GQ:47.6 PL:[47.6, 0.0, 57.5] SR:3 DR:15 LR:-47.5 LO:47.57);ALT=G]chr17:39960688];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	39959094	+	chr17	39960451	+	.	83	49	9648346_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CCTTGGCCTCCCAAAATGCTGGGATTACAGGTGTGAGCCACCG;MAPQ=60;MATEID=9648346_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_39959501_39984501_224C;SPAN=1357;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:124 DP:11 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:49 DR:83 LR:-366.4 LO:366.4);ALT=G[chr17:39960451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
