chr6	34271817	-	chr6	34272975	+	.	3	3	4128485_1	0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=TCTCGAACTCCTGAC;MAPQ=60;MATEID=4128485_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_34251001_34276001_437C;SPAN=1158;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:133 GQ:19.2 PL:[0.0, 19.2, 359.7] SR:3 DR:3 LR:19.53 LO:7.508);ALT=[chr6:34272975[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
