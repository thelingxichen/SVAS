chr17	72729558	+	chr17	72724024	+	.	10	0	9809761_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=9809761_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:72724024(-)-17:72729558(+)__17_72716001_72741001D;SPAN=5534;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:299 GQ:47.9 PL:[0.0, 47.9, 821.9] SR:0 DR:10 LR:48.0 LO:14.5);ALT=]chr17:72729558]T;VARTYPE=BND:DUP-th;JOINTYPE=th
