chr12	108862531	+	chr1	6037971	+	.	8	0	30950_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=30950_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6037971(-)-12:108862531(+)__1_6027001_6052001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:23 GQ:20.3 PL:[20.3, 0.0, 33.5] SR:0 DR:8 LR:-20.18 LO:20.41);ALT=]chr12:108862531]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	6487927	+	chr1	17046951	+	.	0	21	89705_1	30.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=21;MATEID=89705_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17027501_17052501_804C;SPAN=10559024;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:145 GQ:30.2 PL:[30.2, 0.0, 320.6] SR:21 DR:0 LR:-30.04 LO:44.34);ALT=G[chr1:17046951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16151935	+	chr1	16155440	+	GAGGCGGGCCTTCCAAAATA	39	41	82132_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;INSERTION=GAGGCGGGCCTTCCAAAATA;MAPQ=60;MATEID=82132_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_16145501_16170501_444C;SPAN=3505;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:94 GQ:27.5 PL:[199.1, 0.0, 27.5] SR:41 DR:39 LR:-206.3 LO:206.3);ALT=C[chr1:16155440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16376518	+	chr1	16386258	+	.	57	89	83615_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=83615_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_16366001_16391001_170C;SPAN=9740;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:114 DP:112 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:89 DR:57 LR:-336.7 LO:336.7);ALT=T[chr1:16386258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16386334	+	chr1	16376519	+	CACC	0	95	83618_1	99.0	.	EVDNC=ASSMB;INSERTION=CACC;MAPQ=60;MATEID=83618_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_16366001_16391001_275C;SPAN=9815;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:95 DP:124 GQ:19.4 PL:[280.1, 0.0, 19.4] SR:95 DR:0 LR:-293.2 LO:293.2);ALT=]chr1:16386334]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	16942807	+	chr1	149140721	+	CTATATC	2	56	89136_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTATATC;MAPQ=60;MATEID=89136_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_16929501_16954501_423C;SPAN=132197914;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:133 GQ:99 PL:[155.6, 0.0, 165.5] SR:56 DR:2 LR:-155.4 LO:155.5);ALT=T[chr1:149140721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17051748	-	chr1	234912188	+	GCAGAAGCCGGCGGGATGGGGC	212	86	863110_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GCAGAAGCCGGCGGGATGGGGC;MAPQ=60;MATEID=863110_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_234906001_234931001_216C;SPAN=217860440;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:268 DP:91 GQ:72.4 PL:[795.4, 72.4, 0.0] SR:86 DR:212 LR:-795.5 LO:795.5);ALT=[chr1:234912188[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	17216863	-	chr1	149229911	+	.	10	37	530298_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTT;MAPQ=49;MATEID=530298_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_1_149205001_149230001_304C;SPAN=132013048;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:24 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:37 DR:10 LR:-125.4 LO:125.4);ALT=[chr1:149229911[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	144526643	-	chr1	149203979	+	.	8	0	498250_1	0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=498250_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:144526643(-)-1:149203979(-)__1_144525501_144550501D;SPAN=4677336;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:116 GQ:4.8 PL:[0.0, 4.8, 290.4] SR:0 DR:8 LR:5.019 LO:14.16);ALT=[chr1:149203979[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	144896297	+	chr1	144901047	+	GTAACAGG	57	55	499428_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=GTAACAGG;MAPQ=60;MATEID=499428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_144893001_144918001_543C;SPAN=4750;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:94 DP:138 GQ:61.7 PL:[272.9, 0.0, 61.7] SR:55 DR:57 LR:-280.4 LO:280.4);ALT=G[chr1:144901047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	144896341	+	chr1	144906808	+	.	33	0	499429_1	70.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=499429_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:144896341(+)-1:144906808(-)__1_144893001_144918001D;SPAN=10467;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:144 GQ:70.1 PL:[70.1, 0.0, 278.0] SR:0 DR:33 LR:-69.92 LO:77.01);ALT=A[chr1:144906808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	144901180	+	chr1	144906810	+	.	44	45	499448_1	99.0	.	DISC_MAPQ=35;EVDNC=TSI_L;MAPQ=45;MATEID=499448_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_1_144893001_144918001_429C;SPAN=5630;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:162 GQ:99 PL:[203.9, 0.0, 187.4] SR:45 DR:44 LR:-203.7 LO:203.7);ALT=G[chr1:144906810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145067309	+	chr1	145069124	-	.	8	0	502302_1	0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=502302_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:145067309(+)-1:145069124(+)__1_145064501_145089501D;SPAN=1815;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:478 GQ:99 PL:[0.0, 102.9, 1366.0] SR:0 DR:8 LR:103.1 LO:9.211);ALT=G]chr1:145069124];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	145092948	+	chr1	145097095	+	ACCTGTTAAAAG	67	110	500989_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=ACCTGTTAAAAG;MAPQ=60;MATEID=500989_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_145089001_145114001_396C;SPAN=4147;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:164 DP:197 GQ:10.3 PL:[498.4, 10.3, 0.0] SR:110 DR:67 LR:-520.8 LO:520.8);ALT=C[chr1:145097095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145139863	-	chr12	93771888	+	.	38	0	501712_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=501712_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:145139863(-)-12:93771888(-)__1_145138001_145163001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:38 DP:88 GQ:99 PL:[101.6, 0.0, 111.5] SR:0 DR:38 LR:-101.6 LO:101.6);ALT=[chr12:93771888[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	234318646	+	chr1	234319748	+	.	27	27	861032_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=861032_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_234293501_234318501_172C;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:44 DP:0 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:27 DR:27 LR:-128.7 LO:128.7);ALT=A[chr1:234319748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	234607336	+	chr1	234565262	+	.	6	10	861872_1	37.0	.	DISC_MAPQ=43;EVDNC=ASDIS;MAPQ=60;MATEID=861872_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_234587501_234612501_194C;SPAN=42074;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:32 GQ:37.7 PL:[37.7, 0.0, 37.7] SR:10 DR:6 LR:-37.54 LO:37.55);ALT=]chr1:234607336]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	93504293	+	chr12	93505388	+	CCAAATA	72	53	7794589_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCAAATA;MAPQ=60;MATEID=7794589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_93492001_93517001_167C;SPAN=1095;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:23 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:53 DR:72 LR:-293.8 LO:293.8);ALT=A[chr12:93505388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93895672	+	chr12	93894557	+	AAATTAAA	0	47	7795615_1	99.0	.	EVDNC=ASSMB;INSERTION=AAATTAAA;MAPQ=60;MATEID=7795615_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_93884001_93909001_263C;SPAN=1115;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:47 DP:50 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:47 DR:0 LR:-148.5 LO:148.5);ALT=]chr12:93895672]C;VARTYPE=BND:DUP-th;JOINTYPE=th
