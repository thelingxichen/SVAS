chr7	110181968	+	chr7	110188433	+	.	58	39	5130597_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCT;MAPQ=11;MATEID=5130597_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_110176501_110201501_83C;SPAN=6465;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:81 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:39 DR:58 LR:-247.6 LO:247.6);ALT=T[chr7:110188433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	110313150	+	chr7	110608584	+	.	79	28	5131505_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5131505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_110593001_110618001_70C;SPAN=295434;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:45 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:28 DR:79 LR:-267.4 LO:267.4);ALT=C[chr7:110608584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	110650207	+	chr7	110723402	+	.	53	46	5131749_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=5131749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_110715501_110740501_353C;SPAN=73195;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:35 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:46 DR:53 LR:-237.7 LO:237.7);ALT=A[chr7:110723402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
