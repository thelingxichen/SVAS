chr8	137160197	+	chr8	137163899	+	.	43	34	4093886_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=4093886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_137151001_137176001_223C;SPAN=3702;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:68 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:34 DR:43 LR:-201.3 LO:201.3);ALT=C[chr8:137163899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
