chr7	224289	+	chr7	225976	+	.	57	19	4489446_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=GGGGTCGCACGGCGGCTGTCCCCTGAGCCTTCTCTCA;MAPQ=21;MATEID=4489446_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_220501_245501_117C;SPAN=1687;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:55 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:19 DR:57 LR:-221.2 LO:221.2);ALT=A[chr7:225976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	452941	-	chr7	453952	+	.	9	0	4490301_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4490301_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:452941(-)-7:453952(-)__7_441001_466001D;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:112 GQ:0.3 PL:[0.0, 0.3, 270.6] SR:0 DR:9 LR:0.6346 LO:16.56);ALT=[chr7:453952[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	1043202	+	chr7	1041091	+	.	22	0	4493329_1	36.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4493329_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:1041091(-)-7:1043202(+)__7_1029001_1054001D;SPAN=2111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:135 GQ:36.2 PL:[36.2, 0.0, 290.3] SR:0 DR:22 LR:-36.05 LO:47.68);ALT=]chr7:1043202]T;VARTYPE=BND:DUP-th;JOINTYPE=th
