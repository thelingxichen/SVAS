chr4	80360630	+	chr4	80362723	+	.	38	30	2765269_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2765269_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_80335501_80360501_105C;SPAN=2093;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:0 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:30 DR:38 LR:-211.3 LO:211.3);ALT=G[chr4:80362723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	80888062	+	chr4	80894092	+	.	49	27	2766291_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAATAGGGCGTCCG;MAPQ=60;MATEID=2766291_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_80874501_80899501_81C;SPAN=6030;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:69 DP:135 GQ:99 PL:[191.3, 0.0, 135.2] SR:27 DR:49 LR:-191.7 LO:191.7);ALT=G[chr4:80894092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
