chrX	100274978	-	chrX	100276413	+	.	8	0	7483574_1	14.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7483574_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:100274978(-)-23:100276413(-)__23_100254001_100279001D;SPAN=1435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=[chrX:100276413[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	100629623	+	chrX	100641050	+	CCACGTTCAAAGTCATACTCATAGTAGGAGAGTTTGTGCACGGTCAAGAGAAACAGGCGCTTCTTGAAGTTTAGAGGTGATGTTTTCTTTTTCTGTTGGGATCGCTTCAGAAAGATGCTCTCCAGAATCACTGCGGCCATAGCTTCTTCTTTCTGGAGTTCACCTGTGTG	0	32	7484203_1	87.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCACGTTCAAAGTCATACTCATAGTAGGAGAGTTTGTGCACGGTCAAGAGAAACAGGCGCTTCTTGAAGTTTAGAGGTGATGTTTTCTTTTTCTGTTGGGATCGCTTCAGAAAGATGCTCTCCAGAATCACTGCGGCCATAGCTTCTTCTTTCTGGAGTTCACCTGTGTG;MAPQ=60;MATEID=7484203_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_100621501_100646501_43C;SPAN=11427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:68 GQ:77.3 PL:[87.2, 0.0, 77.3] SR:32 DR:0 LR:-87.24 LO:87.24);ALT=C[chrX:100641050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	100630304	+	chrX	100641050	+	.	45	13	7484205_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=7484205_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_100621501_100646501_43C;SPAN=10746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:74 GQ:32.9 PL:[145.1, 0.0, 32.9] SR:13 DR:45 LR:-148.8 LO:148.8);ALT=T[chrX:100641050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	100658977	+	chrX	100662698	+	.	0	23	7484350_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CTGA;MAPQ=60;MATEID=7484350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_100646001_100671001_166C;SPAN=3721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:61 GQ:59.6 PL:[59.6, 0.0, 86.0] SR:23 DR:0 LR:-59.4 LO:59.71);ALT=A[chrX:100662698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	100663307	+	chrX	100666922	+	.	28	5	7484363_1	88.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7484363_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_100646001_100671001_261C;SPAN=3615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:65 GQ:68.3 PL:[88.1, 0.0, 68.3] SR:5 DR:28 LR:-88.13 LO:88.13);ALT=G[chrX:100666922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	100871801	+	chrX	100872872	+	.	25	0	7484578_1	68.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7484578_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:100871801(+)-23:100872872(-)__23_100866501_100891501D;SPAN=1071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:51 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:0 DR:25 LR:-68.79 LO:68.79);ALT=T[chrX:100872872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
