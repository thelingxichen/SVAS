chr12	84593114	+	chr12	84596012	+	.	62	36	5270600_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCCTCA;MAPQ=60;MATEID=5270600_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_84574001_84599001_310C;SPAN=2898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:46 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:36 DR:62 LR:-237.7 LO:237.7);ALT=A[chr12:84596012[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
