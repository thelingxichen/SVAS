chr7	133785003	+	chr7	133798330	+	.	88	59	5290473_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=60;MATEID=5290473_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_133794501_133819501_71C;SPAN=13327;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:118 DP:12 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:59 DR:88 LR:-349.9 LO:349.9);ALT=C[chr7:133798330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
