chr4	61330106	+	chr4	61333187	+	G	56	54	2730827_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=2730827_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_4_61323501_61348501_119C;SPAN=3081;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:18 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:54 DR:56 LR:-303.7 LO:303.7);ALT=T[chr4:61333187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
