chr1	150497311	-	chr1	150498923	+	.	10	0	537312_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=537312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150497311(-)-1:150498923(-)__1_150479001_150504001D;SPAN=1612;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:252 GQ:34.9 PL:[0.0, 34.9, 679.9] SR:0 DR:10 LR:35.26 LO:15.25);ALT=[chr1:150498923[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	150763722	+	chr1	150524662	+	.	46	20	538754_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=538754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150748501_150773501_459C;SPAN=239060;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:57 DP:79 GQ:24.8 PL:[166.7, 0.0, 24.8] SR:20 DR:46 LR:-172.8 LO:172.8);ALT=]chr1:150763722]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	150593722	-	chr5	55447995	+	.	24	41	3437217_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3437217_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_55443501_55468501_178C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:57 DP:89 GQ:51.8 PL:[164.0, 0.0, 51.8] SR:41 DR:24 LR:-167.3 LO:167.3);ALT=[chr5:55447995[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	151741763	-	chr2	190518529	+	.	7	59	544691_1	99.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=GGGAGGGAGGTGGGGGGCAG;MAPQ=60;MATEID=544691_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_1_151728501_151753501_316C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:62 DP:63 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:59 DR:7 LR:-184.8 LO:184.8);ALT=[chr2:190518529[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	190047656	-	chr2	190049206	+	.	8	0	1574871_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1574871_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:190047656(-)-2:190049206(-)__2_190046501_190071501D;SPAN=1550;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:120 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.103 LO:14.04);ALT=[chr2:190049206[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	25996622	-	chr5	55137495	+	.	47	57	3434600_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=G;MAPQ=8;MATEID=3434600_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_55125001_55150001_381C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:82 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:57 DR:47 LR:-257.5 LO:257.5);ALT=[chr5:55137495[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
