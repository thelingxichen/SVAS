chr3	152311738	+	chr3	152313156	+	.	102	57	2412335_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAGGTCACTGTTT;MAPQ=60;MATEID=2412335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_152292001_152317001_4C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:77 GQ:36 PL:[396.0, 36.0, 0.0] SR:57 DR:102 LR:-396.1 LO:396.1);ALT=T[chr3:152313156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
