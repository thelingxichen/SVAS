chr3	33916572	+	chr3	34533798	+	.	70	44	1938553_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTCT;MAPQ=60;MATEID=1938553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_34520501_34545501_271C;SPAN=617226;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:37 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:44 DR:70 LR:-267.4 LO:267.4);ALT=T[chr3:34533798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
