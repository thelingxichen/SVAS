chr8	32680009	+	chr8	32691262	+	.	82	43	5437009_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5437009_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_32658501_32683501_3C;SPAN=11253;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:9 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:43 DR:82 LR:-310.3 LO:310.3);ALT=G[chr8:32691262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
