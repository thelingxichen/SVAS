chr7	120290167	+	chr7	120291387	+	.	17	0	3553263_1	36.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=3553263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:120290167(+)-7:120291387(-)__7_120270501_120295501D;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:72 GQ:36.8 PL:[36.8, 0.0, 135.8] SR:0 DR:17 LR:-36.61 LO:39.93);ALT=G[chr7:120291387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
