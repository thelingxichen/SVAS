chr9	86243875	+	chr9	86258342	+	ACCGGATTCCATGGCTCTGTAACTTGCATGACATTTTACTA	0	12	4305808_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACCGGATTCCATGGCTCTGTAACTTGCATGACATTTTACTA;MAPQ=60;MATEID=4305808_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_86240001_86265001_385C;SPAN=14467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:116 GQ:8.3 PL:[8.3, 0.0, 272.3] SR:12 DR:0 LR:-8.185 LO:23.46);ALT=G[chr9:86258342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	86593215	+	chr9	86595433	+	.	14	0	4307117_1	23.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=4307117_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:86593215(+)-9:86595433(-)__9_86583001_86608001D;SPAN=2218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:0 DR:14 LR:-23.73 LO:30.57);ALT=T[chr9:86595433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	86593215	+	chr9	86595053	+	.	19	0	4307116_1	37.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4307116_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:86593215(+)-9:86595053(-)__9_86583001_86608001D;SPAN=1838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:95 GQ:37.1 PL:[37.1, 0.0, 192.2] SR:0 DR:19 LR:-36.98 LO:43.06);ALT=T[chr9:86595053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
