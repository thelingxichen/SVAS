chr3	28283303	+	chr3	28304779	+	.	7	9	1325204_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1325204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_28273001_28298001_310C;SPAN=21476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:9 DR:7 LR:-21.68 LO:25.03);ALT=G[chr3:28304779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	28382114	+	chr3	28390092	+	.	6	6	1325349_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1325349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_28371001_28396001_241C;SPAN=7978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:123 GQ:3.3 PL:[0.0, 3.3, 303.6] SR:6 DR:6 LR:3.615 LO:16.17);ALT=C[chr3:28390092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
