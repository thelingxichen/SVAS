chr12	45610174	+	chr12	45695796	+	.	0	8	5171913_1	15.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5171913_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_45692501_45717501_298C;SPAN=85622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:8 DR:0 LR:-15.84 LO:18.23);ALT=G[chr12:45695796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	45903153	+	chr12	45909940	+	.	0	63	5172241_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5172241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_45888501_45913501_137C;SPAN=6787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:36 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:63 DR:0 LR:-184.8 LO:184.8);ALT=A[chr12:45909940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	46123922	+	chr12	46124998	+	.	0	4	5172877_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5172877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_46109001_46134001_29C;SPAN=1076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:52 GQ:0.6 PL:[0.0, 0.6, 125.4] SR:4 DR:0 LR:0.8841 LO:7.279);ALT=T[chr12:46124998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	46355642	+	chr12	46384135	+	TCCATGTCTTCATACTTCTTATCTCCCATATTTAGGGTACATACAGTTTTCTTCTTCATTTCTCTTTGGAAAAGGGTTT	2	20	5173292_1	49.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TCCATGTCTTCATACTTCTTATCTCCCATATTTAGGGTACATACAGTTTTCTTCTTCATTTCTCTTTGGAAAAGGGTTT;MAPQ=60;MATEID=5173292_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_46378501_46403501_173C;SPAN=28493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:60 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:20 DR:2 LR:-49.76 LO:50.57);ALT=T[chr12:46384135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	46633678	+	chr12	46636982	+	.	0	7	5174045_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5174045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_46623501_46648501_240C;SPAN=3304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:63 GQ:6.2 PL:[6.2, 0.0, 144.8] SR:7 DR:0 LR:-6.039 LO:13.91);ALT=T[chr12:46636982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	46765164	+	chr12	46766291	+	.	0	6	5174274_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5174274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_46746001_46771001_47C;SPAN=1127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:112 GQ:10.2 PL:[0.0, 10.2, 290.4] SR:6 DR:0 LR:10.54 LO:9.947);ALT=T[chr12:46766291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
