chr8	594397	+	chr8	599415	+	CAA	0	48	3709440_1	99.0	.	EVDNC=ASSMB;INSERTION=CAA;MAPQ=60;MATEID=3709440_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_588001_613001_148C;SPAN=5018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:28 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:48 DR:0 LR:-141.9 LO:141.9);ALT=G[chr8:599415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	625151	+	chr8	626487	+	.	13	0	3709570_1	26.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3709570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:625151(+)-8:626487(-)__8_612501_637501D;SPAN=1336;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.66 LO:29.98);ALT=C[chr8:626487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	642615	+	chr8	665861	+	.	0	23	3709615_1	65.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=3709615_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_661501_686501_45C;SPAN=23246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:23 DR:0 LR:-65.7 LO:65.7);ALT=G[chr8:665861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	642655	+	chr8	681139	+	.	18	0	3709757_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3709757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:642655(+)-8:681139(-)__8_637001_662001D;SPAN=38484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:54 GQ:44.9 PL:[44.9, 0.0, 84.5] SR:0 DR:18 LR:-44.79 LO:45.51);ALT=A[chr8:681139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	666008	+	chr8	681140	+	.	16	7	3709654_1	34.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3709654_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CACA;SCTG=c_8_661501_686501_45C;SPAN=15132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:105 GQ:34.4 PL:[34.4, 0.0, 219.2] SR:7 DR:16 LR:-34.27 LO:42.13);ALT=C[chr8:681140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	963696	+	chr8	967540	+	.	94	0	3710609_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3710609_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:963696(+)-8:967540(-)__8_955501_980501D;SPAN=3844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:30 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:0 DR:94 LR:-277.3 LO:277.3);ALT=T[chr8:967540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	1285858	+	chr8	1284407	+	.	41	0	3711486_1	99.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3711486_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:1284407(-)-8:1285858(+)__8_1274001_1299001D;SPAN=1451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:112 GQ:99 PL:[105.2, 0.0, 164.6] SR:0 DR:41 LR:-105.0 LO:105.8);ALT=]chr8:1285858]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	1521670	+	chr8	1519457	+	.	24	0	3712317_1	54.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=3712317_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:1519457(-)-8:1521670(+)__8_1519001_1544001D;SPAN=2213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:90 GQ:54.8 PL:[54.8, 0.0, 163.7] SR:0 DR:24 LR:-54.84 LO:57.85);ALT=]chr8:1521670]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	1712133	+	chr8	1719095	+	.	10	0	3712719_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3712719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:1712133(+)-8:1719095(-)__8_1715001_1740001D;SPAN=6962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=G[chr8:1719095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	2556847	+	chr8	2537451	+	.	47	0	3715554_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3715554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:2537451(-)-8:2556847(+)__8_2523501_2548501D;SPAN=19396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:61 GQ:6.8 PL:[138.8, 0.0, 6.8] SR:0 DR:47 LR:-145.3 LO:145.3);ALT=]chr8:2556847]T;VARTYPE=BND:DUP-th;JOINTYPE=th
