chr3	190232009	+	chr3	190236296	+	.	6	2	1852143_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1852143_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_190218001_190243001_249C;SPAN=4287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:109 GQ:6.3 PL:[0.0, 6.3, 277.2] SR:2 DR:6 LR:6.424 LO:12.17);ALT=G[chr3:190236296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
