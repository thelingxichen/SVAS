chr6	168830425	+	chr6	168829313	+	.	31	0	3119777_1	86.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3119777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:168829313(-)-6:168830425(+)__6_168829501_168854501D;SPAN=1112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:60 GQ:59.6 PL:[86.0, 0.0, 59.6] SR:0 DR:31 LR:-86.33 LO:86.33);ALT=]chr6:168830425]G;VARTYPE=BND:DUP-th;JOINTYPE=th
