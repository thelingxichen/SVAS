chr1	14438565	+	chr1	14436309	+	.	14	99	74271_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GATT;MAPQ=60;MATEID=74271_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_14430501_14455501_82C;SPAN=2256;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:44 GQ:27 PL:[297.0, 27.0, 0.0] SR:99 DR:14 LR:-297.1 LO:297.1);ALT=]chr1:14438565]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	14438565	+	chr1	14436656	+	TCAGCGTCAAGTAGGAGCTGTACTAAAAATTTATGTAA	85	145	74277_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GTTT;INSERTION=TCAGCGTCAAGTAGGAGCTGTACTAAAAATTTATGTAA;MAPQ=60;MATEID=74277_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_1_14430501_14455501_82C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:199 DP:44 GQ:53.8 PL:[590.8, 53.8, 0.0] SR:145 DR:85 LR:-590.8 LO:590.8);ALT=]chr1:14438565]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	14437074	+	chr1	14438940	+	.	0	86	74282_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=74282_2;MATENM=2;NM=3;NUMPARTS=2;SCTG=c_1_14430501_14455501_323C;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:32 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:86 DR:0 LR:-254.2 LO:254.2);ALT=T[chr1:14438940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
