chr2	60654032	+	chr2	60655437	+	.	0	46	1030870_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GGTC;MAPQ=60;MATEID=1030870_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_60637501_60662501_302C;SPAN=1405;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:46 DP:98 GQ:99 PL:[125.3, 0.0, 112.1] SR:46 DR:0 LR:-125.3 LO:125.3);ALT=C[chr2:60655437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
