chr2	159132848	-	chr2	159134028	+	.	6	2	1452473_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=47;MATEID=1452473_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_159127501_159152501_457C;SPAN=1180;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:163 GQ:17.5 PL:[0.0, 17.5, 429.1] SR:2 DR:6 LR:17.75 LO:12.95);ALT=[chr2:159134028[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	160095988	+	chr2	160100167	+	.	69	95	1456739_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAA;MAPQ=60;MATEID=1456739_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_160083001_160108001_378C;SPAN=4179;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:112 GQ:36 PL:[396.0, 36.0, 0.0] SR:95 DR:69 LR:-396.1 LO:396.1);ALT=A[chr2:160100167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	160149126	+	chr2	160151649	+	.	82	78	1456963_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAGAATTTC;MAPQ=60;MATEID=1456963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_160132001_160157001_263C;SPAN=2523;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:126 DP:72 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:78 DR:82 LR:-373.0 LO:373.0);ALT=C[chr2:160151649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
