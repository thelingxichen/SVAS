chr7	95906652	+	chr7	95926210	+	.	2	3	3465657_1	4.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3465657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_95893001_95918001_177C;SPAN=19558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:45 GQ:4.4 PL:[4.4, 0.0, 103.4] SR:3 DR:2 LR:-4.313 LO:9.938);ALT=T[chr7:95926210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	95906687	+	chr7	95951310	+	.	8	0	3465806_1	15.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=3465806_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:95906687(+)-7:95951310(-)__7_95942001_95967001D;SPAN=44623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:0 DR:8 LR:-15.84 LO:18.23);ALT=T[chr7:95951310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	96318328	+	chr7	96339057	+	.	73	0	3467134_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=3467134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:96318328(+)-7:96339057(-)__7_96334001_96359001D;SPAN=20729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:0 DR:73 LR:-237.7 LO:237.7);ALT=T[chr7:96339057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	96324205	+	chr7	96339000	+	.	92	115	3467135_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=18;MATEID=3467135_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_96334001_96359001_86C;SPAN=14795;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:173 DP:66 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:115 DR:92 LR:-511.6 LO:511.6);ALT=T[chr7:96339000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	96475901	+	chr7	96481995	+	.	134	44	3467757_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCAACTGGAACTTTC;MAPQ=60;MATEID=3467757_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_96456501_96481501_331C;SPAN=6094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:24 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:44 DR:134 LR:-435.7 LO:435.7);ALT=C[chr7:96481995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	96747210	+	chr7	96810322	+	.	0	24	3468646_1	64.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3468646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_96799501_96824501_369C;SPAN=63112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:54 GQ:64.7 PL:[64.7, 0.0, 64.7] SR:24 DR:0 LR:-64.59 LO:64.6);ALT=G[chr7:96810322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	97420483	+	chr7	97402640	+	.	33	44	3470877_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCCT;MAPQ=60;MATEID=3470877_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_97387501_97412501_13C;SPAN=17843;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:33 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:44 DR:33 LR:-184.8 LO:184.8);ALT=]chr7:97420483]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	97599159	+	chr7	97601445	+	.	5	9	3471127_1	5.0	.	DISC_MAPQ=22;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=48;MATEID=3471127_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_97583501_97608501_443C;SPAN=2286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:116 GQ:5 PL:[5.0, 0.0, 275.6] SR:9 DR:5 LR:-4.884 LO:21.06);ALT=T[chr7:97601445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	97688063	+	chr7	97689132	-	.	8	0	3471790_1	3.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3471790_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:97688063(+)-7:97689132(+)__7_97681501_97706501D;SPAN=1069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=T]chr7:97689132];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	97911766	+	chr7	97920417	+	.	4	4	3473098_1	0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CTGCAGG;MAPQ=60;MATEID=3473098_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_97902001_97927001_107C;SPAN=8651;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:4 DR:4 LR:0.9554 LO:14.66);ALT=G[chr7:97920417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
