chr13	39057319	+	chr13	39060202	+	.	58	42	8013961_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGAA;MAPQ=60;MATEID=8013961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_39053001_39078001_357C;SPAN=2883;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:77 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:42 DR:58 LR:-234.4 LO:234.4);ALT=A[chr13:39060202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	39934199	+	chr13	39935481	+	.	76	54	8017564_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AGTCTCACTCTGTCGCC;MAPQ=60;MATEID=8017564_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_39910501_39935501_155C;SPAN=1282;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:100 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:54 DR:76 LR:-340.0 LO:340.0);ALT=C[chr13:39935481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
