chr13	90862855	+	chr13	90864807	+	.	68	59	8213289_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAT;MAPQ=60;MATEID=8213289_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_90846001_90871001_366C;SPAN=1952;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:89 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:59 DR:68 LR:-303.7 LO:303.7);ALT=T[chr13:90864807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
