chr1	233095350	+	chr18	31269079	-	.	52	39	9972450_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GCCT;MAPQ=60;MATEID=9972450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_31262001_31287001_317C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:78 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:39 DR:52 LR:-237.7 LO:237.7);ALT=C]chr18:31269079];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	233295888	-	chr18	31182338	+	.	73	65	9972118_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=9972118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_31164001_31189001_16C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:76 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:65 DR:73 LR:-346.6 LO:346.6);ALT=[chr18:31182338[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr18	31699744	+	chr18	31701578	+	.	71	44	9974133_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=9974133_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_31678501_31703501_285C;SPAN=1834;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:77 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:44 DR:71 LR:-287.2 LO:287.2);ALT=C[chr18:31701578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
