chr18	32621625	+	chr18	32650157	+	.	0	12	6585562_1	29.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6585562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_32634001_32659001_277C;SPAN=28532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:12 DR:0 LR:-29.05 LO:29.82);ALT=G[chr18:32650157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	32870388	+	chr18	32885936	+	.	11	0	6586095_1	25.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6586095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:32870388(+)-18:32885936(-)__18_32879001_32904001D;SPAN=15548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:41 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:0 DR:11 LR:-25.2 LO:26.55);ALT=G[chr18:32885936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	32920728	+	chr18	32924329	+	.	16	0	6586267_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6586267_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:32920728(+)-18:32924329(-)__18_32903501_32928501D;SPAN=3601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:85 GQ:29.9 PL:[29.9, 0.0, 175.1] SR:0 DR:16 LR:-29.79 LO:35.79);ALT=T[chr18:32924329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	33552762	+	chr18	33554857	+	.	8	0	6587828_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6587828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:33552762(+)-18:33554857(-)__18_33540501_33565501D;SPAN=2095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=A[chr18:33554857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	33557563	+	chr18	33558791	+	.	0	6	6587840_1	0	.	EVDNC=ASSMB;HOMSEQ=TTTTCAG;MAPQ=60;MATEID=6587840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_33540501_33565501_251C;SPAN=1228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:70 GQ:0.8 PL:[0.8, 0.0, 169.1] SR:6 DR:0 LR:-0.8413 LO:11.21);ALT=G[chr18:33558791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	33710034	+	chr18	33713200	+	.	0	8	6588034_1	15.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6588034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_33712001_33737001_227C;SPAN=3166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:8 DR:0 LR:-15.03 LO:17.94);ALT=G[chr18:33713200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	33713279	+	chr18	33716270	+	.	0	8	6588037_1	7.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6588037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_33712001_33737001_297C;SPAN=2991;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:8 DR:0 LR:-7.172 LO:15.95);ALT=T[chr18:33716270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34377015	+	chr18	34378412	+	.	3	2	6589612_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6589612_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_34373501_34398501_65C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:89 GQ:10.8 PL:[0.0, 10.8, 237.6] SR:2 DR:3 LR:10.91 LO:6.32);ALT=T[chr18:34378412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34385466	+	chr18	34387810	+	.	2	16	6589638_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6589638_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_34373501_34398501_257C;SPAN=2344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:96 GQ:33.5 PL:[33.5, 0.0, 198.5] SR:16 DR:2 LR:-33.41 LO:40.23);ALT=C[chr18:34387810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34385517	+	chr18	34408690	+	.	10	0	6589716_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6589716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:34385517(+)-18:34408690(-)__18_34398001_34423001D;SPAN=23173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:44 GQ:21.2 PL:[21.2, 0.0, 83.9] SR:0 DR:10 LR:-21.09 LO:23.3);ALT=A[chr18:34408690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34387897	+	chr18	34398857	+	.	0	19	6589717_1	52.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6589717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_34398001_34423001_83C;SPAN=10960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:37 GQ:36.2 PL:[52.7, 0.0, 36.2] SR:19 DR:0 LR:-52.84 LO:52.84);ALT=T[chr18:34398857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34387942	+	chr18	34408683	+	.	12	0	6589719_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6589719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:34387942(+)-18:34408683(-)__18_34398001_34423001D;SPAN=20741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:42 GQ:28.4 PL:[28.4, 0.0, 71.3] SR:0 DR:12 LR:-28.23 LO:29.36);ALT=A[chr18:34408683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	34398938	+	chr18	34408646	+	.	19	19	6589724_1	75.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6589724_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_34398001_34423001_111C;SPAN=9708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:75 GQ:75.5 PL:[75.5, 0.0, 105.2] SR:19 DR:19 LR:-75.41 LO:75.7);ALT=T[chr18:34408646[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
