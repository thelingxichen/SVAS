chr8	26240748	+	chr8	26248759	+	.	0	43	3790268_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=3790268_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_26239501_26264501_45C;SPAN=8011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:102 GQ:99 PL:[114.5, 0.0, 131.0] SR:43 DR:0 LR:-114.3 LO:114.4);ALT=T[chr8:26248759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	26241231	+	chr8	26248752	+	.	51	0	3790270_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3790270_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:26241231(+)-8:26248752(-)__8_26239501_26264501D;SPAN=7521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:131 GQ:99 PL:[133.1, 0.0, 182.6] SR:0 DR:51 LR:-132.9 LO:133.3);ALT=G[chr8:26248752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	26248942	+	chr8	26252744	+	.	3	8	3790295_1	8.0	.	DISC_MAPQ=40;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3790295_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_8_26239501_26264501_1C;SPAN=3802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:91 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:8 DR:3 LR:-8.356 LO:19.82);ALT=G[chr8:26252744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	26248942	+	chr8	26265513	+	CCCTTCGCCACAAGAAGATGGGCAGATCATGTTTGATGTGGAAATGCACACCAGCAGGGACCATAGCTCT	3	13	3790296_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=CCCTTCGCCACAAGAAGATGGGCAGATCATGTTTGATGTGGAAATGCACACCAGCAGGGACCATAGCTCT;MAPQ=60;MATEID=3790296_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_26239501_26264501_1C;SPAN=16571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:13 DR:3 LR:-35.16 LO:36.62);ALT=G[chr8:26265513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	26265892	+	chr8	26267879	+	.	2	3	3789932_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3789932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_26264001_26289001_34C;SPAN=1987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:92 GQ:11.4 PL:[0.0, 11.4, 244.2] SR:3 DR:2 LR:11.72 LO:6.262);ALT=G[chr8:26267879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
