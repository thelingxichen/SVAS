chr14	42675285	+	chr14	42614492	+	.	42	50	8465748_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=TG;MAPQ=60;MATEID=8465748_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_42654501_42679501_87C;SPAN=60793;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:74 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:50 DR:42 LR:-224.5 LO:224.5);ALT=]chr14:42675285]T;VARTYPE=BND:DUP-th;JOINTYPE=th
