chr9	120759409	-	chr9	120760659	+	.	2	3	4418978_1	0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=AGAGGAAAA;MAPQ=60;MATEID=4418978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_120736001_120761001_14C;SPAN=1250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:3 DR:2 LR:6.844 LO:6.647);ALT=[chr9:120760659[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
