chr4	90756846	+	chr4	90758113	+	.	17	22	2084387_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2084387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_90748001_90773001_20C;SPAN=1267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:103 GQ:71.3 PL:[71.3, 0.0, 176.9] SR:22 DR:17 LR:-71.13 LO:73.69);ALT=G[chr4:90758113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	91596798	+	chr4	91602909	+	.	43	35	2086903_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTGTTTTTATCTT;MAPQ=60;MATEID=2086903_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_91581001_91606001_199C;SPAN=6111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:63 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:35 DR:43 LR:-184.8 LO:184.8);ALT=T[chr4:91602909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	91760140	+	chrX	12994394	-	.	21	0	2087126_1	0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=2087126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:91760140(+)-23:12994394(+)__4_91752501_91777501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:21 DP:332 GQ:20.3 PL:[0.0, 20.3, 845.0] SR:0 DR:21 LR:20.63 LO:36.37);ALT=T]chrX:12994394];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chrX	11953199	+	chrX	11959436	+	.	67	49	7365640_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGGTGATTTTTTTT;MAPQ=60;MATEID=7365640_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_23_11931501_11956501_193C;SPAN=6237;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:42 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:49 DR:67 LR:-283.9 LO:283.9);ALT=T[chrX:11959436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	12809738	+	chrX	12817324	+	.	17	20	7366608_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7366608_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_12813501_12838501_5C;SPAN=7586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:20 DR:17 LR:-89.12 LO:89.12);ALT=G[chrX:12817324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	12993328	+	chrX	12995028	+	.	42	0	7366954_1	65.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=7366954_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:12993328(+)-23:12995028(-)__23_12985001_13010001D;SPAN=1700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:270 GQ:65.5 PL:[65.5, 0.0, 590.3] SR:0 DR:42 LR:-65.49 LO:90.09);ALT=G[chrX:12995028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	13707348	+	chrX	13721875	+	.	13	0	7368068_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7368068_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:13707348(+)-23:13721875(-)__23_13720001_13745001D;SPAN=14527;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:30 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:0 DR:13 LR:-34.79 LO:34.79);ALT=C[chrX:13721875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	13707408	+	chrX	13726838	+	.	13	3	7368071_1	43.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7368071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_13720001_13745001_124C;SPAN=19430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:36 GQ:43.1 PL:[43.1, 0.0, 43.1] SR:3 DR:13 LR:-43.06 LO:43.06);ALT=G[chrX:13726838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	13762638	+	chrX	13764437	+	.	0	7	7368010_1	9.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7368010_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_13744501_13769501_109C;SPAN=1799;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=G[chrX:13764437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
