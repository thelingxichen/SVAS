chr8	77337385	+	chr8	77338427	+	.	59	42	5511401_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTT;MAPQ=60;MATEID=5511401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_77322001_77347001_30C;SPAN=1042;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:34 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:42 DR:59 LR:-254.2 LO:254.2);ALT=T[chr8:77338427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
