chr1	51436172	+	chr1	51439562	+	.	34	39	149046_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGTT;MAPQ=60;MATEID=149046_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_51425501_51450501_131C;SPAN=3390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:95 GQ:63.5 PL:[165.8, 0.0, 63.5] SR:39 DR:34 LR:-168.1 LO:168.1);ALT=T[chr1:51439562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	51937463	+	chr1	51984869	+	.	12	0	150639_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=150639_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:51937463(+)-1:51984869(-)__1_51964501_51989501D;SPAN=47406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=A[chr1:51984869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52082859	+	chr1	52135105	+	.	11	0	151204_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=151204_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:52082859(+)-1:52135105(-)__1_52062501_52087501D;SPAN=52246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:0 DR:11 LR:-26.02 LO:26.98);ALT=T[chr1:52135105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52082893	+	chr1	52117662	+	.	2	2	151205_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=151205_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_52062501_52087501_227C;SPAN=34769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:40 GQ:2.3 PL:[2.3, 0.0, 94.7] SR:2 DR:2 LR:-2.367 LO:7.756);ALT=G[chr1:52117662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52306187	+	chr1	52343947	+	.	7	12	151765_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=151765_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_52332001_52357001_207C;SPAN=37760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:47 GQ:36.8 PL:[36.8, 0.0, 76.4] SR:12 DR:7 LR:-36.78 LO:37.57);ALT=C[chr1:52343947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52493022	+	chr1	52520670	+	TTGCAAGCTCCACACCAGGATTTATGAATAATCACCATCAGGGGCAGTCCACTGGCAGCTGCTTCTTTCTTCCCATCTTCCAGTGTCCTCCAATGAATATGATCTCCAAA	0	41	152267_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TTGCAAGCTCCACACCAGGATTTATGAATAATCACCATCAGGGGCAGTCCACTGGCAGCTGCTTCTTTCTTCCCATCTTCCAGTGTCCTCCAATGAATATGATCTCCAAA;MAPQ=60;MATEID=152267_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_52503501_52528501_345C;SPAN=27648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:41 DR:0 LR:-128.7 LO:128.7);ALT=T[chr1:52520670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52494353	+	chr1	52520780	+	.	14	0	152270_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=152270_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:52494353(+)-1:52520780(-)__1_52503501_52528501D;SPAN=26427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:49 GQ:32.9 PL:[32.9, 0.0, 85.7] SR:0 DR:14 LR:-32.94 LO:34.25);ALT=T[chr1:52520780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52507318	+	chr1	52520776	+	.	20	0	152289_1	43.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=152289_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:52507318(+)-1:52520776(-)__1_52503501_52528501D;SPAN=13458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:85 GQ:43.1 PL:[43.1, 0.0, 161.9] SR:0 DR:20 LR:-42.99 LO:46.94);ALT=A[chr1:52520776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	52992047	+	chr1	53018603	+	.	3	5	153715_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=153715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_52969001_52994001_114C;SPAN=26556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:27 GQ:15.8 PL:[15.8, 0.0, 48.8] SR:5 DR:3 LR:-15.79 LO:16.77);ALT=T[chr1:53018603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53068155	+	chr1	53072354	+	.	11	0	153847_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=153847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53068155(+)-1:53072354(-)__1_53067001_53092001D;SPAN=4199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:81 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:0 DR:11 LR:-14.37 LO:22.89);ALT=T[chr1:53072354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53393053	+	chr1	53407465	+	.	11	0	154932_1	12.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=154932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53393053(+)-1:53407465(-)__1_53385501_53410501D;SPAN=14412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:0 DR:11 LR:-12.74 LO:22.52);ALT=C[chr1:53407465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53393137	+	chr1	53413679	+	TTTGTGAAGCCTGGAGCTGAGAATTCAAGAGACTACCCTGACTTGGCAGAAGAAGC	0	20	154934_1	55.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TTTGTGAAGCCTGGAGCTGAGAATTCAAGAGACTACCCTGACTTGGCAGAAGAAGC;MAPQ=60;MATEID=154934_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_53385501_53410501_163C;SPAN=20542;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:40 GQ:41.9 PL:[55.1, 0.0, 41.9] SR:20 DR:0 LR:-55.28 LO:55.28);ALT=G[chr1:53413679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53480715	+	chr1	53493637	+	.	41	15	155368_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAG;MAPQ=60;MATEID=155368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53459001_53484001_286C;SPAN=12922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:43 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:15 DR:41 LR:-141.9 LO:141.9);ALT=G[chr1:53493637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53480761	+	chr1	53504586	+	.	74	0	155369_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=155369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53480761(+)-1:53504586(-)__1_53459001_53484001D;SPAN=23825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:31 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:0 DR:74 LR:-217.9 LO:217.9);ALT=T[chr1:53504586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53493744	+	chr1	53504587	+	.	3	65	155259_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=155259_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53483501_53508501_176C;SPAN=10843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:92 GQ:21.5 PL:[199.7, 0.0, 21.5] SR:65 DR:3 LR:-207.6 LO:207.6);ALT=G[chr1:53504587[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53504718	+	chr1	53513528	+	.	0	26	155173_1	69.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=155173_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53508001_53533001_332C;SPAN=8810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:59 GQ:69.8 PL:[69.8, 0.0, 73.1] SR:26 DR:0 LR:-69.84 LO:69.85);ALT=G[chr1:53513528[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53594099	+	chr1	53595604	+	AATAACCTCGTGAAGGAGGTATTCTTCCCACTTTATAGATAAGGACACTGAGGCTCAGATGCTAAAAGGCTTGTTTACATTTGCACATCTAGAGGGTGACTCCAAAGCCCTGTTCCTGCCCTGTAGCCTTTGCAGATTTCAACCACCCCCGCCCATGCTTCCTGCTCCCCCGCCA	22	95	155483_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CAT;INSERTION=AATAACCTCGTGAAGGAGGTATTCTTCCCACTTTATAGATAAGGACACTGAGGCTCAGATGCTAAAAGGCTTGTTTACATTTGCACATCTAGAGGGTGACTCCAAAGCCCTGTTCCTGCCCTGTAGCCTTTGCAGATTTCAACCACCCCCGCCCATGCTTCCTGCTCCCCCGCCA;MAPQ=60;MATEID=155483_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_1_53581501_53606501_217C;SPAN=1505;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:54 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:95 DR:22 LR:-320.2 LO:320.2);ALT=T[chr1:53595604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53682531	+	chr1	53685933	+	ATTGTAAGGCTTGATGGTGCTGCTTAAAATCTCGATGGAATTTTCTCTTGCACACAGCTTGCACTTCTGGACCATGGAAGCACTGCCACGGCCCCCCTTCAGTGCCACACTGTCCATCAGCCGGATGTACTGCCACTTGTCCGAAATCTCACCACAGTTGCCACATTTCAT	0	37	155827_1	96.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTT;INSERTION=ATTGTAAGGCTTGATGGTGCTGCTTAAAATCTCGATGGAATTTTCTCTTGCACACAGCTTGCACTTCTGGACCATGGAAGCACTGCCACGGCCCCCCTTCAGTGCCACACTGTCCATCAGCCGGATGTACTGCCACTTGTCCGAAATCTCACCACAGTTGCCACATTTCAT;MAPQ=60;MATEID=155827_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_53679501_53704501_28C;SPAN=3402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:96 GQ:96.2 PL:[96.2, 0.0, 135.8] SR:37 DR:0 LR:-96.13 LO:96.52);ALT=C[chr1:53685933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53682590	+	chr1	53686241	+	.	8	0	155828_1	1.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=155828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53682590(+)-1:53686241(-)__1_53679501_53704501D;SPAN=3651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=G[chr1:53686241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53684214	+	chr1	53686241	+	.	27	0	155832_1	65.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=155832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53684214(+)-1:53686241(-)__1_53679501_53704501D;SPAN=2027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:88 GQ:65.3 PL:[65.3, 0.0, 147.8] SR:0 DR:27 LR:-65.29 LO:67.06);ALT=A[chr1:53686241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53684643	+	chr1	53686240	+	.	23	0	155835_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=155835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53684643(+)-1:53686240(-)__1_53679501_53704501D;SPAN=1597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:90 GQ:51.5 PL:[51.5, 0.0, 167.0] SR:0 DR:23 LR:-51.54 LO:54.94);ALT=A[chr1:53686240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53692816	+	chr1	53694543	+	.	2	22	155859_1	60.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=155859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53679501_53704501_26C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:70 GQ:60.2 PL:[60.2, 0.0, 109.7] SR:22 DR:2 LR:-60.26 LO:61.05);ALT=C[chr1:53694543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53694628	+	chr1	53701248	+	.	0	15	155864_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=155864_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53679501_53704501_20C;SPAN=6620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:78 GQ:28.4 PL:[28.4, 0.0, 160.4] SR:15 DR:0 LR:-28.38 LO:33.71);ALT=T[chr1:53701248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53694667	+	chr1	53704105	+	.	9	0	155865_1	10.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=155865_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53694667(+)-1:53704105(-)__1_53679501_53704501D;SPAN=9438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:0 DR:9 LR:-10.2 LO:18.38);ALT=T[chr1:53704105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53699357	+	chr1	53704091	+	.	13	0	155876_1	24.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=155876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53699357(+)-1:53704091(-)__1_53679501_53704501D;SPAN=4734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:69 GQ:24.2 PL:[24.2, 0.0, 143.0] SR:0 DR:13 LR:-24.22 LO:29.08);ALT=G[chr1:53704091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53701347	+	chr1	53704105	+	.	8	0	155889_1	5.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=155889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53701347(+)-1:53704105(-)__1_53679501_53704501D;SPAN=2758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:0 DR:8 LR:-5.276 LO:15.61);ALT=A[chr1:53704105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54395819	+	chr1	54405657	+	.	0	21	157452_1	50.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=157452_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=CC;SCTG=c_1_54390001_54415001_171C;SPAN=9838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:72 GQ:50 PL:[50.0, 0.0, 122.6] SR:21 DR:0 LR:-49.81 LO:51.6);ALT=C[chr1:54405657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54395867	+	chr1	54411223	+	.	36	0	157455_1	96.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=157455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:54395867(+)-1:54411223(-)__1_54390001_54415001D;SPAN=15356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:84 GQ:96.2 PL:[96.2, 0.0, 106.1] SR:0 DR:36 LR:-96.08 LO:96.12);ALT=T[chr1:54411223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54405793	+	chr1	54411225	+	.	13	0	157499_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=157499_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:54405793(+)-1:54411225(-)__1_54390001_54415001D;SPAN=5432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=A[chr1:54411225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54497980	+	chr1	54502283	+	.	8	29	157766_1	97.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=157766_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54488001_54513001_130C;SPAN=4303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:78 GQ:91.1 PL:[97.7, 0.0, 91.1] SR:29 DR:8 LR:-97.71 LO:97.71);ALT=T[chr1:54502283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54502391	+	chr1	54506429	+	.	4	7	157781_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=157781_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54488001_54513001_8C;SPAN=4038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:7 DR:4 LR:-18.43 LO:23.96);ALT=A[chr1:54506429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54506548	+	chr1	54509045	+	.	8	0	157792_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=157792_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:54506548(+)-1:54509045(-)__1_54488001_54513001D;SPAN=2497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:0 DR:8 LR:-6.089 LO:15.75);ALT=A[chr1:54509045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54507480	+	chr1	54509046	+	.	2	9	157794_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=157794_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_54488001_54513001_307C;SPAN=1566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:84 GQ:10.4 PL:[10.4, 0.0, 191.9] SR:9 DR:2 LR:-10.25 LO:20.2);ALT=T[chr1:54509046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54507480	+	chr1	54512940	+	GGAATATAACTATTTTTCCGTCATCGGCTTGAAGATAAAAAGTCCATGAAGAGGTTATGAAGCTCTGTGCGGAGTCCATCATGTCACTCCAGAATGACCTCACCAGAGTTAGAGGAAAGAGTAGGTGCATTTTTGGCATCAGGGACATAAGTTGTTCTTGTCTCAGTTCAGCGAATGGCAGCTGATTCTGGCAACCAAGATGGCAAGCATATTGCTCATCAGATTGGGAATATGCTTCTGTACATG	0	41	157795_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGAATATAACTATTTTTCCGTCATCGGCTTGAAGATAAAAAGTCCATGAAGAGGTTATGAAGCTCTGTGCGGAGTCCATCATGTCACTCCAGAATGACCTCACCAGAGTTAGAGGAAAGAGTAGGTGCATTTTTGGCATCAGGGACATAAGTTGTTCTTGTCTCAGTTCAGCGAATGGCAGCTGATTCTGGCAACCAAGATGGCAAGCATATTGCTCATCAGATTGGGAATATGCTTCTGTACATG;MAPQ=60;MATEID=157795_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_54488001_54513001_307C;SPAN=5460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:87 GQ:98.6 PL:[111.8, 0.0, 98.6] SR:41 DR:0 LR:-111.8 LO:111.8);ALT=T[chr1:54512940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54509198	+	chr1	54511365	+	.	4	15	157800_1	32.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=157800_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_54488001_54513001_307C;SPAN=2167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:76 GQ:32.3 PL:[32.3, 0.0, 151.1] SR:15 DR:4 LR:-32.23 LO:36.67);ALT=G[chr1:54511365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54511460	+	chr1	54512940	+	.	0	32	157817_1	94.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=157817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54512501_54537501_236C;SPAN=1480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:42 GQ:5.3 PL:[94.4, 0.0, 5.3] SR:32 DR:0 LR:-98.59 LO:98.59);ALT=C[chr1:54512940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54511461	+	chr1	54518673	+	.	13	2	157818_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=157818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54512501_54537501_293C;SPAN=7212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:2 DR:13 LR:-23.73 LO:30.57);ALT=T[chr1:54518673[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54513047	+	chr1	54518672	+	.	0	94	157820_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=157820_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54512501_54537501_242C;SPAN=5625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:131 GQ:40.7 PL:[275.0, 0.0, 40.7] SR:94 DR:0 LR:-284.5 LO:284.5);ALT=T[chr1:54518672[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54671119	+	chr1	54675682	+	.	8	0	158249_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=158249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:54671119(+)-1:54675682(-)__1_54659501_54684501D;SPAN=4563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=T[chr1:54675682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54675805	+	chr1	54681813	+	ATTCCAGGAAGGCTATCCTTACCCCTATCCCCATACCCTGTACTTACTGGACAAAGCCAATTTACGACCACACCGCCTTCAACCAGATCAGCTGCGGGCCAAGATGATCCTGTTTGCTTTTGGCAGTGCCCTGGCTCAGGCCCGGCTCCTCTATGG	4	15	158264_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATTCCAGGAAGGCTATCCTTACCCCTATCCCCATACCCTGTACTTACTGGACAAAGCCAATTTACGACCACACCGCCTTCAACCAGATCAGCTGCGGGCCAAGATGATCCTGTTTGCTTTTGGCAGTGCCCTGGCTCAGGCCCGGCTCCTCTATGG;MAPQ=60;MATEID=158264_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_54659501_54684501_207C;SPAN=6008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:74 GQ:36.2 PL:[36.2, 0.0, 141.8] SR:15 DR:4 LR:-36.07 LO:39.69);ALT=G[chr1:54681813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54675805	+	chr1	54678171	+	.	7	8	158263_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=158263_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_54659501_54684501_207C;SPAN=2366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:8 DR:7 LR:-17.4 LO:25.39);ALT=G[chr1:54678171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54678331	+	chr1	54681813	+	.	9	6	158267_1	12.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=158267_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ATGATG;SCTG=c_1_54659501_54684501_207C;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:71 GQ:12.3 PL:[12.3, 0.0, 113.7] SR:6 DR:9 LR:-11.99 LO:17.86);ALT=G[chr1:54681813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	54682018	+	chr1	54683844	+	.	2	32	158276_1	83.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=158276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_54659501_54684501_257C;SPAN=1826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:93 GQ:83.9 PL:[83.9, 0.0, 140.0] SR:32 DR:2 LR:-83.74 LO:84.56);ALT=G[chr1:54683844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	55092274	+	chr1	55095967	+	.	81	64	159466_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=159466_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_55076001_55101001_241C;SPAN=3693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:51 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:64 DR:81 LR:-369.7 LO:369.7);ALT=G[chr1:55095967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
