chr2	4781310	+	chr2	4787357	+	.	59	32	902288_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAGATACTGCA;MAPQ=60;MATEID=902288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_4777501_4802501_200C;SPAN=6047;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:37 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:32 DR:59 LR:-214.6 LO:214.6);ALT=A[chr2:4787357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
