chr1	119401260	+	chr1	79099827	+	.	35	0	472451_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=472451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:79099827(-)-1:119401260(+)__1_119388501_119413501D;SPAN=40301433;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:0 DR:35 LR:-112.2 LO:112.2);ALT=]chr1:119401260]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	133815672	+	chr1	79276449	+	.	17	0	2928012_1	46.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=2928012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:79276449(-)-4:133815672(+)__4_133794501_133819501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:37 GQ:42.8 PL:[46.1, 0.0, 42.8] SR:0 DR:17 LR:-46.1 LO:46.1);ALT=]chr4:133815672]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	79276565	+	chr4	133815788	+	.	12	0	2928013_1	26.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=2928013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:79276565(+)-4:133815788(-)__4_133794501_133819501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:50 GQ:26 PL:[26.0, 0.0, 95.3] SR:0 DR:12 LR:-26.07 LO:28.28);ALT=C[chr4:133815788[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	80221782	+	chr1	80223029	+	.	35	38	373164_1	99.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=373164_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_1_80213001_80238001_47C;SPAN=1247;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:59 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:38 DR:35 LR:-174.9 LO:174.9);ALT=T[chr1:80223029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	133180765	+	chr4	133182990	+	.	29	0	2925584_1	71.0	.	DISC_MAPQ=7;EVDNC=DSCRD;IMPRECISE;MAPQ=7;MATEID=2925584_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:133180765(+)-4:133182990(-)__4_133182001_133207001D;SPAN=2225;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:89 GQ:71.6 PL:[71.6, 0.0, 144.2] SR:0 DR:29 LR:-71.62 LO:72.96);ALT=A[chr4:133182990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
