chr1	186342596	+	chr1	186344010	+	.	0	13	448542_1	18.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=448542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_186322501_186347501_387C;SPAN=1414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:92 GQ:18.2 PL:[18.2, 0.0, 203.0] SR:13 DR:0 LR:-17.99 LO:27.3);ALT=C[chr1:186344010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	186798169	+	chr1	186823416	+	.	6	3	449815_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=449815_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_186812501_186837501_2C;SPAN=25247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:45 GQ:11 PL:[11.0, 0.0, 96.8] SR:3 DR:6 LR:-10.92 LO:15.02);ALT=T[chr1:186823416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	187716106	+	chr1	187722533	+	.	79	53	452440_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=452440_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_187719001_187744001_260C;SPAN=6427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:107 DP:13 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:53 DR:79 LR:-316.9 LO:316.9);ALT=A[chr1:187722533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
