chr5	32167776	+	chr5	32106203	+	.	55	21	3341824_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=58;MATEID=3341824_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32144001_32169001_481C;SPAN=61573;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:60 DP:114 GQ:99 PL:[167.3, 0.0, 107.9] SR:21 DR:55 LR:-167.8 LO:167.8);ALT=]chr5:32167776]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	32350037	-	chr5	32351190	+	.	2	2	3343893_1	0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=CCTGGCTAATTTTTGTATTTTTAGTAGAGA;MAPQ=40;MATEID=3343893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32340001_32365001_169C;SPAN=1153;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:189 GQ:37.9 PL:[0.0, 37.9, 534.7] SR:2 DR:2 LR:38.0 LO:5.008);ALT=[chr5:32351190[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
