chr9	82028164	+	chr9	82033447	+	.	72	40	5902968_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTAAA;MAPQ=60;MATEID=5902968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_82026001_82051001_56C;SPAN=5283;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:17 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:40 DR:72 LR:-280.6 LO:280.6);ALT=A[chr9:82033447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
