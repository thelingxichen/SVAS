chr1	193018981	+	chr1	193028313	+	TTTAATTTTTCAAAATTCTCAGGCTCTAAACTCCATATTTCTTCTACTTGGGCTCCTCGGCA	0	12	467439_1	12.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TTTAATTTTTCAAAATTCTCAGGCTCTAAACTCCATATTTCTTCTACTTGGGCTCCTCGGCA;MAPQ=60;MATEID=467439_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_193011001_193036001_153C;SPAN=9332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:100 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:12 DR:0 LR:-12.52 LO:24.28);ALT=C[chr1:193028313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	193028848	+	chr1	193038161	+	.	9	0	467729_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=467729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:193028848(+)-1:193038161(-)__1_193035501_193060501D;SPAN=9313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:59 GQ:13.7 PL:[13.7, 0.0, 129.2] SR:0 DR:9 LR:-13.72 LO:19.22);ALT=G[chr1:193038161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	193046180	+	chr1	193050492	+	.	3	4	467760_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=467760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_193035501_193060501_143C;SPAN=4312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:84 GQ:2.7 PL:[0.0, 2.7, 207.9] SR:4 DR:3 LR:2.952 LO:10.72);ALT=G[chr1:193050492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	193091462	+	chr1	193094241	+	.	6	3	467660_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=467660_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_193084501_193109501_274C;SPAN=2779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:124 GQ:10.2 PL:[0.0, 10.2, 320.1] SR:3 DR:6 LR:10.49 LO:11.77);ALT=G[chr1:193094241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
