chr2	46447911	-	chr6	109858802	+	.	23	0	4353918_1	66.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4353918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:46447911(-)-6:109858802(-)__6_109858001_109883001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:23 DP:11 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:23 LR:-66.02 LO:66.02);ALT=[chr6:109858802[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	26031699	+	chr5	26003834	+	.	65	32	3304573_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=3304573_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_26019001_26044001_266C;SPAN=27865;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:86 DP:121 GQ:40.1 PL:[251.3, 0.0, 40.1] SR:32 DR:65 LR:-259.5 LO:259.5);ALT=]chr5:26031699]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	26457048	+	chrX	101413096	+	.	8	20	3307024_1	72.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCTTCTTCTTCTTCTTCTTCTTCTTCTTCTT;MAPQ=60;MATEID=3307024_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_26435501_26460501_413C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:25 DP:18 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:20 DR:8 LR:-72.62 LO:72.62);ALT=T[chrX:101413096[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	26796701	+	chr5	26801897	+	.	61	53	3309059_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=3309059_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_5_26778501_26803501_344C;SPAN=5196;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:134 GQ:39.8 PL:[284.0, 0.0, 39.8] SR:53 DR:61 LR:-294.3 LO:294.3);ALT=T[chr5:26801897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	27173645	-	chr6	106832766	+	.	16	13	3311107_1	63.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=CAGTCTCTTTCAAAATCTCTGCTA;MAPQ=60;MATEID=3311107_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_5_27170501_27195501_15C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:108 GQ:63.2 PL:[63.2, 0.0, 198.5] SR:13 DR:16 LR:-63.17 LO:67.09);ALT=[chr6:106832766[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	27936330	+	chr5	27900870	+	.	42	22	3315844_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGAA;MAPQ=60;MATEID=3315844_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_27881001_27906001_89C;SPAN=35460;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:100 GQ:99 PL:[137.9, 0.0, 104.9] SR:22 DR:42 LR:-138.2 LO:138.2);ALT=]chr5:27936330]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	128537737	+	chr6	107321881	+	.	10	0	5279539_1	27.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5279539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:107321881(-)-7:128537737(+)__7_128527001_128552001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:20 GQ:20.9 PL:[27.5, 0.0, 20.9] SR:0 DR:10 LR:-27.64 LO:27.64);ALT=]chr7:128537737]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	108031342	+	chr6	108032403	+	TCCTCCCACTCACTCC	0	56	4349769_1	99.0	.	EVDNC=ASSMB;INSERTION=TCCTCCCACTCACTCC;MAPQ=60;MATEID=4349769_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_6_108020501_108045501_167C;SPAN=1061;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:56 DP:19 GQ:15 PL:[165.0, 15.0, 0.0] SR:56 DR:0 LR:-165.0 LO:165.0);ALT=T[chr6:108032403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	108906232	-	chr11	103792589	+	.	24	24	7166328_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=0;MATEID=7166328_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_103782001_103807001_321C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:31 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:24 DR:24 LR:-125.4 LO:125.4);ALT=[chr11:103792589[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	108906546	+	chr11	103792604	-	.	24	34	4351851_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=0;MATEID=4351851_2;MATENM=2;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_6_108902501_108927501_31C;SECONDARY;SPAN=-1;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:51 DP:42 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:34 DR:24 LR:-148.5 LO:148.5);ALT=T]chr11:103792604];VARTYPE=BND:TRX-hh;JOINTYPE=hh
