chr4	74431940	+	chr4	74454535	-	.	10	0	2753872_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2753872_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:74431940(+)-4:74454535(+)__4_74431001_74456001D;SPAN=22595;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:0 DR:10 LR:-26.24 LO:26.3);ALT=T]chr4:74454535];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	74431980	+	chr4	74480197	+	TAATTATTGTTAATCTATATTGAATGCTTACTATTTTCAGGG	57	88	2754048_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CA;INSERTION=TAATTATTGTTAATCTATATTGAATGCTTACTATTTTCAGGG;MAPQ=60;MATEID=2754048_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_4_74480001_74505001_203C;SECONDARY;SPAN=48217;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:129 DP:15 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:88 DR:57 LR:-382.9 LO:382.9);ALT=A[chr4:74480197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	74454436	-	chr4	74480197	+	.	10	71	2754050_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CA;MAPQ=60;MATEID=2754050_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_4_74480001_74505001_203C;SPAN=25761;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:15 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:71 DR:10 LR:-208.0 LO:208.0);ALT=[chr4:74480197[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	74742064	+	chr4	74744700	+	.	2	5	2754382_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGCA;MAPQ=60;MATEID=2754382_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTTGTT;SCTG=c_4_74725001_74750001_181C;SPAN=2636;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:66 GQ:4.6 PL:[0.0, 4.6, 127.4] SR:5 DR:2 LR:4.871 LO:5.612);ALT=G[chr4:74744700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
