chr3	8325639	+	chr3	8326812	+	.	46	26	1278472_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1278472_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_8305501_8330501_69C;SPAN=1173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:11 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:26 DR:46 LR:-174.9 LO:174.9);ALT=A[chr3:8326812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
