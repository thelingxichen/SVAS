chr11	8933472	-	chr11	8934595	+	.	11	0	4752356_1	16.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4752356_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:8933472(-)-11:8934595(-)__11_8918001_8943001D;SPAN=1123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:0 DR:11 LR:-16.26 LO:23.36);ALT=[chr11:8934595[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	8983732	+	chr11	8985756	+	.	0	10	4752467_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4752467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_8967001_8992001_248C;SPAN=2024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:10 DR:0 LR:-7.543 LO:19.68);ALT=T[chr11:8985756[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	9300106	-	chr11	9301571	+	.	9	0	4753548_1	9.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=4753548_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:9300106(-)-11:9301571(-)__11_9285501_9310501D;SPAN=1465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:0 DR:9 LR:-9.661 LO:18.26);ALT=[chr11:9301571[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	9525796	+	chr11	9526800	+	.	71	32	4754820_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=TGAGCCACCA;MAPQ=60;MATEID=4754820_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_9506001_9531001_317C;SPAN=1004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:37 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:32 DR:71 LR:-270.7 LO:270.7);ALT=A[chr11:9526800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	9685827	+	chr11	9715691	+	.	10	10	4755335_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4755335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_9677501_9702501_209C;SPAN=29864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:48 GQ:29.9 PL:[29.9, 0.0, 86.0] SR:10 DR:10 LR:-29.91 LO:31.44);ALT=T[chr11:9715691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10251848	-	chr11	10363271	+	.	22	0	4757117_1	62.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=4757117_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:10251848(-)-11:10363271(-)__11_10363501_10388501D;SPAN=111423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:0 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:0 DR:22 LR:-62.72 LO:62.72);ALT=[chr11:10363271[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	10260049	+	chr11	10261314	+	.	78	75	4757027_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4757027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_10241001_10266001_335C;SPAN=1265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:37 GQ:33 PL:[363.0, 33.0, 0.0] SR:75 DR:78 LR:-363.1 LO:363.1);ALT=T[chr11:10261314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10292746	+	chr11	10293835	+	.	97	55	4757052_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CAGCAATCTTGATTCTTT;MAPQ=60;MATEID=4757052_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_10290001_10315001_213C;SPAN=1089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:37 GQ:33 PL:[363.0, 33.0, 0.0] SR:55 DR:97 LR:-363.1 LO:363.1);ALT=T[chr11:10293835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10546922	+	chr11	10552190	+	.	3	4	4757773_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4757773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_10535001_10560001_318C;SPAN=5268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:75 GQ:3.6 PL:[0.0, 3.6, 188.1] SR:4 DR:3 LR:3.814 LO:8.777);ALT=T[chr11:10552190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10552298	+	chr11	10555563	+	.	2	16	4757783_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4757783_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_10535001_10560001_362C;SPAN=3265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:97 GQ:29.9 PL:[29.9, 0.0, 204.8] SR:16 DR:2 LR:-29.84 LO:37.44);ALT=T[chr11:10555563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10555775	+	chr11	10562668	+	.	21	0	4757791_1	60.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4757791_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:10555775(+)-11:10562668(-)__11_10535001_10560001D;SPAN=6893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:34 GQ:20.6 PL:[60.2, 0.0, 20.6] SR:0 DR:21 LR:-61.05 LO:61.05);ALT=A[chr11:10562668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10773006	+	chr11	10774217	+	.	0	6	4758136_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=4758136_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_10755501_10780501_92C;SPAN=1211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:6 DR:0 LR:3.764 LO:10.62);ALT=T[chr11:10774217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10819430	+	chr11	10820537	+	.	24	8	4758431_1	72.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4758431_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_10804501_10829501_355C;SPAN=1107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:73 GQ:72.8 PL:[72.8, 0.0, 102.5] SR:8 DR:24 LR:-72.65 LO:72.97);ALT=T[chr11:10820537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	10828966	+	chr11	10830406	+	.	10	0	4758642_1	13.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4758642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:10828966(+)-11:10830406(-)__11_10829001_10854001D;SPAN=1440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:0 DR:10 LR:-12.96 LO:20.79);ALT=A[chr11:10830406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	11822988	+	chr11	11824631	+	GGTTC	108	66	4761109_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GGTTC;MAPQ=60;MATEID=4761109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_11809001_11834001_256C;SPAN=1643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:55 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:66 DR:108 LR:-392.8 LO:392.8);ALT=A[chr11:11824631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	11863771	+	chr11	11901722	+	.	0	9	4761296_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4761296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_11882501_11907501_70C;SPAN=37951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:9 DR:0 LR:-21.31 LO:22.09);ALT=G[chr11:11901722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
