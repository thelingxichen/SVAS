chr2	112638432	+	chr2	112641519	+	.	13	8	946585_1	33.0	.	DISC_MAPQ=19;EVDNC=ASDIS;HOMSEQ=CTGTAT;MAPQ=60;MATEID=946585_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_112626501_112651501_404C;SPAN=3087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:8 DR:13 LR:-33.63 LO:38.73);ALT=T[chr2:112641519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	113342227	+	chr2	113343551	+	.	0	6	949027_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=949027_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_113337001_113362001_339C;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:122 GQ:12.9 PL:[0.0, 12.9, 320.1] SR:6 DR:0 LR:13.25 LO:9.719);ALT=G[chr2:113343551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	113343943	+	chr2	113346441	+	.	4	55	949035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=949035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_113337001_113362001_319C;SPAN=2498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:108 GQ:99 PL:[162.2, 0.0, 99.5] SR:55 DR:4 LR:-163.0 LO:163.0);ALT=G[chr2:113346441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	113591154	+	chr2	113593760	+	TCATCTGTTTAGGGCCATCAGCTTCAAAGAACAAGTCATCCTCATTGCCA	0	15	949726_1	27.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTGTAATAA;INSERTION=TCATCTGTTTAGGGCCATCAGCTTCAAAGAACAAGTCATCCTCATTGCCA;MAPQ=60;MATEID=949726_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_113582001_113607001_223C;SPAN=2606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:81 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:15 DR:0 LR:-27.57 LO:33.43);ALT=T[chr2:113593760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	113591193	+	chr2	113594294	+	.	17	0	949727_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=949727_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:113591193(+)-2:113594294(-)__2_113582001_113607001D;SPAN=3101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:94 GQ:30.8 PL:[30.8, 0.0, 195.8] SR:0 DR:17 LR:-30.65 LO:37.69);ALT=T[chr2:113594294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114151301	+	chr2	114153615	+	.	16	0	951320_1	39.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=951320_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:114151301(+)-2:114153615(-)__2_114145501_114170501D;SPAN=2314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:0 DR:16 LR:-39.54 LO:40.27);ALT=T[chr2:114153615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114647821	+	chr2	114670747	+	.	26	0	953560_1	63.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=953560_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:114647821(+)-2:114670747(-)__2_114635501_114660501D;SPAN=22926;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:83 GQ:63.5 PL:[63.5, 0.0, 136.1] SR:0 DR:26 LR:-63.34 LO:64.87);ALT=A[chr2:114670747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114647903	+	chr2	114674461	+	TACAAAACTAGGATATGCTGGAAATACAGAACCACAGTTTATCATCCCTTCCT	25	74	953563_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GTA;INSERTION=TACAAAACTAGGATATGCTGGAAATACAGAACCACAGTTTATCATCCCTTCCT;MAPQ=60;MATEID=953563_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_114635501_114660501_55C;SPAN=26558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:50 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:74 DR:25 LR:-250.9 LO:250.9);ALT=A[chr2:114674461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114674585	+	chr2	114684920	+	.	2	20	953734_1	59.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=953734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_114684501_114709501_327C;SPAN=10335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:49 GQ:59.3 PL:[59.3, 0.0, 59.3] SR:20 DR:2 LR:-59.35 LO:59.35);ALT=G[chr2:114684920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114688974	+	chr2	114691854	+	.	0	9	953749_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=953749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_114684501_114709501_316C;SPAN=2880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:63 GQ:12.8 PL:[12.8, 0.0, 138.2] SR:9 DR:0 LR:-12.64 LO:18.94);ALT=G[chr2:114691854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114697680	+	chr2	114699761	+	.	2	6	953772_1	7.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=953772_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_114684501_114709501_301C;SPAN=2081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:6 DR:2 LR:-6.901 LO:15.9);ALT=G[chr2:114699761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114699936	+	chr2	114709054	+	.	8	7	953780_1	18.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=953780_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_114684501_114709501_336C;SPAN=9118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:7 DR:8 LR:-18.7 LO:24.04);ALT=G[chr2:114709054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114699975	+	chr2	114709294	+	.	9	0	953781_1	12.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=953781_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:114699975(+)-2:114709294(-)__2_114684501_114709501D;SPAN=9319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=A[chr2:114709294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114709148	+	chr2	114714936	+	AATATTGTCCTCTCTGGAGGTTCAACCATGTTCAGGGACTTTGGACGTCGCTTGCAAAGAGATTTGAAAAGAACTGTAGATGCCCGGCTGAAATTAAGTGAGGAATTGAGTGGTGGTAGATTGAAGCCAAAACCTATTGATGTACAAGTCATTACACACCACATGCAGCGATATGCAGTTTGGTTTGGAGGATCAATGCTGGCTTCCAC	0	25	953795_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATATTGTCCTCTCTGGAGGTTCAACCATGTTCAGGGACTTTGGACGTCGCTTGCAAAGAGATTTGAAAAGAACTGTAGATGCCCGGCTGAAATTAAGTGAGGAATTGAGTGGTGGTAGATTGAAGCCAAAACCTATTGATGTACAAGTCATTACACACCACATGCAGCGATATGCAGTTTGGTTTGGAGGATCAATGCTGGCTTCCAC;MAPQ=60;MATEID=953795_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_114684501_114709501_351C;SPAN=5788;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:36 GQ:13.4 PL:[72.8, 0.0, 13.4] SR:25 DR:0 LR:-74.96 LO:74.96);ALT=G[chr2:114714936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114709422	+	chr2	114713198	+	.	2	14	953677_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=18;MATEID=953677_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_114709001_114734001_328C;SPAN=3776;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:14 DR:2 LR:-26.17 LO:31.35);ALT=G[chr2:114713198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	114713283	+	chr2	114714936	+	.	6	12	953688_1	35.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=953688_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_114709001_114734001_328C;SPAN=1653;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:76 GQ:35.6 PL:[35.6, 0.0, 147.8] SR:12 DR:6 LR:-35.53 LO:39.47);ALT=G[chr2:114714936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
