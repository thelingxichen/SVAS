chr21	14816840	+	chr21	14818167	+	AAGTGCTACTACT	45	28	7114665_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;INSERTION=AAGTGCTACTACT;MAPQ=60;MATEID=7114665_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_21_14798001_14823001_224C;SPAN=1327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:39 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:28 DR:45 LR:-181.5 LO:181.5);ALT=T[chr21:14818167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	14889907	+	chr21	14888793	+	.	11	0	7114975_1	17.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=7114975_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:14888793(-)-21:14889907(+)__21_14871501_14896501D;SPAN=1114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=]chr21:14889907]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	15460780	+	chr21	15461865	+	AATAATTCATATA	0	7	7116682_1	13.0	.	EVDNC=ASSMB;INSERTION=AATAATTCATATA;MAPQ=60;MATEID=7116682_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_21_15459501_15484501_285C;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:37 GQ:13.1 PL:[13.1, 0.0, 75.8] SR:7 DR:0 LR:-13.08 LO:15.67);ALT=T[chr21:15461865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	15893586	+	chr21	15918531	+	.	24	0	7117587_1	69.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7117587_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:15893586(+)-21:15918531(-)__21_15900501_15925501D;SPAN=24945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:35 GQ:13.7 PL:[69.8, 0.0, 13.7] SR:0 DR:24 LR:-71.71 LO:71.71);ALT=T[chr21:15918531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
