chrX	10738666	+	chrX	10788675	+	.	34	2	7364014_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GATCACCTATTGAAAAATATGTTATAGTTTTCTGACTAAACTCATCAAGGCTAGTGTTTACGTAGGTAGTC;MAPQ=60;MATEID=7364014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_10780001_10805001_162C;SPAN=50009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:1 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:2 DR:34 LR:-105.6 LO:105.6);ALT=C[chrX:10788675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
