chr1	118087003	+	chr1	117941213	+	ATC	55	43	469955_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=ATC;MAPQ=60;MATEID=469955_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_118065501_118090501_366C;SPAN=145790;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:44 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:43 DR:55 LR:-227.8 LO:227.8);ALT=]chr1:118087003]T;VARTYPE=BND:DUP-th;JOINTYPE=th
