chr19	5488255	+	chr19	5487054	+	.	32	35	10129311_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCCCAGGCTGGAGTGCAGTGGCGC;MAPQ=60;MATEID=10129311_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5463501_5488501_141C;SPAN=1201;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:169 GQ:99 PL:[162.2, 0.0, 248.0] SR:35 DR:32 LR:-162.2 LO:163.2);ALT=]chr19:5488255]G;VARTYPE=BND:DUP-th;JOINTYPE=th
