chr3	170506477	-	chr3	170507590	+	.	10	0	2483139_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2483139_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:170506477(-)-3:170507590(-)__3_170495501_170520501D;SPAN=1113;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:156 GQ:9.1 PL:[0.0, 9.1, 396.0] SR:0 DR:10 LR:9.254 LO:17.38);ALT=[chr3:170507590[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
