chr1	50039956	+	chr1	50148301	+	.	11	10	248643_1	30.0	.	DISC_MAPQ=52;EVDNC=ASDIS;MAPQ=60;MATEID=248643_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_50127001_50152001_6C;SPAN=108345;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:71 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:10 DR:11 LR:-30.28 LO:34.4);ALT=T[chr1:50148301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	50403662	+	chr1	50206695	+	.	3	10	249177_1	19.0	.	DISC_MAPQ=25;EVDNC=TSI_L;HOMSEQ=AGCAGAAGGCAAGAAATAACTA;MAPQ=14;MATEID=249177_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_1_50200501_50225501_20C;SPAN=196967;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:10 DR:3 LR:-19.29 LO:25.9);ALT=]chr1:50403662]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	50763767	-	chr1	50765164	+	.	10	0	251078_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=251078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:50763767(-)-1:50765164(-)__1_50739501_50764501D;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-13.77 LO:20.98);ALT=[chr1:50765164[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	51350985	-	chr9	115594722	+	.	7	15	5968185_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACACACACACACTCTCTCTCTCTCTCTCTC;MAPQ=60;MATEID=5968185_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_9_115591001_115616001_14C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:33 GQ:24.2 PL:[53.9, 0.0, 24.2] SR:15 DR:7 LR:-54.29 LO:54.29);ALT=[chr9:115594722[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	51743372	+	chrX	103003940	+	.	2	8	11335112_1	29.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=CTCCCAAAGTGCTGGGATTACAGGCGTGAGC;MAPQ=43;MATEID=11335112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_102998001_103023001_313C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:10 DP:5 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:8 DR:2 LR:-29.71 LO:29.71);ALT=C[chrX:103003940[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	114898112	+	chr9	114662191	+	.	9	5	5966360_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=5966360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_114880501_114905501_292C;SPAN=235921;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:5 DR:9 LR:-20.5 LO:21.66);ALT=]chr9:114898112]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	103000383	+	chrX	102832619	+	TAATGTACTAACATATAAATATTAAT	0	56	11335128_1	99.0	.	EVDNC=ASSMB;INSERTION=TAATGTACTAACATATAAATATTAAT;MAPQ=60;MATEID=11335128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_102998001_103023001_202C;SPAN=167764;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:56 DP:46 GQ:15 PL:[165.0, 15.0, 0.0] SR:56 DR:0 LR:-165.0 LO:165.0);ALT=]chrX:103000383]T;VARTYPE=BND:DUP-th;JOINTYPE=th
