chr1	77672467	+	chr1	77685033	+	.	11	0	209553_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=209553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:77672467(+)-1:77685033(-)__1_77665001_77690001D;SPAN=12566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:0 DR:11 LR:-16.53 LO:23.43);ALT=G[chr1:77685033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	77685338	+	chr1	77686471	+	.	6	3	209574_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=209574_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_77665001_77690001_205C;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:61 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:3 DR:6 LR:-6.581 LO:14.02);ALT=G[chr1:77686471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	78207479	+	chr1	78225406	+	.	15	0	211109_1	31.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=211109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:78207479(+)-1:78225406(-)__1_78204001_78229001D;SPAN=17927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:68 GQ:31.1 PL:[31.1, 0.0, 133.4] SR:0 DR:15 LR:-31.09 LO:34.72);ALT=A[chr1:78225406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	78409956	+	chr1	78411191	+	.	0	5	211631_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=211631_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_78400001_78425001_157C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:5 DR:0 LR:5.711 LO:8.577);ALT=T[chr1:78411191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	78422387	+	chr1	78425869	+	.	5	6	211975_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=211975_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_78424501_78449501_95C;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:6 DR:5 LR:-13.67 LO:17.51);ALT=T[chr1:78425869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	78426180	+	chr1	78428454	+	.	14	7	211981_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=211981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_78424501_78449501_384C;SPAN=2274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:75 GQ:39.2 PL:[39.2, 0.0, 141.5] SR:7 DR:14 LR:-39.1 LO:42.43);ALT=C[chr1:78428454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	78435701	+	chr1	78444569	+	.	0	10	212007_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=212007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_78424501_78449501_182C;SPAN=8868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:10 DR:0 LR:-14.59 LO:21.18);ALT=T[chr1:78444569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	79115609	+	chr1	79120698	+	.	10	0	213370_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=213370_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:79115609(+)-1:79120698(-)__1_79110501_79135501D;SPAN=5089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:0 DR:10 LR:-12.69 LO:20.72);ALT=T[chr1:79120698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	133815668	+	chr1	79276448	+	.	13	0	2216195_1	32.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=2216195_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:79276448(-)-4:133815668(+)__4_133794501_133819501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:39 GQ:32.3 PL:[32.3, 0.0, 62.0] SR:0 DR:13 LR:-32.35 LO:32.87);ALT=]chr4:133815668]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	80221782	+	chr1	80223029	+	.	5	14	215615_1	41.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=215615_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_1_80213001_80238001_249C;SPAN=1247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:43 GQ:41.3 PL:[41.3, 0.0, 61.1] SR:14 DR:5 LR:-41.17 LO:41.42);ALT=T[chr1:80223029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
