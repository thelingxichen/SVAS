chr13	76100778	+	chr13	76111898	+	AAACTGTGGAATCGTCATTTCAAAGCACTTGGTCTTTACTTGGCCTGAATGATCTGCCACTTTTAGCATCACTGCAACGTAAGGATACTTAAGAGATCTGCAAGTGTCTGAGCTCACAGCCATACCCAGTTTCCACTGAAAATCTACAAGCTGGTTGGTG	26	138	5558341_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=AAACTGTGGAATCGTCATTTCAAAGCACTTGGTCTTTACTTGGCCTGAATGATCTGCCACTTTTAGCATCACTGCAACGTAAGGATACTTAAGAGATCTGCAAGTGTCTGAGCTCACAGCCATACCCAGTTTCCACTGAAAATCTACAAGCTGGTTGGTG;MAPQ=60;MATEID=5558341_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_76097001_76122001_110C;SPAN=11120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:149 DP:177 GQ:14.8 PL:[458.8, 14.8, 0.0] SR:138 DR:26 LR:-475.2 LO:475.2);ALT=G[chr13:76111898[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	76100778	+	chr13	76104250	+	.	4	107	5558340_1	99.0	.	DISC_MAPQ=45;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5558340_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_13_76097001_76122001_110C;SPAN=3472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:259 GQ:99 PL:[296.3, 0.0, 332.6] SR:107 DR:4 LR:-296.2 LO:296.4);ALT=G[chr13:76104250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	76104547	+	chr13	76111900	+	.	78	0	5558358_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5558358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:76104547(+)-13:76111900(-)__13_76097001_76122001D;SPAN=7353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:96 GQ:0.5 PL:[231.5, 0.0, 0.5] SR:0 DR:78 LR:-245.5 LO:245.5);ALT=A[chr13:76111900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	76124000	+	chr13	76134884	+	CACCA	16	3	5558184_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CACCA;MAPQ=60;MATEID=5558184_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_76121501_76146501_305C;SPAN=10884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:102 GQ:32 PL:[32.0, 0.0, 213.5] SR:3 DR:16 LR:-31.78 LO:39.7);ALT=T[chr13:76134884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	76124000	+	chr13	76140828	+	.	8	0	5558185_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5558185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:76124000(+)-13:76140828(-)__13_76121501_76146501D;SPAN=16828;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:116 GQ:4.8 PL:[0.0, 4.8, 290.4] SR:0 DR:8 LR:5.019 LO:14.16);ALT=T[chr13:76140828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	76135017	+	chr13	76140829	+	.	0	9	5558219_1	6.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5558219_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_76121501_76146501_274C;SPAN=5812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:9 DR:0 LR:-6.139 LO:17.59);ALT=G[chr13:76140829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
