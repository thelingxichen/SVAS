chr1	29026716	-	chr1	29027878	+	.	8	0	150177_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=150177_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:29026716(-)-1:29027878(-)__1_29008001_29033001D;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:162 GQ:17.2 PL:[0.0, 17.2, 425.8] SR:0 DR:8 LR:17.48 LO:12.97);ALT=[chr1:29027878[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
