chr9	71650863	+	chr9	71661301	+	.	14	16	4259556_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4259556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_71638001_71663001_78C;SPAN=10438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:102 GQ:48.5 PL:[48.5, 0.0, 197.0] SR:16 DR:14 LR:-48.29 LO:53.49);ALT=A[chr9:71661301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	71661398	+	chr9	71668055	+	.	0	19	4259609_1	48.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=25;MATEID=4259609_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_71638001_71663001_227C;SPAN=6657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:53 GQ:48.5 PL:[48.5, 0.0, 78.2] SR:19 DR:0 LR:-48.36 LO:48.79);ALT=G[chr9:71668055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	71738122	+	chr9	71743355	+	.	46	35	4259850_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=4259850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_71736001_71761001_363C;SPAN=5233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:58 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:35 DR:46 LR:-184.8 LO:184.8);ALT=C[chr9:71743355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	72373620	+	chr9	72374765	+	.	0	15	4262447_1	21.0	.	EVDNC=ASSMB;HOMSEQ=TCAC;MAPQ=60;MATEID=4262447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_72373001_72398001_336C;SPAN=1145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:103 GQ:21.8 PL:[21.8, 0.0, 226.4] SR:15 DR:0 LR:-21.61 LO:31.71);ALT=C[chr9:72374765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	72860526	+	chr9	72854182	+	.	11	0	4264040_1	16.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=4264040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:72854182(-)-9:72860526(+)__9_72838501_72863501D;SPAN=6344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:0 DR:11 LR:-15.99 LO:23.29);ALT=]chr9:72860526]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	72874179	+	chr9	72879220	+	.	0	12	4263644_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4263644_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_72863001_72888001_101C;SPAN=5041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:101 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:12 DR:0 LR:-12.25 LO:24.22);ALT=T[chr9:72879220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	72892389	+	chr9	72893405	+	.	0	4	4263854_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4263854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_72887501_72912501_253C;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:98 GQ:13.2 PL:[0.0, 13.2, 264.0] SR:4 DR:0 LR:13.35 LO:6.151);ALT=G[chr9:72893405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	72895816	+	chr9	72897337	+	.	0	8	4263870_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4263870_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_72887501_72912501_114C;SPAN=1521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:8 DR:0 LR:-0.1283 LO:14.81);ALT=G[chr9:72897337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
