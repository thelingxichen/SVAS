chr2	1536483	+	chr2	1529454	+	.	38	23	895065_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CCCCAAATCCCCC;MAPQ=48;MATEID=895065_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_1519001_1544001_59C;SPAN=7029;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:31 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:23 DR:38 LR:-174.9 LO:174.9);ALT=]chr2:1536483]C;VARTYPE=BND:DUP-th;JOINTYPE=th
