chr1	71447114	+	chr6	157944020	+	.	0	26	4463136_1	75.0	.	EVDNC=ASSMB;HOMSEQ=TTTCTTTTCTTT;MAPQ=60;MATEID=4463136_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_157927001_157952001_164C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:26 DP:9 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:26 DR:0 LR:-75.92 LO:75.92);ALT=T[chr6:157944020[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	157559511	+	chr6	157641364	-	.	32	0	4462263_1	92.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4462263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:157559511(+)-6:157641364(+)__6_157633001_157658001D;SPAN=81853;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:32 DP:0 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=N]chr6:157641364];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	157734424	+	chr6	157733133	+	.	7	26	4462993_1	71.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=CTCACC;MAPQ=19;MATEID=4462993_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_6_157731001_157756001_129C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:140 GQ:71 PL:[71.0, 0.0, 269.0] SR:26 DR:7 LR:-71.0 LO:77.48);ALT=]chr6:157734424]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	158908130	+	chr12	117819265	-	.	12	0	4465288_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4465288_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:158908130(+)-12:117819265(+)__6_158907001_158932001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=A]chr12:117819265];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	117086884	+	chr12	117088194	+	.	148	67	7847408_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGTGGCTCAGGCCTATAATCCCAGCACTT;MAPQ=60;MATEID=7847408_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_12_117085501_117110501_372C;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:187 DP:29 GQ:50.5 PL:[554.5, 50.5, 0.0] SR:67 DR:148 LR:-554.5 LO:554.5);ALT=T[chr12:117088194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
