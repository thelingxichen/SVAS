chr12	90687033	+	chr12	90363383	+	.	79	59	7789402_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCTAGG;MAPQ=60;MATEID=7789402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_90674501_90699501_123C;SPAN=323650;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:53 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:59 DR:79 LR:-313.6 LO:313.6);ALT=]chr12:90687033]G;VARTYPE=BND:DUP-th;JOINTYPE=th
