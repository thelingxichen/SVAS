chr4	122604633	+	chr4	122605831	+	.	0	8	2180641_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2180641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_122598001_122623001_58C;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:8 DR:0 LR:2.31 LO:14.49);ALT=C[chr4:122605831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	122605927	+	chr4	122607442	+	.	0	14	2180651_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2180651_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_122598001_122623001_348C;SPAN=1515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:116 GQ:14.9 PL:[14.9, 0.0, 265.7] SR:14 DR:0 LR:-14.79 LO:28.36);ALT=C[chr4:122607442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	122605975	+	chr4	122618040	+	.	10	0	2180652_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2180652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:122605975(+)-4:122618040(-)__4_122598001_122623001D;SPAN=12065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:114 GQ:2.3 PL:[2.3, 0.0, 272.9] SR:0 DR:10 LR:-2.125 LO:18.79);ALT=T[chr4:122618040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	122607584	+	chr4	122618048	+	.	23	0	2180664_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2180664_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:122607584(+)-4:122618048(-)__4_122598001_122623001D;SPAN=10464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:99 GQ:49.1 PL:[49.1, 0.0, 191.0] SR:0 DR:23 LR:-49.1 LO:53.83);ALT=T[chr4:122618048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	123301080	+	chr4	123302205	-	.	2	3	2183060_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=2183060_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_123284001_123309001_136C;SPAN=1125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:90 GQ:7.8 PL:[0.0, 7.8, 234.3] SR:3 DR:2 LR:7.878 LO:8.37);ALT=G]chr4:123302205];VARTYPE=BND:INV-hh;JOINTYPE=hh
