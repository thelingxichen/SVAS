chr3	177294510	+	chr3	177297474	+	.	56	42	1806591_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1806591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_177282001_177307001_340C;SPAN=2964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:76 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:42 DR:56 LR:-247.6 LO:247.6);ALT=A[chr3:177297474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	177381310	+	chr3	177385458	+	.	25	0	1807092_1	61.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=1807092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:177381310(+)-3:177385458(-)__3_177380001_177405001D;SPAN=4148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:77 GQ:61.7 PL:[61.7, 0.0, 124.4] SR:0 DR:25 LR:-61.66 LO:62.85);ALT=T[chr3:177385458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
