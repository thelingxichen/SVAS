chr22	16853977	+	chr22	16848555	+	.	12	0	10828124_1	0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=10828124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:16848555(-)-22:16853977(+)__22_16831501_16856501D;SPAN=5422;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:12 DP:152 GQ:1.3 PL:[0.0, 1.3, 369.6] SR:0 DR:12 LR:1.569 LO:21.98);ALT=]chr22:16853977]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	17047117	+	chr22	17044030	+	.	9	0	10830473_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=10830473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:17044030(-)-22:17047117(+)__22_17027501_17052501D;SPAN=3087;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:191 GQ:21.7 PL:[0.0, 21.7, 505.0] SR:0 DR:9 LR:22.04 LO:14.41);ALT=]chr22:17047117]A;VARTYPE=BND:DUP-th;JOINTYPE=th
