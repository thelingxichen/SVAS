chr5	83947993	+	chr5	83954951	+	.	14	0	3579483_1	30.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3579483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:83947993(+)-5:83954951(-)__5_83937001_83962001D;SPAN=6958;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:57 GQ:30.8 PL:[30.8, 0.0, 106.7] SR:0 DR:14 LR:-30.77 LO:33.16);ALT=T[chr5:83954951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	84303728	+	chr5	169899776	-	.	3	40	3581223_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATAAAAAGGAATGAATTAACAGCATTTGTAGTGACCTG;MAPQ=60;MATEID=3581223_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_84280001_84305001_13C;SPAN=85596048;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:42 DP:41 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:40 DR:3 LR:-122.1 LO:122.1);ALT=G]chr5:169899776];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	169597468	-	chr5	169598756	+	CTCTG	106	96	3922216_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTCTG;MAPQ=60;MATEID=3922216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_169589001_169614001_381C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:223 DP:133 GQ:60.1 PL:[660.1, 60.1, 0.0] SR:96 DR:106 LR:-660.2 LO:660.2);ALT=[chr5:169598756[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	170129990	+	chr5	170131367	+	.	38	0	3924128_1	99.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=3924128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:170129990(+)-5:170131367(-)__5_170128001_170153001D;SPAN=1377;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:38 DP:48 GQ:3.5 PL:[112.4, 0.0, 3.5] SR:0 DR:38 LR:-118.5 LO:118.5);ALT=G[chr5:170131367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
