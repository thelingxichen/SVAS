chr6	37007057	+	chr6	36996778	+	.	64	60	4142255_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4142255_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_36995001_37020001_292C;SPAN=10279;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:106 DP:149 GQ:52.1 PL:[309.5, 0.0, 52.1] SR:60 DR:64 LR:-320.0 LO:320.0);ALT=]chr6:37007057]G;VARTYPE=BND:DUP-th;JOINTYPE=th
