chrX	42512048	+	chrX	42513870	+	.	22	0	11114875_1	41.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=11114875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:42512048(+)-23:42513870(-)__23_42507501_42532501D;SPAN=1822;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:117 GQ:41 PL:[41.0, 0.0, 242.3] SR:0 DR:22 LR:-40.92 LO:49.2);ALT=A[chrX:42513870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	42512290	+	chrX	42513871	+	.	58	152	11114876_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=45;MATEID=11114876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_42507501_42532501_144C;SPAN=1581;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:187 DP:67 GQ:50.5 PL:[554.5, 50.5, 0.0] SR:152 DR:58 LR:-554.5 LO:554.5);ALT=A[chrX:42513871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
