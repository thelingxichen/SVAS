chr3	3873165	+	chr7	45589198	-	.	9	0	1809085_1	7.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=1809085_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:3873165(+)-7:45589198(+)__3_3871001_3896001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=A]chr7:45589198];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	4066937	+	chr3	4069556	+	.	0	69	1809792_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACAAAATATATAT;MAPQ=60;MATEID=1809792_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_4067001_4092001_227C;SPAN=2619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:13 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:69 DR:0 LR:-204.7 LO:204.7);ALT=T[chr3:4069556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44873537	+	chr7	44545137	+	A	49	22	4757691_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4757691_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_44541001_44566001_320C;SPAN=328400;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:89 GQ:28.7 PL:[187.1, 0.0, 28.7] SR:22 DR:49 LR:-193.8 LO:193.8);ALT=]chr7:44873537]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	44895446	+	chr7	44896478	-	.	8	0	4760099_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4760099_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44895446(+)-7:44896478(+)__7_44884001_44909001D;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:176 GQ:21.1 PL:[0.0, 21.1, 468.7] SR:0 DR:8 LR:21.27 LO:12.68);ALT=T]chr7:44896478];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	45274348	+	chr7	45276143	-	.	2	3	4764581_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGTCTTCCTTTACCTCCCTGAAT;MAPQ=60;MATEID=4764581_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_45276001_45301001_483C;SPAN=1795;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:77 GQ:7.5 PL:[0.0, 7.5, 201.3] SR:3 DR:2 LR:7.657 LO:6.577);ALT=A]chr7:45276143];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	46057422	+	chr7	46056327	+	.	5	2	4769735_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=35;MATEID=4769735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_46035501_46060501_9C;SPAN=1095;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:210 GQ:40.3 PL:[0.0, 40.3, 590.8] SR:2 DR:5 LR:40.39 LO:6.514);ALT=]chr7:46057422]G;VARTYPE=BND:DUP-th;JOINTYPE=th
