chr4	13481152	+	chr4	13485700	+	.	0	9	1907303_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1907303_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_13475001_13500001_100C;SPAN=4548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:52 GQ:15.8 PL:[15.8, 0.0, 108.2] SR:9 DR:0 LR:-15.62 LO:19.77);ALT=T[chr4:13485700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
