chr1	102892536	-	chr1	102970102	+	.	11	0	438234_1	23.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=438234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:102892536(-)-1:102970102(-)__1_102875501_102900501D;SPAN=77566;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:0 DR:11 LR:-23.31 LO:25.67);ALT=[chr1:102970102[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	103096385	+	chr12	2089842	+	.	58	127	7331314_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;MAPQ=0;MATEID=7331314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_2082501_2107501_352C;SPAN=-1;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:174 DP:67 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:127 DR:58 LR:-514.9 LO:514.9);ALT=C[chr12:2089842[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	76526512	+	chr2	76528894	+	.	102	79	1101247_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GTTTTCCATGTTTT;MAPQ=60;MATEID=1101247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_76513501_76538501_242C;SPAN=2382;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:155 DP:34 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:79 DR:102 LR:-458.8 LO:458.8);ALT=T[chr2:76528894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	76773553	+	chr2	76775453	+	TTATTCTTTTA	52	43	1101772_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TTATTCTTTTA;MAPQ=60;MATEID=1101772_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_76758501_76783501_166C;SPAN=1900;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:24 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:43 DR:52 LR:-227.8 LO:227.8);ALT=T[chr2:76775453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	77007953	-	chr2	77023870	+	.	11	0	1104414_1	1.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=1104414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:77007953(-)-2:77023870(-)__2_77003501_77028501D;SPAN=15917;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:128 GQ:1.7 PL:[1.7, 0.0, 308.6] SR:0 DR:11 LR:-1.633 LO:20.57);ALT=[chr2:77023870[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	77316383	+	chr9	118236416	+	.	10	50	1104203_1	99.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=CTTGTCTCTACCCCTTCT;MAPQ=60;MATEID=1104203_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_77297501_77322501_447C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:70 GQ:5.7 PL:[181.5, 5.7, 0.0] SR:50 DR:10 LR:-188.3 LO:188.3);ALT=T[chr9:118236416[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	77632026	+	chr17	35736509	+	.	16	47	1105383_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1105383_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_77616001_77641001_397C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:49 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:47 DR:16 LR:-155.1 LO:155.1);ALT=T[chr17:35736509[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	77841755	+	chr2	77843151	+	.	79	54	1105785_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1105785_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_77836501_77861501_119C;SPAN=1396;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:85 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:54 DR:79 LR:-323.5 LO:323.5);ALT=A[chr2:77843151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	77847438	+	chr2	77851850	+	.	53	46	1105800_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1105800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_77836501_77861501_252C;SPAN=4412;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:78 GQ:21 PL:[231.0, 21.0, 0.0] SR:46 DR:53 LR:-231.1 LO:231.1);ALT=T[chr2:77851850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	138364741	+	chr12	2994185	-	.	69	30	1374378_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=1374378_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_138351501_138376501_67C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:59 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:30 DR:69 LR:-277.3 LO:277.3);ALT=T]chr12:2994185];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	28226476	+	chr3	54428355	+	.	36	0	7504129_1	96.0	.	DISC_MAPQ=7;EVDNC=DSCRD;IMPRECISE;MAPQ=7;MATEID=7504129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:54428355(-)-12:28226476(+)__12_28224001_28249001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:83 GQ:96.5 PL:[96.5, 0.0, 103.1] SR:0 DR:36 LR:-96.35 LO:96.37);ALT=]chr12:28226476]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	54512690	-	chr9	118004803	+	.	13	31	2030286_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TATATATATATAT;MAPQ=60;MATEID=2030286_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_54488001_54513001_188C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:36 DP:27 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:31 DR:13 LR:-105.6 LO:105.6);ALT=[chr9:118004803[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	56607729	+	chr3	56621585	+	.	81	36	2038660_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=2038660_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_56619501_56644501_197C;SPAN=13856;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:43 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:36 DR:81 LR:-310.3 LO:310.3);ALT=A[chr3:56621585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57524041	+	chr3	57522647	+	CTATGATTAGTGA	16	35	2043473_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;INSERTION=CTATGATTAGTGA;MAPQ=60;MATEID=2043473_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57501501_57526501_335C;SPAN=1394;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:43 DP:120 GQ:99 PL:[109.4, 0.0, 182.0] SR:35 DR:16 LR:-109.4 LO:110.4);ALT=]chr3:57524041]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	57522710	+	chr3	57524052	+	ATAATCACCTGA	0	33	2043474_1	74.0	.	EVDNC=ASSMB;INSERTION=ATAATCACCTGA;MAPQ=60;MATEID=2043474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57501501_57526501_170C;SPAN=1342;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:126 GQ:74.9 PL:[74.9, 0.0, 230.0] SR:33 DR:0 LR:-74.8 LO:79.24);ALT=T[chr3:57524052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57991849	+	chr17	35587296	-	.	8	0	2046259_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2046259_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:57991849(+)-17:35587296(+)__3_57967001_57992001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=G]chr17:35587296];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	58946234	+	chr21	47677372	+	.	11	13	10818311_1	62.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=CAGCAAGGCTCTGTCTCAAAAAAAAAAAAAAAAA;MAPQ=35;MATEID=10818311_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_21_47677001_47702001_387C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:22 DP:13 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:13 DR:11 LR:-62.72 LO:62.72);ALT=A[chr21:47677372[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	59763595	+	chr3	59746779	+	.	3	6	2053484_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2053484_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_59755501_59780501_273C;SPAN=16816;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:69 GQ:7.7 PL:[7.7, 0.0, 159.5] SR:6 DR:3 LR:-7.714 LO:16.06);ALT=]chr3:59763595]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	60123979	+	chr3	60352336	+	.	86	58	2055193_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGATG;MAPQ=60;MATEID=2055193_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_60343501_60368501_77C;SPAN=228357;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:13 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:58 DR:86 LR:-333.4 LO:333.4);ALT=G[chr3:60352336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60276268	+	chr3	60389793	+	.	51	35	2055187_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGG;MAPQ=60;MATEID=2055187_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_60368001_60393001_25C;SPAN=113525;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:9 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:35 DR:51 LR:-211.3 LO:211.3);ALT=G[chr3:60389793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60363255	+	chr3	60667236	+	.	9	0	2055447_1	20.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2055447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:60363255(+)-3:60667236(-)__3_60662001_60687001D;SPAN=303981;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:35 GQ:20.3 PL:[20.3, 0.0, 63.2] SR:0 DR:9 LR:-20.23 LO:21.53);ALT=C[chr3:60667236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60363538	+	chr3	60667237	+	.	10	30	2055448_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=52;MATEID=2055448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_60662001_60687001_399C;SPAN=303699;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:30 DR:10 LR:-102.3 LO:102.3);ALT=T[chr3:60667237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60412920	+	chr3	60532343	+	.	0	35	2055252_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2055252_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_3_60392501_60417501_18C;SPAN=119423;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:6 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:35 DR:0 LR:-102.3 LO:102.3);ALT=T[chr3:60532343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60587837	+	chr3	60655441	+	C	70	46	2055290_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=2055290_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_60564001_60589001_222C;SPAN=67604;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:9 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:46 DR:70 LR:-277.3 LO:277.3);ALT=C[chr3:60655441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	61069019	-	chr4	86099305	+	.	11	37	2056871_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;MAPQ=13;MATEID=2056871_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_61054001_61079001_409C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:121 GQ:99 PL:[112.7, 0.0, 178.7] SR:37 DR:11 LR:-112.5 LO:113.3);ALT=[chr4:86099305[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr17	35071989	+	chr7	147472325	+	.	6	25	9620322_1	89.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=ATATATATATTTATATATAT;MAPQ=60;MATEID=9620322_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_17_35059501_35084501_198C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:31 DP:23 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:25 DR:6 LR:-89.12 LO:89.12);ALT=]chr17:35071989]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	148072866	+	chr7	148076324	+	.	41	55	5319441_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=ATC;MAPQ=60;MATEID=5319441_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_148053501_148078501_60C;SPAN=3458;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:21 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:55 DR:41 LR:-227.8 LO:227.8);ALT=C[chr7:148076324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	117082012	+	chr9	117083382	+	.	91	47	5971666_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=5971666_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_117061001_117086001_8C;SPAN=1370;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:112 DP:23 GQ:30 PL:[330.0, 30.0, 0.0] SR:47 DR:91 LR:-330.1 LO:330.1);ALT=G[chr9:117083382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	1730110	-	chr17	36594951	+	.	35	43	7329119_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGGCGTGGTGGCTCACACCTGTAATGCCAGCACTTTGGGAGGTTGAGGCGGGC;MAPQ=60;MATEID=7329119_2;MATENM=3;NM=2;NUMPARTS=2;SCTG=c_12_1715001_1740001_19C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:89 GQ:10.8 PL:[237.6, 10.8, 0.0] SR:43 DR:35 LR:-243.8 LO:243.8);ALT=[chr17:36594951[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	3837747	+	chr12	3451947	+	CA	60	28	7339259_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CA;MAPQ=60;MATEID=7339259_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_3430001_3455001_68C;SPAN=385800;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:91 GQ:4.5 PL:[227.7, 4.5, 0.0] SR:28 DR:60 LR:-237.3 LO:237.3);ALT=]chr12:3837747]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	27861632	+	chr12	27668868	+	.	37	16	7500094_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=7500094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_27856501_27881501_257C;SPAN=192764;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:100 GQ:99 PL:[118.1, 0.0, 124.7] SR:16 DR:37 LR:-118.2 LO:118.2);ALT=]chr12:27861632]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	28026953	+	chr15	84491260	-	.	9	0	7501673_1	4.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=7501673_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:28026953(+)-15:84491260(+)__12_28003501_28028501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:93 GQ:4.7 PL:[4.7, 0.0, 219.2] SR:0 DR:9 LR:-4.513 LO:17.32);ALT=C]chr15:84491260];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	28027143	-	chr15	84491119	+	.	22	0	7501675_1	50.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=7501675_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:28027143(-)-15:84491119(-)__12_28003501_28028501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:80 GQ:50.9 PL:[50.9, 0.0, 143.3] SR:0 DR:22 LR:-50.95 LO:53.38);ALT=[chr15:84491119[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr17	2719930	+	chr17	2721218	+	.	104	117	9473625_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=9473625_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_2719501_2744501_295C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:184 DP:37 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:117 DR:104 LR:-544.6 LO:544.6);ALT=T[chr17:2721218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3063342	+	chr17	37133744	+	CACACACATATGTATATATATACACACATATGTATACAC	4	96	9475546_1	99.0	.	DISC_MAPQ=48;EVDNC=TSI_L;INSERTION=CACACACATATGTATATATATACACACATATGTATACAC;MAPQ=60;MATEID=9475546_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACACACA;SCTG=c_17_3062501_3087501_119C;SPAN=34070402;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:56 GQ:26.1 PL:[175.6, 26.1, 0.0] SR:96 DR:4 LR:-175.6 LO:175.6);ALT=T[chr17:37133744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	37133794	+	chr17	3063358	+	TATGTATAT	6	63	9475547_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=TATGTATAT;MAPQ=60;MATEID=9475547_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_3062501_3087501_119C;SPAN=34070436;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:51 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:63 DR:6 LR:-204.7 LO:204.7);ALT=]chr17:37133794]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	3510197	-	chr17	3512185	+	.	8	0	9476900_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=9476900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:3510197(-)-17:3512185(-)__17_3503501_3528501D;SPAN=1988;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:0 DR:8 LR:5.561 LO:14.1);ALT=[chr17:3512185[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	3734815	+	chr17	3735843	+	.	95	81	9478145_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TGAACCCGGGAGGCGGAGGTTGCAGTGAGCC;MAPQ=60;MATEID=9478145_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_17_3724001_3749001_30C;SPAN=1028;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:170 DP:23 GQ:46 PL:[505.0, 46.0, 0.0] SR:81 DR:95 LR:-505.0 LO:505.0);ALT=C[chr17:3735843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36172710	+	chr17	36015933	+	.	8	0	9626540_1	9.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=9626540_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:36015933(-)-17:36172710(+)__17_36162001_36187001D;SPAN=156777;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:0 DR:8 LR:-9.34 LO:16.4);ALT=]chr17:36172710]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	36524997	+	chr17	36526080	+	G	0	58	9629620_1	99.0	.	EVDNC=ASSMB;INSERTION=G;MAPQ=60;MATEID=9629620_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36505001_36530001_176C;SPAN=1083;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:165 GQ:99 PL:[146.9, 0.0, 252.5] SR:58 DR:0 LR:-146.8 LO:148.3);ALT=A[chr17:36526080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
