chr15	23671476	+	chr15	23675251	+	.	54	0	8785674_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=8785674_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:23671476(+)-15:23675251(-)__15_23667001_23692001D;SPAN=3775;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:54 DP:123 GQ:99 PL:[145.1, 0.0, 151.7] SR:0 DR:54 LR:-144.9 LO:144.9);ALT=G[chr15:23675251[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	24613911	+	chr15	24508056	+	.	8	0	8789025_1	8.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=8789025_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:24508056(-)-15:24613911(+)__15_24500001_24525001D;SPAN=105855;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=]chr15:24613911]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	24587511	+	chr15	24802174	-	.	4	6	8789664_1	8.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=8789664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_24573501_24598501_0C;SPAN=214663;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:6 DR:4 LR:-8.306 LO:17.99);ALT=C]chr15:24802174];VARTYPE=BND:INV-hh;JOINTYPE=hh
