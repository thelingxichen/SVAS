chr13	90862855	+	chr13	90864807	+	.	37	25	5593260_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAT;MAPQ=60;MATEID=5593260_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_90846001_90871001_285C;SPAN=1952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:59 GQ:2.7 PL:[148.5, 2.7, 0.0] SR:25 DR:37 LR:-155.5 LO:155.5);ALT=T[chr13:90864807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
