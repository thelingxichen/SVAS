chr2	125051756	+	chr2	125053240	-	.	59	57	1314546_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1314546_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_125048001_125073001_155C;SPAN=1484;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:124 GQ:12.8 PL:[286.7, 0.0, 12.8] SR:57 DR:59 LR:-301.4 LO:301.4);ALT=C]chr2:125053240];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	125051760	-	chr2	125052915	+	GTAGG	34	44	1314547_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTAGG;MAPQ=60;MATEID=1314547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_125048001_125073001_385C;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:67 DP:137 GQ:99 PL:[184.1, 0.0, 147.8] SR:44 DR:34 LR:-184.3 LO:184.3);ALT=[chr2:125052915[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	125766561	+	chr2	125768248	+	.	99	102	1317427_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1317427_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_125758501_125783501_64C;SPAN=1687;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:180 DP:139 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:102 DR:99 LR:-534.7 LO:534.7);ALT=C[chr2:125768248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	125768401	+	chr2	125766562	+	TCTATACTCACTACTACACTAT	0	83	1317429_1	99.0	.	EVDNC=ASSMB;INSERTION=TCTATACTCACTACTACACTAT;MAPQ=60;MATEID=1317429_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_125758501_125783501_113C;SPAN=1839;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:83 DP:146 GQ:99 PL:[234.5, 0.0, 119.0] SR:83 DR:0 LR:-236.4 LO:236.4);ALT=]chr2:125768401]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	125770948	+	chr8	118679719	-	.	11	6	5645811_1	37.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=5645811_2;MATENM=1;NM=6;NUMPARTS=2;SCTG=c_8_118678001_118703001_130C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:46 GQ:37.1 PL:[37.1, 0.0, 73.4] SR:6 DR:11 LR:-37.05 LO:37.75);ALT=A]chr8:118679719];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	125771009	-	chr8	118679601	+	ATTTTATTT	2	28	1317450_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTTTATTT;MAPQ=60;MATEID=1317450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_125758501_125783501_297C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:20 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:28 DR:2 LR:-85.82 LO:85.82);ALT=[chr8:118679601[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	126443251	+	chr2	126451832	+	.	192	44	1319794_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAAC;MAPQ=60;MATEID=1319794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_126420001_126445001_2C;SPAN=8581;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:210 DP:14 GQ:56.8 PL:[623.8, 56.8, 0.0] SR:44 DR:192 LR:-623.9 LO:623.9);ALT=C[chr2:126451832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117627975	+	chr17	46935421	+	.	20	0	9688610_1	50.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=9688610_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:117627975(+)-17:46935421(-)__17_46917501_46942501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:57 GQ:50.6 PL:[50.6, 0.0, 86.9] SR:0 DR:20 LR:-50.58 LO:51.13);ALT=T[chr17:46935421[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	118503476	-	chr8	118506369	+	.	10	0	5644804_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5644804_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:118503476(-)-8:118506369(-)__8_118482001_118507001D;SPAN=2893;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:124 GQ:0.3 PL:[0.0, 0.3, 300.3] SR:0 DR:10 LR:0.5846 LO:18.41);ALT=[chr8:118506369[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	46617220	+	chr17	46615632	+	.	29	79	9687001_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGA;MAPQ=60;MATEID=9687001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46599001_46624001_25C;SPAN=1588;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:105 DP:136 GQ:19.4 PL:[309.8, 0.0, 19.4] SR:79 DR:29 LR:-324.9 LO:324.9);ALT=]chr17:46617220]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	46615803	+	chr17	46617221	+	.	0	71	9687004_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AAG;MAPQ=60;MATEID=9687004_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46599001_46624001_26C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:71 DP:144 GQ:99 PL:[195.5, 0.0, 152.6] SR:71 DR:0 LR:-195.6 LO:195.6);ALT=G[chr17:46617221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47166552	+	chr17	47171633	+	CCCTC	132	119	9689820_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=CCCTC;MAPQ=60;MATEID=9689820_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_47162501_47187501_95C;SPAN=5081;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:226 DP:40 GQ:61 PL:[670.0, 61.0, 0.0] SR:119 DR:132 LR:-670.1 LO:670.1);ALT=T[chr17:47171633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
