chr12	60412349	+	chr12	60413509	+	.	25	41	5214151_1	99.0	.	DISC_MAPQ=25;EVDNC=ASDIS;HOMSEQ=GAAT;MAPQ=53;MATEID=5214151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_60392501_60417501_155C;SPAN=1160;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:42 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:41 DR:25 LR:-155.1 LO:155.1);ALT=T[chr12:60413509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	60521845	+	chr12	60525036	+	.	55	39	5214031_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGTCTA;MAPQ=60;MATEID=5214031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_60515001_60540001_183C;SPAN=3191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:45 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:39 DR:55 LR:-224.5 LO:224.5);ALT=A[chr12:60525036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
