chr8	78645247	+	chr8	78544926	+	TAAATCAGATA	41	13	5513473_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TAAATCAGATA;MAPQ=60;MATEID=5513473_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_78620501_78645501_359C;SPAN=100321;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:47 DP:33 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:13 DR:41 LR:-138.6 LO:138.6);ALT=]chr8:78645247]T;VARTYPE=BND:DUP-th;JOINTYPE=th
