chr9	66469907	-	chr9	66478641	+	.	53	0	4237978_1	87.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=4237978_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:66469907(-)-9:66478641(-)__9_66468501_66493501D;SPAN=8734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:325 GQ:87.1 PL:[87.1, 0.0, 701.0] SR:0 DR:53 LR:-86.9 LO:114.9);ALT=[chr9:66478641[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
