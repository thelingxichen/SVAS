chr8	132277700	+	chr8	132280534	+	.	60	0	5703985_1	99.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5703985_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:132277700(+)-8:132280534(-)__8_132275501_132300501D;SPAN=2834;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:23 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=T[chr8:132280534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
