chrX	34059778	+	chrX	34062705	+	ATTATAGTAT	5	15	7395907_1	42.0	.	DISC_MAPQ=24;EVDNC=ASDIS;INSERTION=ATTATAGTAT;MAPQ=24;MATEID=7395907_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_34055001_34080001_142C;SPAN=2927;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:9 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:15 DR:5 LR:-42.91 LO:42.91);ALT=C[chrX:34062705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
