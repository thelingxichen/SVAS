chr10	85522715	+	chr10	85523906	+	.	61	45	4646810_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4646810_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_10_85505001_85530001_292C;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:21 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:45 DR:61 LR:-250.9 LO:250.9);ALT=C[chr10:85523906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85899398	+	chr10	85903750	+	.	11	0	4647417_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4647417_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:85899398(+)-10:85903750(-)__10_85897001_85922001D;SPAN=4352;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=A[chr10:85903750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85899398	+	chr10	85901334	+	.	35	0	4647416_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4647416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:85899398(+)-10:85901334(-)__10_85897001_85922001D;SPAN=1936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:95 GQ:89.9 PL:[89.9, 0.0, 139.4] SR:0 DR:35 LR:-89.8 LO:90.41);ALT=A[chr10:85901334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85901386	+	chr10	85902410	+	.	0	47	4647419_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4647419_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ATAT;SCTG=c_10_85897001_85922001_74C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:78 GQ:54.8 PL:[134.0, 0.0, 54.8] SR:47 DR:0 LR:-135.8 LO:135.8);ALT=G[chr10:85902410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85901386	+	chr10	85903751	+	AATATGCCACCAAAACAAGAATTGGGATCCGGCGTGGGAGAACTGGCCAAGAACTCAAAGAGGCAGCATTGGAACCATCGATGGAAAAAATATTTAAAA	0	77	4647420_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AATATGCCACCAAAACAAGAATTGGGATCCGGCGTGGGAGAACTGGCCAAGAACTCAAAGAGGCAGCATTGGAACCATCGATGGAAAAAATATTTAAAA;MAPQ=60;MATEID=4647420_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_85897001_85922001_74C;SPAN=2365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:74 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:77 DR:0 LR:-227.8 LO:227.8);ALT=G[chr10:85903751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85902510	+	chr10	85903751	+	.	2	19	4647421_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4647421_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_10_85897001_85922001_74C;SPAN=1241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:64 GQ:52.1 PL:[52.1, 0.0, 101.6] SR:19 DR:2 LR:-51.98 LO:52.91);ALT=A[chr10:85903751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85908596	+	chr10	85909810	+	.	4	4	4647427_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4647427_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_85897001_85922001_180C;SPAN=1214;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:61 GQ:3.5 PL:[3.5, 0.0, 142.1] SR:4 DR:4 LR:-3.28 LO:11.59);ALT=T[chr10:85909810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	85910637	+	chr10	85912020	+	.	0	13	4647431_1	29.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4647431_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_85897001_85922001_73C;SPAN=1383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:51 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:13 DR:0 LR:-29.1 LO:31.04);ALT=G[chr10:85912020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
