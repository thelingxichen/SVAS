chr6	166733746	+	chr6	166738022	+	TGCATATGGGATGTACGACAGGCTA	0	22	3114572_1	47.0	.	EVDNC=ASSMB;INSERTION=TGCATATGGGATGTACGACAGGCTA;MAPQ=60;MATEID=3114572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_166722501_166747501_209C;SPAN=4276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:94 GQ:47.3 PL:[47.3, 0.0, 179.3] SR:22 DR:0 LR:-47.16 LO:51.57);ALT=T[chr6:166738022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166741847	+	chr6	166743648	+	GGCTAACGCAGCAAGATTGCCGAGGGTATAAAACACTGCAAAAAGCTTTATGCCGCCCGGAAGCCACAGCAATCCAGTTC	0	41	3114595_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGCTAACGCAGCAAGATTGCCGAGGGTATAAAACACTGCAAAAAGCTTTATGCCGCCCGGAAGCCACAGCAATCCAGTTC;MAPQ=60;MATEID=3114595_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_166722501_166747501_352C;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:77 GQ:71.6 PL:[114.5, 0.0, 71.6] SR:41 DR:0 LR:-115.0 LO:115.0);ALT=T[chr6:166743648[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166741847	+	chr6	166755905	+	GGCTAACGCAGCAAGATTGCCGAGGGTATAAAACACTGCAAAAAGCTTTATGCCGCCCGGAAGCCACAGCAATCCAGTTCCAAGAATAGAAAAGAAAACGCCACATACGAAGCAGATGGCAAACCATTTCAATCTGGTGTTGAAACTAAGGGATGAGGCATCCAGG	5	35	3114751_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=GGCTAACGCAGCAAGATTGCCGAGGGTATAAAACACTGCAAAAAGCTTTATGCCGCCCGGAAGCCACAGCAATCCAGTTCCAAGAATAGAAAAGAAAACGCCACATACGAAGCAGATGGCAAACCATTTCAATCTGGTGTTGAAACTAAGGGATGAGGCATCCAGG;MAPQ=60;MATEID=3114751_2;MATENM=2;NM=0;NUMPARTS=4;SCTG=c_6_166747001_166772001_327C;SPAN=14058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:35 DR:5 LR:-117.0 LO:117.0);ALT=T[chr6:166755905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166743125	+	chr6	166755955	+	.	16	0	3114753_1	36.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3114753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:166743125(+)-6:166755955(-)__6_166747001_166772001D;SPAN=12830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:0 DR:16 LR:-36.83 LO:38.71);ALT=T[chr6:166755955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166743737	+	chr6	166755905	+	.	28	15	3114601_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=3114601_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_6_166722501_166747501_332C;SPAN=12168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:28 GQ:9 PL:[99.0, 9.0, 0.0] SR:15 DR:28 LR:-99.02 LO:99.02);ALT=T[chr6:166755905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166779643	+	chr6	166796310	+	.	24	0	3114813_1	68.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3114813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:166779643(+)-6:166796310(-)__6_166796001_166821001D;SPAN=16667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:38 GQ:22.7 PL:[68.9, 0.0, 22.7] SR:0 DR:24 LR:-70.17 LO:70.17);ALT=A[chr6:166796310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	166780380	+	chr6	166796294	+	GTA	0	19	3114814_1	54.0	.	EVDNC=ASSMB;INSERTION=GTA;MAPQ=60;MATEID=3114814_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_166796001_166821001_182C;SPAN=15914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:30 GQ:18.2 PL:[54.5, 0.0, 18.2] SR:19 DR:0 LR:-55.59 LO:55.59);ALT=C[chr6:166796294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	167343281	+	chr6	167352383	+	GGCTTGGTGGAAGGCACTGGATTTTGGGTATCACTCCATATACTCTGGCAAGGGCATCTTTAAAATCTGCAACTTGGTAGTAATTGATGGATGGTTTTATCCCCAATTTTAGAAGCACA	3	70	3116257_1	99.0	.	DISC_MAPQ=51;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GGCTTGGTGGAAGGCACTGGATTTTGGGTATCACTCCATATACTCTGGCAAGGGCATCTTTAAAATCTGCAACTTGGTAGTAATTGATGGATGGTTTTATCCCCAATTTTAGAAGCACA;MAPQ=60;MATEID=3116257_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_167335001_167360001_258C;SPAN=9102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:113 GQ:68.6 PL:[203.9, 0.0, 68.6] SR:70 DR:3 LR:-207.3 LO:207.3);ALT=T[chr6:167352383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	167801544	+	chr6	167802735	+	.	7	21	3117542_1	68.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=TCCTGAGGTGTGTGAGGGTTGTGTGTGTGTCCTGAGGTGTGTGAGG;MAPQ=60;MATEID=3117542_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_167800501_167825501_141C;SPAN=1191;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:101 GQ:68.6 PL:[68.6, 0.0, 174.2] SR:21 DR:7 LR:-68.37 LO:71.02);ALT=G[chr6:167802735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
