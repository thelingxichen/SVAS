chr1	75772648	+	chr12	41847723	-	.	7	40	355154_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;MAPQ=21;MATEID=355154_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_75754001_75779001_34C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:72 GQ:36.8 PL:[135.8, 0.0, 36.8] SR:40 DR:7 LR:-138.6 LO:138.6);ALT=C]chr12:41847723];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	40881999	+	chr12	40883637	+	.	62	12	7559683_1	99.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=GTGACAGAGATAACTGGACTATCAGCTGGAGTGACAGGGACAA;MAPQ=0;MATEID=7559683_2;MATENM=2;NM=3;NUMPARTS=2;REPSEQ=AA;SCTG=c_12_40866001_40891001_69C;SECONDARY;SPAN=1638;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:34 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:12 DR:62 LR:-208.0 LO:208.0);ALT=A[chr12:40883637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
