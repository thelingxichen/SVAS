chr16	10837789	+	chr16	10840998	+	.	12	0	6107928_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6107928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:10837789(+)-16:10840998(-)__16_10829001_10854001D;SPAN=3209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:100 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:0 DR:12 LR:-12.52 LO:24.28);ALT=G[chr16:10840998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	10971240	+	chr16	10989137	+	.	0	8	6108708_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6108708_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_10951501_10976501_19C;SPAN=17897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.86 LO:17.27);ALT=G[chr16:10989137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11647545	+	chr16	11650367	+	.	4	62	6110802_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6110802_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_16_11637501_11662501_343C;SPAN=2822;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:121 GQ:99 PL:[175.4, 0.0, 116.0] SR:62 DR:4 LR:-175.8 LO:175.8);ALT=A[chr16:11650367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11647598	+	chr16	11680739	+	.	30	0	6111321_1	86.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6111321_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:11647598(+)-16:11680739(-)__16_11662001_11687001D;SPAN=33141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:48 GQ:29.9 PL:[86.0, 0.0, 29.9] SR:0 DR:30 LR:-87.48 LO:87.48);ALT=G[chr16:11680739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11650592	+	chr16	11680740	+	.	41	2	6111323_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6111323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_11662001_11687001_344C;SPAN=30148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:50 GQ:0.3 PL:[122.1, 0.3, 0.0] SR:2 DR:41 LR:-129.5 LO:129.5);ALT=C[chr16:11680740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11931972	+	chr16	11933552	+	.	18	2	6112037_1	53.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6112037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_11907001_11932001_12C;SPAN=1580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:48 GQ:53 PL:[53.0, 0.0, 62.9] SR:2 DR:18 LR:-53.02 LO:53.07);ALT=T[chr16:11933552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11935860	+	chr16	11940358	+	.	0	23	6112169_1	51.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6112169_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_11931501_11956501_28C;SPAN=4498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:92 GQ:51.2 PL:[51.2, 0.0, 170.0] SR:23 DR:0 LR:-51.0 LO:54.69);ALT=G[chr16:11940358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11941663	+	chr16	11945263	+	AATCTGACCCTCAGTTCTTTACTTGGAATTTTCCATAATACCACCATTAAAAATAAACTTTCATTCTCATTCAAAAGCAACCCATAATTGTTTTTCCTGGACTTGCAATGCGTCAAGAGAGCGTCCACTGCCTTTCTA	34	97	6112200_1	99.0	.	DISC_MAPQ=46;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=AATCTGACCCTCAGTTCTTTACTTGGAATTTTCCATAATACCACCATTAAAAATAAACTTTCATTCTCATTCAAAAGCAACCCATAATTGTTTTTCCTGGACTTGCAATGCGTCAAGAGAGCGTCCACTGCCTTTCTA;MAPQ=60;MATEID=6112200_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_11931501_11956501_414C;SPAN=3600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:100 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:97 DR:34 LR:-320.2 LO:320.2);ALT=C[chr16:11945263[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	11967029	+	chr16	11969612	+	.	4	4	6111845_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCTTACC;MAPQ=60;MATEID=6111845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_11956001_11981001_318C;SPAN=2583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:81 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:4 DR:4 LR:-1.162 LO:13.11);ALT=C[chr16:11969612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	12070694	+	chr16	12121173	+	.	9	0	6112576_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6112576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:12070694(+)-16:12121173(-)__16_12103001_12128001D;SPAN=50479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=C[chr16:12121173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	12875262	+	chr16	12897564	+	.	36	5	6115578_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6115578_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_12862501_12887501_303C;SPAN=22302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:5 DR:36 LR:-115.5 LO:115.5);ALT=T[chr16:12897564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
