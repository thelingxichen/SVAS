chr4	145316447	+	chr4	145319906	+	.	45	70	2970338_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=0;MATEID=2970338_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_145309501_145334501_385C;SECONDARY;SPAN=3459;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:40 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:70 DR:45 LR:-307.0 LO:307.0);ALT=C[chr4:145319906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
