chr8	21770023	+	chr8	21771050	+	.	36	11	3775883_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3775883_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_21756001_21781001_127C;SPAN=1027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:80 GQ:83.9 PL:[110.3, 0.0, 83.9] SR:11 DR:36 LR:-110.6 LO:110.6);ALT=T[chr8:21771050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
