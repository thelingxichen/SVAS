chr5	90499775	+	chr5	90502096	+	.	135	107	3603746_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTA;MAPQ=60;MATEID=3603746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_90478501_90503501_13C;SPAN=2321;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:192 DP:38 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:107 DR:135 LR:-567.7 LO:567.7);ALT=A[chr5:90502096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
