chr16	51958353	+	chr16	51935211	+	.	4	5	9315992_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATGTGA;MAPQ=60;MATEID=9315992_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_51940001_51965001_30C;SPAN=23142;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:5 DR:4 LR:-7.443 LO:16.0);ALT=]chr16:51958353]A;VARTYPE=BND:DUP-th;JOINTYPE=th
