chr15	99574554	+	chr15	99575609	+	.	124	20	9102394_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CACTGCAACCTCCGCCTCCCAGGTTCAAGTGATTCTCCTGCCTCAGCCTCCCGAGCAGCTGGGATTACAGGC;MAPQ=60;MATEID=9102394_2;MATENM=2;NM=5;NUMPARTS=2;SCTG=c_15_99568001_99593001_353C;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:141 DP:11 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:20 DR:124 LR:-415.9 LO:415.9);ALT=C[chr15:99575609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	100467009	+	chr15	100468647	+	.	8	0	9106361_1	9.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=9106361_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100467009(+)-15:100468647(-)__15_100450001_100475001D;SPAN=1638;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=G[chr15:100468647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
