chr4	186441637	+	chr4	186444074	+	.	0	93	3119757_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AA;MAPQ=60;MATEID=3119757_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_186420501_186445501_314C;SPAN=2437;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:32 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:93 DR:0 LR:-274.0 LO:274.0);ALT=A[chr4:186444074[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	187093524	+	chr4	187098241	+	.	13	0	3123011_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3123011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:187093524(+)-4:187098241(-)__4_187082001_187107001D;SPAN=4717;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:0 DR:13 LR:-22.32 LO:28.48);ALT=A[chr4:187098241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	187353484	+	chr4	187357165	+	.	65	36	3124824_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GCACACACGGCATTACCCAC;MAPQ=60;MATEID=3124824_2;MATENM=5;NM=3;NUMPARTS=2;SCTG=c_4_187351501_187376501_160C;SPAN=3681;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:97 DP:332 GQ:99 PL:[230.5, 0.0, 573.8] SR:36 DR:65 LR:-230.3 LO:238.4);ALT=C[chr4:187357165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
