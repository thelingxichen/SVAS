chr5	101992	+	chr5	100804	+	.	56	0	3138708_1	99.0	.	DISC_MAPQ=9;EVDNC=DSCRD;IMPRECISE;MAPQ=9;MATEID=3138708_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:100804(-)-5:101992(+)__5_98001_123001D;SPAN=1188;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:244 GQ:99 PL:[118.9, 0.0, 472.1] SR:0 DR:56 LR:-118.8 LO:130.7);ALT=]chr5:101992]T;VARTYPE=BND:DUP-th;JOINTYPE=th
