chr2	28518706	+	chr2	28488879	+	TCT	95	63	947023_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TCT;MAPQ=60;MATEID=947023_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_28518001_28543001_61C;SPAN=29827;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:132 DP:41 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:63 DR:95 LR:-389.5 LO:389.5);ALT=]chr2:28518706]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	28546933	+	chr2	28519797	+	.	86	49	947035_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=947035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_28518001_28543001_408C;SPAN=27136;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:112 DP:52 GQ:30 PL:[330.0, 30.0, 0.0] SR:49 DR:86 LR:-330.1 LO:330.1);ALT=]chr2:28546933]C;VARTYPE=BND:DUP-th;JOINTYPE=th
