chr11	50067304	-	chr11	50325635	+	ATGTCTAAAAGATGTCTAAAAGCCAGATA	79	30	4860799_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=ATGTCTAAAAGATGTCTAAAAGCCAGATA;MAPQ=60;MATEID=4860799_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_50323001_50348001_3C;SPAN=258331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:12 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:30 DR:79 LR:-293.8 LO:293.8);ALT=[chr11:50325635[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
