chr11	4968130	+	chr11	4976692	+	.	10	0	6629269_1	26.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6629269_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:4968130(+)-11:4976692(-)__11_4949001_4974001D;SPAN=8562;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:24 GQ:26.6 PL:[26.6, 0.0, 29.9] SR:0 DR:10 LR:-26.51 LO:26.53);ALT=C[chr11:4976692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
