chr2	236425722	+	chr2	236600479	+	.	0	51	1767242_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1767242_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_236596501_236621501_21C;SPAN=174757;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:51 DP:47 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:51 DR:0 LR:-148.5 LO:148.5);ALT=T[chr2:236600479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
