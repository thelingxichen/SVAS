chr18	5209639	+	chr18	5210659	+	ATATGTATACATATATACATAAATATAAATATATTTATAAAAAATATAAATATATTTAGCATGT	40	99	9873132_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATATGTATACATATATACATAAATATAAATATATTTATAAAAAATATAAATATATTTAGCATGT;MAPQ=60;MATEID=9873132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_5194001_5219001_192C;SPAN=1020;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:122 DP:35 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:99 DR:40 LR:-359.8 LO:359.8);ALT=T[chr18:5210659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
