chr2	122363756	+	chr2	122406948	+	.	7	3	971665_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=971665_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_122402001_122427001_315C;SPAN=43192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:36 GQ:23.3 PL:[23.3, 0.0, 62.9] SR:3 DR:7 LR:-23.26 LO:24.32);ALT=T[chr2:122406948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	122489781	+	chr2	122493189	+	.	0	23	972243_1	51.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=972243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_122475501_122500501_331C;SPAN=3408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:89 GQ:51.8 PL:[51.8, 0.0, 164.0] SR:23 DR:0 LR:-51.81 LO:55.07);ALT=C[chr2:122493189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	122513422	+	chr2	122514814	+	.	21	15	971966_1	57.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=971966_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_122500001_122525001_151C;SPAN=1392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:94 GQ:57.2 PL:[57.2, 0.0, 169.4] SR:15 DR:21 LR:-57.06 LO:60.23);ALT=G[chr2:122514814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	122513439	+	chr2	122516285	+	.	8	0	971967_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=971967_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:122513439(+)-2:122516285(-)__2_122500001_122525001D;SPAN=2846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=C[chr2:122516285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	122516382	+	chr2	122518982	+	.	0	7	971981_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=971981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_122500001_122525001_326C;SPAN=2600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:7 DR:0 LR:-3.059 LO:13.4);ALT=G[chr2:122518982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
