chr4	165861260	-	chr4	165869118	+	.	8	0	2315930_1	12.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2315930_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:165861260(-)-4:165869118(-)__4_165840501_165865501D;SPAN=7858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=[chr4:165869118[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	166024268	+	chr4	166033921	+	.	8	0	2316574_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2316574_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:166024268(+)-4:166033921(-)__4_166012001_166037001D;SPAN=9653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:0 DR:8 LR:5.561 LO:14.1);ALT=G[chr4:166033921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
