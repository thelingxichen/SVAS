chr7	91402536	-	chr7	91404185	+	.	9	0	3451375_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3451375_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:91402536(-)-7:91404185(-)__7_91385001_91410001D;SPAN=1649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:0 DR:9 LR:-1.533 LO:16.86);ALT=[chr7:91404185[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	91570461	+	chr7	91603023	+	.	0	7	3452018_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=3452018_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_91556501_91581501_310C;SPAN=32562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:64 GQ:5.9 PL:[5.9, 0.0, 147.8] SR:7 DR:0 LR:-5.768 LO:13.86);ALT=G[chr7:91603023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	92463006	+	chr7	92465789	+	.	60	3	3455068_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=3455068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_92438501_92463501_345C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:53 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:3 DR:60 LR:-178.2 LO:178.2);ALT=T[chr7:92465789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112178163	+	chr7	92976835	+	.	28	25	4689873_1	99.0	.	DISC_MAPQ=4;EVDNC=ASDIS;MAPQ=60;MATEID=4689873_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_10_112161001_112186001_206C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:33 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:25 DR:28 LR:-135.3 LO:135.3);ALT=]chr10:112178163]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	93416941	+	chr7	93422992	+	.	62	30	3458153_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAATCATCATTCTT;MAPQ=60;MATEID=3458153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_93418501_93443501_141C;SPAN=6051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:27 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:30 DR:62 LR:-214.6 LO:214.6);ALT=T[chr7:93422992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	93628652	+	chr7	93633594	+	.	8	0	3458589_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3458589_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:93628652(+)-7:93633594(-)__7_93614501_93639501D;SPAN=4942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:0 DR:8 LR:2.581 LO:14.46);ALT=T[chr7:93633594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	111572124	+	chr10	111578217	+	.	29	16	4689216_1	18.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TAAAGCCATGTTCT;MAPQ=60;MATEID=4689216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_111548501_111573501_0C;SPAN=6093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:443 GQ:18.9 PL:[18.9, 0.0, 1055.0] SR:16 DR:29 LR:-18.62 LO:80.42);ALT=T[chr10:111578217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	111651585	+	chr10	111667449	+	CGCAGAGCCATCGAATCCAGAGACAAAAGCCCGCCGACAGTCACATGGAGCAATATACTCACT	0	18	4688894_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CGCAGAGCCATCGAATCCAGAGACAAAAGCCCGCCGACAGTCACATGGAGCAATATACTCACT;MAPQ=60;MATEID=4688894_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_111646501_111671501_257C;SPAN=15864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:61 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:18 DR:0 LR:-42.89 LO:44.34);ALT=C[chr10:111667449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	111667576	+	chr10	111674769	+	.	2	12	4688921_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4688921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_111646501_111671501_291C;SPAN=7193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:31 GQ:34.7 PL:[38.0, 0.0, 34.7] SR:12 DR:2 LR:-37.82 LO:37.82);ALT=G[chr10:111674769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	111667627	+	chr10	111683155	+	.	29	0	4688922_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4688922_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:111667627(+)-10:111683155(-)__10_111646501_111671501D;SPAN=15528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:25 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=G[chr10:111683155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112058548	+	chr10	112063225	+	.	3	8	4689396_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4689396_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_112063001_112088001_165C;SPAN=4677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:26 GQ:26 PL:[26.0, 0.0, 35.9] SR:8 DR:3 LR:-25.97 LO:26.07);ALT=C[chr10:112063225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112058567	+	chr10	112064508	+	.	8	0	4689397_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4689397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:112058567(+)-10:112064508(-)__10_112063001_112088001D;SPAN=5941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:21 GQ:20.9 PL:[20.9, 0.0, 27.5] SR:0 DR:8 LR:-20.72 LO:20.82);ALT=A[chr10:112064508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112063347	+	chr10	112064506	+	.	0	16	4689398_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4689398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_112063001_112088001_87C;SPAN=1159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:60 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:16 DR:0 LR:-36.56 LO:38.57);ALT=T[chr10:112064506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112327590	+	chr10	112328693	+	.	10	0	4689940_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4689940_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:112327590(+)-10:112328693(-)__10_112308001_112333001D;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:43 GQ:21.5 PL:[21.5, 0.0, 80.9] SR:0 DR:10 LR:-21.36 LO:23.41);ALT=G[chr10:112328693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112328771	+	chr10	112337179	+	TGGGCAGAAATGGATCTGGAAAAAGTAACTTTTTTTATGCAATTCAGTTTGTTCTCAGTGATGAGTTTAGTCATCTTCGTCCAGAACAGCGGTTGGCTTTATTGCAT	0	16	4689946_1	45.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TGGGCAGAAATGGATCTGGAAAAAGTAACTTTTTTTATGCAATTCAGTTTGTTCTCAGTGATGAGTTTAGTCATCTTCGTCCAGAACAGCGGTTGGCTTTATTGCAT;MAPQ=60;MATEID=4689946_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_112308001_112333001_228C;SPAN=8408;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:27 GQ:19.1 PL:[45.5, 0.0, 19.1] SR:16 DR:0 LR:-46.04 LO:46.04);ALT=G[chr10:112337179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112631770	+	chr10	112635722	+	.	9	0	4690474_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4690474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:112631770(+)-10:112635722(-)__10_112626501_112651501D;SPAN=3952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:59 GQ:13.7 PL:[13.7, 0.0, 129.2] SR:0 DR:9 LR:-13.72 LO:19.22);ALT=C[chr10:112635722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112631811	+	chr10	112640989	+	.	10	0	4690475_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4690475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:112631811(+)-10:112640989(-)__10_112626501_112651501D;SPAN=9178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:0 DR:10 LR:-17.57 LO:22.03);ALT=A[chr10:112640989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112655846	+	chr10	112657784	+	.	3	4	4690551_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4690551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_112651001_112676001_290C;SPAN=1938;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:48 GQ:0.2 PL:[0.2, 0.0, 115.7] SR:4 DR:3 LR:-0.1996 LO:7.424);ALT=G[chr10:112657784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	112679468	+	chr10	112723879	+	.	43	0	4690626_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4690626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:112679468(+)-10:112723879(-)__10_112700001_112725001D;SPAN=44411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:20 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=T[chr10:112723879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
