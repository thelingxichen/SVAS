chr12	46264007	+	chr12	46372954	-	G	66	32	7581208_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=7581208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_46256001_46281001_453C;SPAN=108947;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:96 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:32 DR:66 LR:-283.9 LO:283.9);ALT=C]chr12:46372954];VARTYPE=BND:INV-hh;JOINTYPE=hh
