chr1	158867533	+	chr1	158869982	+	.	75	94	578116_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAT;MAPQ=60;MATEID=578116_2;MATENM=10;NM=0;NUMPARTS=2;SCTG=c_1_158858001_158883001_64C;SPAN=2449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:142 DP:37 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:94 DR:75 LR:-419.2 LO:419.2);ALT=T[chr1:158869982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	158867581	+	chr1	158870245	+	.	18	0	578122_1	49.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=578122_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:158867581(+)-1:158870245(-)__1_158858001_158883001D;SPAN=2664;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:36 GQ:36.5 PL:[49.7, 0.0, 36.5] SR:0 DR:18 LR:-49.75 LO:49.75);ALT=T[chr1:158870245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159013730	+	chr1	159018118	+	.	8	0	577623_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=577623_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159013730(+)-1:159018118(-)__1_159005001_159030001D;SPAN=4388;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:114 GQ:4.2 PL:[0.0, 4.2, 283.8] SR:0 DR:8 LR:4.477 LO:14.23);ALT=C[chr1:159018118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159428669	+	chr1	159494967	-	.	11	0	579694_1	16.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=579694_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159428669(+)-1:159494967(+)__1_159470501_159495501D;SPAN=66298;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:0 DR:11 LR:-16.53 LO:23.43);ALT=G]chr1:159494967];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	159738428	+	chr1	224528411	+	.	12	0	581422_1	16.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=581422_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159738428(+)-1:224528411(-)__1_159715501_159740501D;SPAN=64789983;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:0 DR:12 LR:-16.31 LO:25.12);ALT=C[chr1:224528411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	223974373	-	chr1	223975409	+	.	9	0	838951_1	9.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=838951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:223974373(-)-1:223975409(-)__1_223954501_223979501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=[chr1:223975409[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	224815674	+	chr1	224818308	+	.	62	62	841330_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=841330_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_224812001_224837001_81C;SPAN=2634;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:24 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:62 DR:62 LR:-307.0 LO:307.0);ALT=G[chr1:224818308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	225248324	+	chr1	225133358	+	.	15	0	842237_1	46.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=842237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:225133358(-)-1:225248324(+)__1_225228501_225253501D;SPAN=114966;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:16 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:0 DR:15 LR:-46.21 LO:46.21);ALT=]chr1:225248324]A;VARTYPE=BND:DUP-th;JOINTYPE=th
