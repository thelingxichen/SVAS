chr12	57001806	-	chr12	57002862	+	.	10	0	7632902_1	0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=7632902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57001806(-)-12:57002862(-)__12_56987001_57012001D;SPAN=1056;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:133 GQ:2.7 PL:[0.0, 2.7, 326.7] SR:0 DR:10 LR:3.023 LO:18.09);ALT=[chr12:57002862[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
