chr11	117005284	+	chr11	117080764	-	.	78	0	5017516_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5017516_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:117005284(+)-11:117080764(+)__11_117061001_117086001D;SPAN=75480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:46 GQ:21 PL:[231.0, 21.0, 0.0] SR:0 DR:78 LR:-231.1 LO:231.1);ALT=C]chr11:117080764];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	117105095	+	chr11	117109315	+	.	3	6	5017446_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5017446_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_117085501_117110501_47C;SPAN=4220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:6 DR:3 LR:-9.39 LO:18.21);ALT=G[chr11:117109315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	117109827	+	chr11	117115160	+	ACTGACTTTAAGACAGCTGATTCAGAGGTAAACACAGATCAAGATATTGAAAAGAATTT	0	9	5018098_1	18.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ACTGACTTTAAGACAGCTGATTCAGAGGTAAACACAGATCAAGATATTGAAAAGAATTT;MAPQ=60;MATEID=5018098_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_117110001_117135001_352C;SPAN=5333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:9 DR:0 LR:-18.87 LO:20.92);ALT=G[chr11:117115160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	117209384	+	chr11	117214880	+	.	0	14	5017743_1	26.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5017743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_117208001_117233001_358C;SPAN=5496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:14 DR:0 LR:-26.17 LO:31.35);ALT=G[chr11:117214880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	117214993	+	chr11	117222505	+	.	0	10	5017756_1	6.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5017756_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_117208001_117233001_80C;SPAN=7512;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:99 GQ:6.2 PL:[6.2, 0.0, 233.9] SR:10 DR:0 LR:-6.189 LO:19.44);ALT=G[chr11:117222505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	117920353	+	chr15	57019272	-	.	9	0	5958719_1	21.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=5958719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:117920353(+)-15:57019272(+)__15_57011501_57036501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:29 GQ:21.8 PL:[21.8, 0.0, 48.2] SR:0 DR:9 LR:-21.85 LO:22.41);ALT=C]chr15:57019272];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	118065133	+	chr11	118067450	+	.	5	7	5020061_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5020061_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_118041001_118066001_27C;SPAN=2317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:7 DR:5 LR:-23.85 LO:25.91);ALT=C[chr11:118067450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118067538	+	chr11	118068713	+	.	2	3	5019934_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5019934_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_11_118065501_118090501_272C;SPAN=1175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:98 GQ:9.9 PL:[0.0, 9.9, 257.4] SR:3 DR:2 LR:10.05 LO:8.181);ALT=T[chr11:118068713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118081429	+	chr11	118083121	+	.	2	25	5019968_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5019968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_118065501_118090501_310C;SPAN=1692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:110 GQ:59.3 PL:[59.3, 0.0, 207.8] SR:25 DR:2 LR:-59.33 LO:63.94);ALT=T[chr11:118083121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118081474	+	chr11	118095666	+	.	16	0	5020186_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5020186_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118081474(+)-11:118095666(-)__11_118090001_118115001D;SPAN=14192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.0 LO:39.93);ALT=C[chr11:118095666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118083277	+	chr11	118095656	+	CAGTAACACTGGCAGCAGGATGAGTTTCAGTGGGCAAAACATGCTGCTCTCAACTTTCAAAT	50	24	5020188_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CAGTAACACTGGCAGCAGGATGAGTTTCAGTGGGCAAAACATGCTGCTCTCAACTTTCAAAT;MAPQ=60;MATEID=5020188_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_118090001_118115001_112C;SPAN=12379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:40 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:24 DR:50 LR:-188.1 LO:188.1);ALT=C[chr11:118095656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118085602	+	chr11	118095656	+	.	10	8	5020189_1	32.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5020189_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_11_118090001_118115001_112C;SPAN=10054;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:40 GQ:32 PL:[32.0, 0.0, 65.0] SR:8 DR:10 LR:-32.08 LO:32.69);ALT=C[chr11:118095656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118230432	+	chr11	118239344	+	.	9	0	5020506_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5020506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118230432(+)-11:118239344(-)__11_118237001_118262001D;SPAN=8912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=G[chr11:118239344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118230432	+	chr11	118235753	+	.	12	0	5020468_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5020468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118230432(+)-11:118235753(-)__11_118212501_118237501D;SPAN=5321;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:93 GQ:14.6 PL:[14.6, 0.0, 209.3] SR:0 DR:12 LR:-14.42 LO:24.68);ALT=G[chr11:118235753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118235916	+	chr11	118239345	+	.	0	9	5020507_1	16.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5020507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_118237001_118262001_13C;SPAN=3429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:9 DR:0 LR:-16.43 LO:20.02);ALT=G[chr11:118239345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118272432	+	chr11	118277651	+	.	91	19	5020821_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5020821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_118261501_118286501_322C;SPAN=5219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:140 GQ:47.9 PL:[292.1, 0.0, 47.9] SR:19 DR:91 LR:-302.2 LO:302.2);ALT=G[chr11:118277651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118272452	+	chr11	118279712	+	.	17	0	5020823_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5020823_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118272452(+)-11:118279712(-)__11_118261501_118286501D;SPAN=7260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:122 GQ:23.3 PL:[23.3, 0.0, 270.8] SR:0 DR:17 LR:-23.06 LO:35.58);ALT=G[chr11:118279712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118443267	+	chr11	118451960	+	.	5	2	5021230_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5021230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_118433001_118458001_94C;SPAN=8693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:97 GQ:6.3 PL:[0.0, 6.3, 247.5] SR:2 DR:5 LR:6.474 LO:10.33);ALT=T[chr11:118451960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	118657233	+	chr11	118661804	+	.	24	0	5022320_1	56.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5022320_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:118657233(+)-11:118661804(-)__11_118653501_118678501D;SPAN=4571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:86 GQ:56 PL:[56.0, 0.0, 151.7] SR:0 DR:24 LR:-55.92 LO:58.42);ALT=A[chr11:118661804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	119077325	+	chr11	119103156	+	.	0	10	5023762_1	22.0	.	EVDNC=ASSMB;HOMSEQ=AGGTG;MAPQ=60;MATEID=5023762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_119070001_119095001_287C;SPAN=25831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:41 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:10 DR:0 LR:-21.9 LO:23.65);ALT=G[chr11:119103156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	56996465	+	chr15	56999276	+	.	0	12	5958721_1	33.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=TTAC;MAPQ=60;MATEID=5958721_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_15_57011501_57036501_20C;SPAN=2811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:0 GQ:3 PL:[33.0, 3.0, 0.0] SR:12 DR:0 LR:-33.01 LO:33.01);ALT=C[chr15:56999276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	56996511	+	chr15	57025651	+	.	19	0	5958722_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5958722_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:56996511(+)-15:57025651(-)__15_57011501_57036501D;SPAN=29140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:31 GQ:18.2 PL:[54.5, 0.0, 18.2] SR:0 DR:19 LR:-55.13 LO:55.13);ALT=A[chr15:57025651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
