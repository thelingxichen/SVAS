chrX	64949586	+	chr5	25910065	+	.	8	0	7437146_1	19.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7437146_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:25910065(-)-23:64949586(+)__23_64925001_64950001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:0 DR:8 LR:-19.36 LO:19.88);ALT=]chrX:64949586]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chrX	64947773	+	chrX	64949298	+	.	0	8	7437175_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=7437175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_64925001_64950001_285C;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:8 DR:0 LR:-12.05 LO:17.05);ALT=T[chrX:64949298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	64953143	+	chrX	64955128	+	.	4	8	7437285_1	17.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7437285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_64949501_64974501_245C;SPAN=1985;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:8 DR:4 LR:-17.89 LO:23.8);ALT=G[chrX:64955128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	65235393	+	chrX	65236904	+	.	6	4	7437518_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7437518_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_65219001_65244001_277C;SPAN=1511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:59 GQ:7.1 PL:[7.1, 0.0, 135.8] SR:4 DR:6 LR:-7.123 LO:14.13);ALT=G[chrX:65236904[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	65235394	+	chrX	65238664	+	.	17	2	7437519_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7437519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_65219001_65244001_92C;SPAN=3270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:63 GQ:42.5 PL:[42.5, 0.0, 108.5] SR:2 DR:17 LR:-42.35 LO:44.03);ALT=G[chrX:65238664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	65235427	+	chrX	65239964	+	.	8	0	7437520_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7437520_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:65235427(+)-23:65239964(-)__23_65219001_65244001D;SPAN=4537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:0 DR:8 LR:-8.798 LO:16.28);ALT=C[chrX:65239964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
