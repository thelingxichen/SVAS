chr2	52749686	+	chr2	52785271	+	ATTTA	0	87	998883_1	99.0	.	EVDNC=ASSMB;INSERTION=ATTTA;MAPQ=60;MATEID=998883_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_52748501_52773501_41C;SPAN=35585;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:18 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:87 DR:0 LR:-257.5 LO:257.5);ALT=A[chr2:52785271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	53625772	+	chr2	53628000	+	.	74	71	1002814_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAATTATAT;MAPQ=60;MATEID=1002814_2;MATENM=1;NM=6;NUMPARTS=2;SCTG=c_2_53606001_53631001_145C;SPAN=2228;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:119 DP:40 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:71 DR:74 LR:-353.2 LO:353.2);ALT=T[chr2:53628000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	54111588	+	chr14	40317397	-	.	15	34	1004336_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;HOMSEQ=GGATCACAAGGTCAAGAGATTGAGACCATCCTGGCCAACATG;MAPQ=49;MATEID=1004336_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_2_54096001_54121001_230C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:97 GQ:99 PL:[135.5, 0.0, 99.2] SR:34 DR:15 LR:-135.8 LO:135.8);ALT=C]chr14:40317397];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	54565493	+	chr2	54567474	+	TAA	0	105	1006357_1	99.0	.	EVDNC=ASSMB;INSERTION=TAA;MAPQ=60;MATEID=1006357_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_54561501_54586501_307C;SPAN=1981;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:42 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:105 DR:0 LR:-310.3 LO:310.3);ALT=G[chr2:54567474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	39987479	+	chr14	39992269	+	.	14	0	8455636_1	13.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=8455636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:39987479(+)-14:39992269(-)__14_39984001_40009001D;SPAN=4790;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:120 GQ:13.7 PL:[13.7, 0.0, 277.7] SR:0 DR:14 LR:-13.7 LO:28.14);ALT=T[chr14:39992269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
