chr13	104703629	+	chr13	104705265	-	.	9	0	8294449_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=8294449_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:104703629(+)-13:104705265(+)__13_104688501_104713501D;SPAN=1636;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:148 GQ:10.3 PL:[0.0, 10.3, 379.5] SR:0 DR:9 LR:10.39 LO:15.43);ALT=G]chr13:104705265];VARTYPE=BND:INV-hh;JOINTYPE=hh
