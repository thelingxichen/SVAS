chr3	143150495	+	chr3	143151628	+	.	56	33	2376151_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CCCGGCTAATTTTT;MAPQ=60;MATEID=2376151_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_143129001_143154001_226C;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:68 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:33 DR:56 LR:-241.0 LO:241.0);ALT=T[chr3:143151628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
