chr12	93258765	+	chr12	93322819	+	CTGAAGAGCTTTCATTATTGACGTCCACTGTGTTTATAGGAGTTGCTGATGAATCTAAATCAGAACCTTGAGAGCCAACTCTCCCAGGAGT	4	14	5289712_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTGAAGAGCTTTCATTATTGACGTCCACTGTGTTTATAGGAGTTGCTGATGAATCTAAATCAGAACCTTGAGAGCCAACTCTCCCAGGAGT;MAPQ=60;MATEID=5289712_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_93320501_93345501_9C;SPAN=64054;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:28 GQ:22.1 PL:[45.2, 0.0, 22.1] SR:14 DR:4 LR:-45.63 LO:45.63);ALT=T[chr12:93322819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93805090	+	chr12	93835623	+	.	64	0	5291480_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5291480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:93805090(+)-12:93835623(-)__12_93835001_93860001D;SPAN=30533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:28 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=C[chr12:93835623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93861376	+	chr12	93870729	+	.	23	0	5291576_1	53.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5291576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:93861376(+)-12:93870729(-)__12_93859501_93884501D;SPAN=9353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:84 GQ:53.3 PL:[53.3, 0.0, 149.0] SR:0 DR:23 LR:-53.17 LO:55.76);ALT=T[chr12:93870729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93861376	+	chr12	93863001	+	.	13	0	5291575_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5291575_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:93861376(+)-12:93863001(-)__12_93859501_93884501D;SPAN=1625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:81 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:0 DR:13 LR:-20.97 LO:28.08);ALT=T[chr12:93863001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93863131	+	chr12	93873163	+	ATGGAGCTTTATATTGTGTTTGTCATAAATCTACGTATTCTCCTCTACCAGATGACTATAATT	0	44	5291581_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGGAGCTTTATATTGTGTTTGTCATAAATCTACGTATTCTCCTCTACCAGATGACTATAATT;MAPQ=60;MATEID=5291581_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_93859501_93884501_218C;SPAN=10032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:72 GQ:46.7 PL:[125.9, 0.0, 46.7] SR:44 DR:0 LR:-127.6 LO:127.6);ALT=A[chr12:93873163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	93964993	+	chr12	93966459	+	.	0	12	5291750_1	23.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5291750_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_93957501_93982501_314C;SPAN=1466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:12 DR:0 LR:-23.36 LO:27.2);ALT=G[chr12:93966459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	94071249	+	chr12	94072545	+	.	6	4	5292107_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5292107_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_94055501_94080501_82C;SPAN=1296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:4 DR:6 LR:0.4634 LO:12.88);ALT=G[chr12:94072545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
