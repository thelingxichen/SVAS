chr18	59046408	+	chr18	59144128	+	.	4	7	10037488_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=10037488_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_59143001_59168001_213C;SPAN=97720;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:7 DR:4 LR:-22.12 LO:22.58);ALT=A[chr18:59144128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
