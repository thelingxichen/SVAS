chr7	11875806	+	chr7	11878592	+	.	121	82	4545587_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=4545587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_11858001_11883001_292C;SPAN=2786;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:160 DP:91 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:82 DR:121 LR:-475.3 LO:475.3);ALT=A[chr7:11878592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
