chr1	4125146	+	chr1	4126426	+	.	0	4	23386_1	0	.	EVDNC=ASSMB;HOMSEQ=CACACAC;MAPQ=60;MATEID=23386_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_4116001_4141001_195C;SPAN=1280;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:122 GQ:19.5 PL:[0.0, 19.5, 333.3] SR:4 DR:0 LR:19.85 LO:5.767);ALT=C[chr1:4126426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	4138728	+	chr1	4137605	+	.	58	0	23441_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=23441_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:4137605(-)-1:4138728(+)__1_4116001_4141001D;SPAN=1123;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:255 GQ:99 PL:[122.5, 0.0, 495.5] SR:0 DR:58 LR:-122.4 LO:135.1);ALT=]chr1:4138728]C;VARTYPE=BND:DUP-th;JOINTYPE=th
