chr4	138687340	+	chr4	138688934	+	TT	0	10	2943845_1	0	.	EVDNC=ASSMB;INSERTION=TT;MAPQ=60;MATEID=2943845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_138670001_138695001_317C;SPAN=1594;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:162 GQ:10.6 PL:[0.0, 10.6, 412.6] SR:10 DR:0 LR:10.88 LO:17.21);ALT=T[chr4:138688934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	138966211	+	chr4	138967219	+	T	0	102	2944974_1	99.0	.	EVDNC=ASSMB;INSERTION=T;MAPQ=60;MATEID=2944974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_138964001_138989001_179C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:37 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:102 DR:0 LR:-300.4 LO:300.4);ALT=G[chr4:138967219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	139388970	-	chr4	139390014	+	.	11	0	2946288_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2946288_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:139388970(-)-4:139390014(-)__4_139380501_139405501D;SPAN=1044;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:132 GQ:0.8 PL:[0.8, 0.0, 317.6] SR:0 DR:11 LR:-0.549 LO:20.42);ALT=[chr4:139390014[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	139468878	+	chr4	139473240	+	.	96	86	2947096_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=AGAGTGAACAGGCAACC;MAPQ=55;MATEID=2947096_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=CC;SCTG=c_4_139454001_139479001_114C;SECONDARY;SPAN=4362;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:175 DP:84 GQ:47.2 PL:[518.2, 47.2, 0.0] SR:86 DR:96 LR:-518.2 LO:518.2);ALT=C[chr4:139473240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
