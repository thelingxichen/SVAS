chr11	13023198	+	chr18	53590863	-	.	28	39	10026880_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CATTAGATTCTCATAAGGAGCATGCAGCCTAG;MAPQ=60;MATEID=10026880_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_18_53581501_53606501_252C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:47 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:39 DR:28 LR:-184.8 LO:184.8);ALT=G]chr18:53590863];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	13565922	+	chr20	37970249	+	.	6	28	6646058_1	89.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CCTGCCTCAGCCTCCCAAGTAGATGG;MAPQ=60;MATEID=6646058_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_13548501_13573501_86C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:30 DP:8 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:28 DR:6 LR:-89.12 LO:89.12);ALT=G[chr20:37970249[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	37970324	+	chr11	13566291	+	.	6	27	10528954_1	74.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCCACCATGCCTGGCTAATTTTTGTATTTTTAGTAG;MAPQ=60;MATEID=10528954_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_37950501_37975501_94C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:92 GQ:74.3 PL:[74.3, 0.0, 146.9] SR:27 DR:6 LR:-74.11 LO:75.49);ALT=]chr20:37970324]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	13681970	+	chr11	13683767	+	.	69	52	6646192_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=6646192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_13671001_13696001_75C;SPAN=1797;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:20 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:52 DR:69 LR:-316.9 LO:316.9);ALT=T[chr11:13683767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	53560582	+	chr18	70639656	+	.	53	0	10065661_1	99.0	.	DISC_MAPQ=6;EVDNC=DSCRD;IMPRECISE;MAPQ=6;MATEID=10065661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:53560582(+)-18:70639656(-)__18_70633501_70658501D;SPAN=17079074;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:49 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:0 DR:53 LR:-155.1 LO:155.1);ALT=A[chr18:70639656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
