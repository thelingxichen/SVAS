chr1	179263071	+	chr1	179271810	+	.	5	6	424672_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=424672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_179266501_179291501_194C;SPAN=8739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:52 GQ:9.2 PL:[9.2, 0.0, 114.8] SR:6 DR:5 LR:-9.019 LO:14.54);ALT=G[chr1:179271810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	180047809	+	chr1	180049652	+	.	3	3	427517_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=427517_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_180026001_180051001_125C;SPAN=1843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:99 GQ:10.2 PL:[0.0, 10.2, 260.7] SR:3 DR:3 LR:10.32 LO:8.158);ALT=T[chr1:180049652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
