chr4	37651123	+	chr4	37687822	+	.	15	10	1941717_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1941717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_37681001_37706001_234C;SPAN=36699;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:43 GQ:47.9 PL:[47.9, 0.0, 54.5] SR:10 DR:15 LR:-47.77 LO:47.81);ALT=C[chr4:37687822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	37828426	+	chr4	37831583	+	.	9	0	1941921_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1941921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:37828426(+)-4:37831583(-)__4_37828001_37853001D;SPAN=3157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=C[chr4:37831583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	37831754	+	chr4	37836238	+	.	0	7	1941928_1	8.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1941928_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_37828001_37853001_270C;SPAN=4484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:54 GQ:8.6 PL:[8.6, 0.0, 120.8] SR:7 DR:0 LR:-8.477 LO:14.41);ALT=G[chr4:37836238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	37892971	+	chr4	37903621	+	.	8	5	1942068_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=1942068_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_37901501_37926501_136C;SPAN=10650;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:5 DR:8 LR:-22.39 LO:22.75);ALT=T[chr4:37903621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
