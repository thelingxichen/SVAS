chr1	72766324	+	chr1	72811840	+	.	110	97	344172_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=344172_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_72789501_72814501_3C;SPAN=45516;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:170 DP:19 GQ:46 PL:[505.0, 46.0, 0.0] SR:97 DR:110 LR:-505.0 LO:505.0);ALT=G[chr1:72811840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	73757095	+	chr11	38903326	+	.	8	0	6754690_1	13.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6754690_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:73757095(+)-11:38903326(-)__11_38881501_38906501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=C[chr11:38903326[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	51265173	+	chr8	51409780	+	.	58	54	5466830_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=5466830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_51401001_51426001_6C;SPAN=144607;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:10 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:54 DR:58 LR:-267.4 LO:267.4);ALT=A[chr8:51409780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	52051329	-	chr11	68196393	+	.	4	19	6884949_1	52.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=6884949_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_11_68183501_68208501_285C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:74 GQ:52.7 PL:[52.7, 0.0, 125.3] SR:19 DR:4 LR:-52.57 LO:54.28);ALT=[chr11:68196393[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	52731482	+	chr11	38812658	+	.	36	23	5468960_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=ATAA;MAPQ=60;MATEID=5468960_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_52724001_52749001_227C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:39 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:23 DR:36 LR:-148.5 LO:148.5);ALT=A[chr11:38812658[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	38760453	+	chr11	38761728	-	.	11	0	6753835_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6753835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:38760453(+)-11:38761728(+)__11_38759001_38784001D;SPAN=1275;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:99 GQ:9.5 PL:[9.5, 0.0, 230.6] SR:0 DR:11 LR:-9.49 LO:21.86);ALT=T]chr11:38761728];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	67868407	-	chr11	67869498	+	.	8	0	6879044_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6879044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67868407(-)-11:67869498(-)__11_67865001_67890001D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:203 GQ:28.3 PL:[0.0, 28.3, 547.9] SR:0 DR:8 LR:28.59 LO:12.18);ALT=[chr11:67869498[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	68201970	-	chr16	12002671	+	.	8	0	9151795_1	15.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=9151795_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68201970(-)-16:12002671(-)__16_11980501_12005501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=[chr16:12002671[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
