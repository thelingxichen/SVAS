chr6	32778708	+	chr6	32779821	+	ACGCCACCACGCAAGGCTAATTTTTTGTGTTTTTAGTAGAGACGGGG	100	182	4120868_1	99.0	.	DISC_MAPQ=38;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=ACGCCACCACGCAAGGCTAATTTTTTGTGTTTTTAGTAGAGACGGGG;MAPQ=60;MATEID=4120868_2;MATENM=1;NM=10;NUMPARTS=3;SCTG=c_6_32756501_32781501_14C;SPAN=1113;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:261 DP:31 GQ:70.3 PL:[772.3, 70.3, 0.0] SR:182 DR:100 LR:-772.4 LO:772.4);ALT=C[chr6:32779821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32853410	+	chr6	32779821	+	.	38	122	4121402_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=4121402_2;MATENM=2;NM=1;NUMPARTS=3;REPSEQ=GGGG;SCTG=c_6_32830001_32855001_294C;SPAN=73589;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:68 GQ:36 PL:[396.0, 36.0, 0.0] SR:122 DR:38 LR:-396.1 LO:396.1);ALT=]chr6:32853410]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32868228	+	chr6	32883493	-	.	2	3	4121815_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGGTAA;MAPQ=60;MATEID=4121815_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32879001_32904001_316C;SPAN=15265;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:5 DP:52 GQ:2.6 PL:[2.6, 0.0, 121.4] SR:3 DR:2 LR:-2.417 LO:9.606);ALT=C]chr6:32883493];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	33026738	+	chr6	33028600	+	.	43	0	4123553_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4123553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:33026738(+)-6:33028600(-)__6_33026001_33051001D;SPAN=1862;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:11 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=T[chr6:33028600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
