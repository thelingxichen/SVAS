chr8	95835789	+	chr8	95837120	+	.	0	5	3978117_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3978117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_95819501_95844501_215C;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:78 GQ:4.5 PL:[0.0, 4.5, 198.0] SR:5 DR:0 LR:4.627 LO:8.689);ALT=G[chr8:95837120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	95908157	+	chr8	95970219	+	.	7	1	3978596_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAGGT;MAPQ=60;MATEID=3978596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_95966501_95991501_349C;SPAN=62062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:48 GQ:10.1 PL:[10.1, 0.0, 105.8] SR:1 DR:7 LR:-10.1 LO:14.8);ALT=T[chr8:95970219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	96146259	+	chr8	96166258	+	.	5	5	3979336_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3979336_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_96162501_96187501_305C;SPAN=19999;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:5 DR:5 LR:-21.04 LO:21.94);ALT=G[chr8:96166258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
