chr19	15014164	+	chr19	14962883	+	.	22	0	10180105_1	59.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=10180105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14962883(-)-19:15014164(+)__19_14994001_15019001D;SPAN=51281;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:47 GQ:53.3 PL:[59.9, 0.0, 53.3] SR:0 DR:22 LR:-59.9 LO:59.9);ALT=]chr19:15014164]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	14963098	+	chr19	15014280	+	.	16	0	10180106_1	36.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=10180106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14963098(+)-19:15014280(-)__19_14994001_15019001D;SPAN=51182;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:61 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:0 DR:16 LR:-36.29 LO:38.43);ALT=G[chr19:15014280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15046392	+	chr19	15049478	+	.	46	50	10180811_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=10180811_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_15043001_15068001_313C;SPAN=3086;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:70 GQ:21 PL:[231.0, 21.0, 0.0] SR:50 DR:46 LR:-231.1 LO:231.1);ALT=T[chr19:15049478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15965990	+	chr19	15967283	-	.	10	0	10185223_1	0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=10185223_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:15965990(+)-19:15967283(+)__19_15949501_15974501D;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:177 GQ:14.8 PL:[0.0, 14.8, 458.8] SR:0 DR:10 LR:14.94 LO:16.81);ALT=G]chr19:15967283];VARTYPE=BND:INV-hh;JOINTYPE=hh
