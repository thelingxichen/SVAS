chr9	83967925	+	chr9	83970684	+	.	47	39	4298543_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTTATAGC;MAPQ=60;MATEID=4298543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_83961501_83986501_138C;SPAN=2759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:39 DR:47 LR:-208.0 LO:208.0);ALT=C[chr9:83970684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	84324363	+	chr9	84326927	+	.	128	47	4300292_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TAAAATGGCTCTAGC;MAPQ=60;MATEID=4300292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_84304501_84329501_398C;SPAN=2564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:152 DP:897 GQ:99 PL:[258.9, 0.0, 1919.0] SR:47 DR:128 LR:-258.7 LO:332.3);ALT=C[chr9:84326927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
