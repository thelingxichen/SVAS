chr6	82460190	+	chr6	82461306	+	.	5	3	2919459_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2919459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_82442501_82467501_131C;SPAN=1116;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:93 GQ:1.8 PL:[0.0, 1.8, 227.7] SR:3 DR:5 LR:2.089 LO:12.67);ALT=T[chr6:82461306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	82950561	+	chr6	82957277	+	.	0	8	2920671_1	11.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=2920671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_82957001_82982001_278C;SPAN=6716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:8 DR:0 LR:-10.97 LO:16.77);ALT=C[chr6:82957277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
