chr16	29669312	-	chr16	29670574	+	.	9	0	9258140_1	8.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=9258140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:29669312(-)-16:29670574(-)__16_29645001_29670001D;SPAN=1262;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-7.764 LO:17.89);ALT=[chr16:29670574[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
