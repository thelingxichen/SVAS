chr17	29447482	+	chr12	145803	+	.	30	0	7315287_1	59.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7315287_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:145803(-)-17:29447482(+)__12_122501_147501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:145 GQ:59.9 PL:[59.9, 0.0, 290.9] SR:0 DR:30 LR:-59.75 LO:68.49);ALT=]chr17:29447482]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	66002065	+	chr16	24423747	+	.	36	0	9779643_1	99.0	.	DISC_MAPQ=8;EVDNC=DSCRD;IMPRECISE;MAPQ=8;MATEID=9779643_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:24423747(-)-17:66002065(+)__17_65978501_66003501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:65 GQ:55.1 PL:[101.3, 0.0, 55.1] SR:0 DR:36 LR:-101.9 LO:101.9);ALT=]chr17:66002065]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	25340111	+	chr16	25343128	+	.	182	118	9234294_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=9234294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_25333001_25358001_29C;SPAN=3017;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:248 DP:42 GQ:67 PL:[736.0, 67.0, 0.0] SR:118 DR:182 LR:-736.1 LO:736.1);ALT=G[chr16:25343128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29494702	+	chr17	29456776	+	G	61	45	9591705_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=9591705_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_29449001_29474001_546C;SPAN=37926;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:82 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:45 DR:61 LR:-244.3 LO:244.3);ALT=]chr17:29494702]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	29591282	+	chr17	29532860	+	.	60	16	9591938_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTA;MAPQ=60;MATEID=9591938_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_29571501_29596501_120C;SPAN=58422;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:59 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:16 DR:60 LR:-204.7 LO:204.7);ALT=]chr17:29591282]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	30433479	+	chr17	65925559	+	AGCAACAGTCACAGGC	0	10	9596509_1	14.0	.	EVDNC=ASSMB;INSERTION=AGCAACAGTCACAGGC;MAPQ=60;MATEID=9596509_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30429001_30454001_365C;SPAN=35492080;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:10 DR:0 LR:-13.77 LO:20.98);ALT=C[chr17:65925559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66660493	-	chr17	66690167	+	.	47	13	9781991_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=19;MATEID=9781991_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_66640001_66665001_155C;SPAN=29674;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:54 DP:84 GQ:46.7 PL:[155.6, 0.0, 46.7] SR:13 DR:47 LR:-158.6 LO:158.6);ALT=[chr17:66690167[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	66690062	+	chr17	66767168	-	.	34	36	9782455_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=9782455_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_66762501_66787501_41C;SPAN=77106;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:61 DP:74 GQ:3.3 PL:[184.8, 3.3, 0.0] SR:36 DR:34 LR:-193.0 LO:193.0);ALT=A]chr17:66767168];VARTYPE=BND:INV-hh;JOINTYPE=hh
