chrX	144422077	+	chrX	144424506	+	.	53	43	7546580_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7546580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_144403001_144428001_190C;SPAN=2429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:19 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:43 DR:53 LR:-221.2 LO:221.2);ALT=G[chrX:144424506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
