chr2	221278223	-	chr5	39787751	+	G	19	40	3385413_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=3385413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_39763501_39788501_343C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:92 GQ:71 PL:[150.2, 0.0, 71.0] SR:40 DR:19 LR:-151.5 LO:151.5);ALT=[chr5:39787751[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	222232064	+	chr2	222230960	+	.	36	0	1706211_1	91.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=1706211_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:222230960(-)-2:222232064(+)__2_222215001_222240001D;SPAN=1104;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:101 GQ:91.7 PL:[91.7, 0.0, 151.1] SR:0 DR:36 LR:-91.47 LO:92.34);ALT=]chr2:222232064]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	130625059	+	chr5	39787751	+	G	27	79	3385508_1	99.0	.	DISC_MAPQ=8;EVDNC=ASDIS;INSERTION=G;MAPQ=34;MATEID=3385508_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_39763501_39788501_418C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:92 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:79 DR:27 LR:-274.0 LO:274.0);ALT=]chr10:130625059]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	40020850	+	chr22	29065259	+	.	12	27	10865002_1	87.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=10865002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_29057001_29082001_291C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:32 DP:67 GQ:74.3 PL:[87.5, 0.0, 74.3] SR:27 DR:12 LR:-87.53 LO:87.53);ALT=G[chr22:29065259[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	40845844	-	chr5	40851278	+	.	49	47	3389996_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAA;MAPQ=60;MATEID=3389996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_40841501_40866501_442C;SPAN=5434;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:85 DP:121 GQ:43.4 PL:[248.0, 0.0, 43.4] SR:47 DR:49 LR:-255.7 LO:255.7);ALT=[chr5:40851278[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	40848797	+	chr5	40851277	+	.	8	0	3390011_1	9.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3390011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:40848797(+)-5:40851277(-)__5_40841501_40866501D;SPAN=2480;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=T[chr5:40851277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	9122379	+	chr9	9532385	+	CT	61	33	5778827_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CT;MAPQ=60;MATEID=5778827_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_9530501_9555501_23C;SPAN=410006;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:8 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:33 DR:61 LR:-237.7 LO:237.7);ALT=T[chr9:9532385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	18918573	+	chr9	9472190	+	.	8	25	5778759_1	85.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=T;MAPQ=41;MATEID=5778759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_9457001_9482001_5C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:2 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:25 DR:8 LR:-85.82 LO:85.82);ALT=]chr11:18918573]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	9557816	+	chr9	9786265	+	.	83	52	5778844_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5778844_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_9775501_9800501_15C;SPAN=228449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:10 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:52 DR:83 LR:-340.0 LO:340.0);ALT=T[chr9:9786265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	129647116	+	chr9	10208236	+	.	29	0	6594799_1	82.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=6594799_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:10208236(-)-10:129647116(+)__10_129629501_129654501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:51 GQ:39.2 PL:[82.1, 0.0, 39.2] SR:0 DR:29 LR:-82.61 LO:82.61);ALT=]chr10:129647116]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	10208403	+	chr10	129647274	+	.	13	0	6594801_1	31.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6594801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:10208403(+)-10:129647274(-)__10_129629501_129654501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:44 GQ:31.1 PL:[31.1, 0.0, 74.0] SR:0 DR:13 LR:-30.99 LO:32.03);ALT=A[chr10:129647274[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	49808791	+	chr10	130186863	+	.	8	0	6597156_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6597156_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:130186863(-)-12:49808791(+)__10_130168501_130193501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=]chr12:49808791]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	18963939	+	chr11	18986247	+	CAGACGATGGCTGAAGGTTTTCCTTTGGAGA	15	63	6656458_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;INSERTION=CAGACGATGGCTGAAGGTTTTCCTTTGGAGA;MAPQ=60;MATEID=6656458_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_11_18963001_18988001_140C;SPAN=22308;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:86 GQ:3.3 PL:[214.5, 3.3, 0.0] SR:63 DR:15 LR:-224.8 LO:224.8);ALT=A[chr11:18986247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
