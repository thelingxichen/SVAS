chr11	58304493	-	chr11	58305977	+	.	8	0	6825826_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6825826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:58304493(-)-11:58305977(-)__11_58285501_58310501D;SPAN=1484;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:102 GQ:0.9 PL:[0.0, 0.9, 247.5] SR:0 DR:8 LR:1.226 LO:14.63);ALT=[chr11:58305977[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
