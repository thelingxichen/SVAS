chr2	21045871	+	chr2	21060956	+	TT	85	71	931164_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TT;MAPQ=60;MATEID=931164_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_21021001_21046001_115C;SPAN=15085;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:126 DP:15 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:71 DR:85 LR:-373.0 LO:373.0);ALT=C[chr2:21060956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
