chr2	212280144	+	chr4	150245257	+	.	12	23	1666022_1	91.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=T;MAPQ=36;MATEID=1666022_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_212268001_212293001_393C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:76 GQ:91.7 PL:[91.7, 0.0, 91.7] SR:23 DR:12 LR:-91.64 LO:91.65);ALT=T[chr4:150245257[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	149990582	+	chr4	149992578	+	.	53	44	2986950_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AACA;MAPQ=60;MATEID=2986950_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_149989001_150014001_22C;SPAN=1996;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:83 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:44 DR:53 LR:-244.3 LO:244.3);ALT=A[chr4:149992578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
