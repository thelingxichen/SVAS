chr21	40799339	+	chr21	40800829	-	.	0	4	10789100_1	0	.	EVDNC=ASSMB;HOMSEQ=GGTGGCTCACGCCTGTAATCCCA;MAPQ=60;MATEID=10789100_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40792501_40817501_203C;SPAN=1490;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:141 GQ:24.6 PL:[0.0, 24.6, 389.4] SR:4 DR:0 LR:25.0 LO:5.515);ALT=A]chr21:40800829];VARTYPE=BND:INV-hh;JOINTYPE=hh
