chr2	134966717	+	chr2	134970131	+	.	70	26	1005489_1	88.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGAACTGGCTTATTTTT;MAPQ=60;MATEID=1005489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_134946001_134971001_73C;SPAN=3414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:723 GQ:88.3 PL:[88.3, 0.0, 1666.0] SR:26 DR:70 LR:-88.01 LO:173.6);ALT=T[chr2:134970131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	135810057	+	chr2	135815579	+	.	14	3	1007149_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1007149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_135803501_135828501_47C;SPAN=5522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:85 GQ:29.9 PL:[29.9, 0.0, 175.1] SR:3 DR:14 LR:-29.79 LO:35.79);ALT=T[chr2:135815579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136289204	+	chr2	136360069	+	.	13	10	1008575_1	43.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1008575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136342501_136367501_185C;SPAN=70865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:48 GQ:43.1 PL:[43.1, 0.0, 72.8] SR:10 DR:13 LR:-43.11 LO:43.54);ALT=G[chr2:136360069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136499585	+	chr2	136511729	+	TGATGAACAGTCTACACAGATGGCTGCAAGTTGGGAAGATGATAAAGTTACAGAAGCATCTTCAAACAGTTTTGTTGCTATTAAAATCGATACCAAAAGTGAAGCCTGCCTACAGTTTTCACAAATCT	5	54	1008989_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGGTGA;INSERTION=TGATGAACAGTCTACACAGATGGCTGCAAGTTGGGAAGATGATAAAGTTACAGAAGCATCTTCAAACAGTTTTGTTGCTATTAAAATCGATACCAAAAGTGAAGCCTGCCTACAGTTTTCACAAATCT;MAPQ=60;MATEID=1008989_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_136489501_136514501_128C;SPAN=12144;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:110 GQ:99 PL:[151.7, 0.0, 115.4] SR:54 DR:5 LR:-152.0 LO:152.0);ALT=A[chr2:136511729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136499585	+	chr2	136505834	+	.	34	34	1008988_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGGTGA;MAPQ=60;MATEID=1008988_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_136489501_136514501_128C;SPAN=6249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:121 GQ:99 PL:[149.0, 0.0, 142.4] SR:34 DR:34 LR:-148.8 LO:148.8);ALT=A[chr2:136505834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136505939	+	chr2	136511729	+	TGAAGCCTGCCTACAGTTTTCACAAATCT	2	22	1009005_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGGTGA;INSERTION=TGAAGCCTGCCTACAGTTTTCACAAATCT;MAPQ=60;MATEID=1009005_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_136489501_136514501_128C;SPAN=5790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:85 GQ:56.3 PL:[56.3, 0.0, 148.7] SR:22 DR:2 LR:-56.2 LO:58.56);ALT=G[chr2:136511729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136511847	+	chr2	136513085	+	.	2	15	1009033_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1009033_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136489501_136514501_127C;SPAN=1238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:103 GQ:28.4 PL:[28.4, 0.0, 219.8] SR:15 DR:2 LR:-28.21 LO:36.95);ALT=G[chr2:136513085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136513262	+	chr2	136519386	+	.	3	56	1009117_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1009117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136514001_136539001_36C;SPAN=6124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:46 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:56 DR:3 LR:-171.6 LO:171.6);ALT=G[chr2:136519386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136528306	+	chr2	136529989	+	.	8	3	1009161_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1009161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136514001_136539001_271C;SPAN=1683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:3 DR:8 LR:-9.661 LO:18.26);ALT=G[chr2:136529989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136602256	+	chr2	136603807	+	.	2	2	1009318_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1009318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136587501_136612501_130C;SPAN=1551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:87 GQ:10.2 PL:[0.0, 10.2, 231.0] SR:2 DR:2 LR:10.37 LO:6.36);ALT=T[chr2:136603807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136664978	+	chr2	136668952	+	AATGCCTCCACCAGCATGAGGAGGGGCTCCAAAGCGGAAGGAATCAATGTAAGCCTTAATTTTCTCCAAAT	3	30	1009489_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AATGCCTCCACCAGCATGAGGAGGGGCTCCAAAGCGGAAGGAATCAATGTAAGCCTTAATTTTCTCCAAAT;MAPQ=60;MATEID=1009489_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_136661001_136686001_313C;SPAN=3974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:72 GQ:83 PL:[89.6, 0.0, 83.0] SR:30 DR:3 LR:-89.43 LO:89.43);ALT=C[chr2:136668952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136691562	+	chr2	136700948	+	.	0	17	1009745_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1009745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136685501_136710501_183C;SPAN=9386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:76 GQ:35.6 PL:[35.6, 0.0, 147.8] SR:17 DR:0 LR:-35.53 LO:39.47);ALT=T[chr2:136700948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136691581	+	chr2	136718965	+	.	10	0	1009746_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1009746_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:136691581(+)-2:136718965(-)__2_136685501_136710501D;SPAN=27384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:24 GQ:26.6 PL:[26.6, 0.0, 29.9] SR:0 DR:10 LR:-26.51 LO:26.53);ALT=A[chr2:136718965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136719070	+	chr2	136736843	+	.	0	22	1009656_1	60.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1009656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_136734501_136759501_29C;SPAN=17773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:44 GQ:44.3 PL:[60.8, 0.0, 44.3] SR:22 DR:0 LR:-60.81 LO:60.81);ALT=T[chr2:136736843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136736939	+	chr2	136742972	+	GTTTTTCTTGTGATTGTATCATTGAAGATATTCCATATCTCTCTTTAGCATAAT	18	33	1009665_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTTTTCTTGTGATTGTATCATTGAAGATATTCCATATCTCTCTTTAGCATAAT;MAPQ=60;MATEID=1009665_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_136734501_136759501_222C;SPAN=6033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:93 GQ:99 PL:[116.9, 0.0, 107.0] SR:33 DR:18 LR:-116.8 LO:116.8);ALT=G[chr2:136742972[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136741068	+	chr2	136743030	+	.	14	0	1009675_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1009675_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:136741068(+)-2:136743030(-)__2_136734501_136759501D;SPAN=1962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:106 GQ:17.6 PL:[17.6, 0.0, 238.7] SR:0 DR:14 LR:-17.5 LO:28.95);ALT=T[chr2:136743030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	136873517	+	chr2	136875657	+	.	26	0	1010027_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1010027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:136873517(+)-2:136875657(-)__2_136857001_136882001D;SPAN=2140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:100 GQ:58.7 PL:[58.7, 0.0, 184.1] SR:0 DR:26 LR:-58.73 LO:62.34);ALT=C[chr2:136875657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
