chrX	40440350	+	chrX	40450484	+	.	18	0	7404401_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7404401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:40440350(+)-23:40450484(-)__23_40449501_40474501D;SPAN=10134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:30 GQ:21.5 PL:[51.2, 0.0, 21.5] SR:0 DR:18 LR:-51.95 LO:51.95);ALT=G[chrX:40450484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	40440357	+	chrX	40448237	+	.	38	15	7404362_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGTG;MAPQ=60;MATEID=7404362_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_23_40425001_40450001_25C;SPAN=7880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:66 GQ:15.2 PL:[143.9, 0.0, 15.2] SR:15 DR:38 LR:-149.8 LO:149.8);ALT=G[chrX:40448237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	40448369	+	chrX	40450486	+	.	0	23	7404379_1	51.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=7404379_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_23_40425001_40450001_25C;SPAN=2117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:30 GQ:2.3 PL:[51.7, 0.0, 2.3] SR:23 DR:0 LR:-54.91 LO:54.91);ALT=G[chrX:40450486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	40450618	+	chrX	40456501	+	.	0	8	7404405_1	13.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7404405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_40449501_40474501_113C;SPAN=5883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:8 DR:0 LR:-13.4 LO:17.42);ALT=G[chrX:40456501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	40460133	+	chrX	40464812	+	.	4	7	7404424_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7404424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_40449501_40474501_209C;SPAN=4679;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:44 GQ:24.5 PL:[24.5, 0.0, 80.6] SR:7 DR:4 LR:-24.39 LO:26.15);ALT=G[chrX:40464812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	41198338	+	chrX	41200733	+	.	2	9	7405744_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AAAGGT;MAPQ=60;MATEID=7405744_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_41184501_41209501_105C;SPAN=2395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:9 DR:2 LR:-16.43 LO:20.02);ALT=T[chrX:41200733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
