chr9	113013744	+	chr9	113018692	+	.	111	56	4393134_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4393134_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_112994001_113019001_356C;SPAN=4948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:131 DP:155 GQ:15.4 PL:[405.9, 15.4, 0.0] SR:56 DR:111 LR:-418.5 LO:418.5);ALT=T[chr9:113018692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	113024576	+	chr9	113037094	+	TTATTATTATTAT	24	27	4392824_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TTATTATTATTAT;MAPQ=60;MATEID=4392824_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_113018501_113043501_251C;SPAN=12518;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:85 GQ:86 PL:[119.0, 0.0, 86.0] SR:27 DR:24 LR:-119.2 LO:119.2);ALT=T[chr9:113037094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	113037287	+	chr9	113029970	+	.	53	41	4392839_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=4392839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_113018501_113043501_328C;SPAN=7317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:97 GQ:3 PL:[240.9, 3.0, 0.0] SR:41 DR:53 LR:-253.2 LO:253.2);ALT=]chr9:113037287]A;VARTYPE=BND:DUP-th;JOINTYPE=th
