chr16	1787978	+	chr16	1786539	+	.	20	0	9119108_1	49.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=9119108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1786539(-)-16:1787978(+)__16_1764001_1789001D;SPAN=1439;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:63 GQ:49.1 PL:[49.1, 0.0, 101.9] SR:0 DR:20 LR:-48.95 LO:50.04);ALT=]chr16:1787978]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	1789744	+	chr16	1788455	+	.	10	0	9118926_1	16.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=9118926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1788455(-)-16:1789744(+)__16_1788501_1813501D;SPAN=1289;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:63 GQ:16.1 PL:[16.1, 0.0, 134.9] SR:0 DR:10 LR:-15.94 LO:21.55);ALT=]chr16:1789744]A;VARTYPE=BND:DUP-th;JOINTYPE=th
