chr18	2674144	+	chr18	2688390	+	.	0	9	6527733_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6527733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_2670501_2695501_91C;SPAN=14246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:9 DR:0 LR:-16.98 LO:20.21);ALT=G[chr18:2688390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3247908	+	chr18	3253230	+	.	107	9	6528746_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6528746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_3234001_3259001_228C;SPAN=5322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:151 GQ:38.6 PL:[325.7, 0.0, 38.6] SR:9 DR:107 LR:-338.3 LO:338.3);ALT=G[chr18:3253230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3247935	+	chr18	3253884	+	.	24	0	6528748_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6528748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:3247935(+)-18:3253884(-)__18_3234001_3259001D;SPAN=5949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:78 GQ:58.1 PL:[58.1, 0.0, 130.7] SR:0 DR:24 LR:-58.09 LO:59.65);ALT=G[chr18:3253884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3254049	+	chr18	3255743	+	.	13	39	6528761_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=13;MATEID=6528761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_3234001_3259001_270C;SPAN=1694;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:58 GQ:2.4 PL:[145.2, 2.4, 0.0] SR:39 DR:13 LR:-152.1 LO:152.1);ALT=G[chr18:3255743[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3262235	+	chr18	3272881	+	.	106	17	6528628_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6528628_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_3258501_3283501_75C;SPAN=10646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:97 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:17 DR:106 LR:-412.6 LO:412.6);ALT=G[chr18:3272881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3262268	+	chr18	3277248	+	.	15	0	6528629_1	35.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6528629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:3262268(+)-18:3277248(-)__18_3258501_3283501D;SPAN=14980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:51 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.7 LO:36.92);ALT=C[chr18:3277248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	3273081	+	chr18	3277249	+	.	4	88	6528649_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6528649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_3258501_3283501_205C;SPAN=4168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:66 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:88 DR:4 LR:-267.4 LO:267.4);ALT=G[chr18:3277249[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
