chr9	44761503	+	chr9	47166979	+	.	0	20	4220483_1	49.0	.	EVDNC=ASSMB;HOMSEQ=GAAACCCCGTCTC;MAPQ=57;MATEID=4220483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_44761501_44786501_678C;SPAN=2405476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:60 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:20 DR:0 LR:-49.76 LO:50.57);ALT=C[chr9:47166979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
