chr5	89821156	+	chr5	89825318	+	.	10	0	2526504_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2526504_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:89821156(+)-5:89825318(-)__5_89817001_89842001D;SPAN=4162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:0 DR:10 LR:-17.3 LO:21.94);ALT=G[chr5:89825318[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	90499775	+	chr5	90502096	+	.	71	43	2527373_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTA;MAPQ=60;MATEID=2527373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_90478501_90503501_112C;SPAN=2321;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:22 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:43 DR:71 LR:-270.7 LO:270.7);ALT=A[chr5:90502096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
