chr5	102873209	-	chrX	107025423	+	.	9	7	3651443_1	47.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATAAATATATATATATAAATATATATATA;MAPQ=60;MATEID=3651443_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_5_102851001_102876001_117C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:21 GQ:1.1 PL:[47.3, 0.0, 1.1] SR:7 DR:9 LR:-49.3 LO:49.3);ALT=[chrX:107025423[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	103854288	+	chr5	103860327	+	.	51	27	3654870_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AATAAAATTATTAA;MAPQ=60;MATEID=3654870_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_103855501_103880501_58C;SPAN=6039;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:37 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:27 DR:51 LR:-191.4 LO:191.4);ALT=A[chr5:103860327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
