chr9	94384636	+	chr1	219648974	+	.	19	29	829805_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGAAAGAAAGAGAGAAAGAAAGAGAGAAAGAAAGA;MAPQ=46;MATEID=829805_2;MATENM=0;NM=14;NUMPARTS=2;SCTG=c_1_219642501_219667501_46C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:40 DP:12 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:29 DR:19 LR:-118.8 LO:118.8);ALT=]chr9:94384636]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	219897105	+	chrX	45536829	-	.	2	55	11133402_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=11133402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_45521001_45546001_1C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:79 GQ:31.4 PL:[160.1, 0.0, 31.4] SR:55 DR:2 LR:-165.0 LO:165.0);ALT=A]chrX:45536829];VARTYPE=BND:TRX-hh;JOINTYPE=hh
