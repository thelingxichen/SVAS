chr3	133503782	+	chr3	133505083	+	.	103	96	2333729_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AACAATACTATTTTTT;MAPQ=60;MATEID=2333729_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_133500501_133525501_147C;SPAN=1301;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:162 DP:42 GQ:43.6 PL:[478.6, 43.6, 0.0] SR:96 DR:103 LR:-478.6 LO:478.6);ALT=T[chr3:133505083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
