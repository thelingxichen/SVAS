chr2	89043877	+	chr3	189959380	-	.	13	0	2566252_1	33.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=2566252_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:89043877(+)-3:189959380(+)__3_189948501_189973501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:36 GQ:33.2 PL:[33.2, 0.0, 53.0] SR:0 DR:13 LR:-33.16 LO:33.44);ALT=C]chr3:189959380];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	89831994	+	chr2	89833326	+	.	0	38	1166847_1	33.0	.	EVDNC=ASSMB;HOMSEQ=TGATGATTCCATTCGA;MAPQ=60;MATEID=1166847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_89817001_89842001_100C;SPAN=1332;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:38 DP:340 GQ:33.3 PL:[33.3, 0.0, 792.5] SR:38 DR:0 LR:-33.32 LO:75.63);ALT=A[chr2:89833326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	90296133	+	chr2	90294967	+	.	16	0	1163486_1	12.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=1163486_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:90294967(-)-2:90296133(+)__2_90282501_90307501D;SPAN=1166;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:150 GQ:12.2 PL:[12.2, 0.0, 352.1] SR:0 DR:16 LR:-12.18 LO:31.5);ALT=]chr2:90296133]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	186581033	+	chr3	186585285	+	.	110	74	2552097_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAAAAATATTGCAAATAG;MAPQ=60;MATEID=2552097_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_3_186567501_186592501_446C;SPAN=4252;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:143 DP:50 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:74 DR:110 LR:-422.5 LO:422.5);ALT=G[chr3:186585285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	187085160	-	chr22	30993411	+	.	11	14	2553730_1	42.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=CACCAATCAGCACCCTGTGTCTAGCTCA;MAPQ=22;MATEID=2553730_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_187082001_187107001_209C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:76 GQ:42.2 PL:[42.2, 0.0, 141.2] SR:14 DR:11 LR:-42.13 LO:45.17);ALT=[chr22:30993411[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	187766589	-	chr3	187768477	+	.	9	0	2556582_1	12.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2556582_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:187766589(-)-3:187768477(-)__3_187768001_187793001D;SPAN=1888;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=[chr3:187768477[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	188596563	+	chr3	188597836	-	.	2	12	2560429_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAA;MAPQ=60;MATEID=2560429_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_188576501_188601501_67C;SPAN=1273;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:122 GQ:13.4 PL:[13.4, 0.0, 280.7] SR:12 DR:2 LR:-13.16 LO:28.03);ALT=A]chr3:188597836];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	189159362	+	chr3	188912760	+	.	3	6	2562640_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2562640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_189140001_189165001_299C;SPAN=246602;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:6 DR:3 LR:-3.059 LO:13.4);ALT=]chr3:189159362]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	189363422	+	chr3	189370900	+	.	118	105	2563202_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=54;MATEID=2563202_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_3_189360501_189385501_227C;SPAN=7478;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:181 DP:47 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:105 DR:118 LR:-534.7 LO:534.7);ALT=T[chr3:189370900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	189737348	+	chr3	189740525	+	.	111	100	2564519_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CTCA;MAPQ=60;MATEID=2564519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_189728001_189753001_91C;SPAN=3177;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:168 DP:38 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:100 DR:111 LR:-498.4 LO:498.4);ALT=A[chr3:189740525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	86954348	+	chr22	31700285	+	.	4	2	8656840_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8656840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_86950501_86975501_91C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:2 DR:4 LR:4.677 LO:6.851);ALT=T[chr22:31700285[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr15	77951478	+	chr15	77654406	+	TG	83	42	9000517_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TG;MAPQ=60;MATEID=9000517_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_77934501_77959501_70C;SPAN=297072;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:83 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:42 DR:83 LR:-316.9 LO:316.9);ALT=]chr15:77951478]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	78892128	+	chr22	31416873	+	.	36	66	9006549_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAATCCTAGCACTTTGGGAGGCCAAGGC;MAPQ=60;MATEID=9006549_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_78890001_78915001_522C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:50 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:66 DR:36 LR:-280.6 LO:280.6);ALT=C[chr22:31416873[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
