chr22	36702256	+	chr22	36782505	+	.	8	0	10882833_1	20.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=10882833_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36702256(+)-22:36782505(-)__22_36774501_36799501D;SPAN=80249;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:23 GQ:20.3 PL:[20.3, 0.0, 33.5] SR:0 DR:8 LR:-20.18 LO:20.41);ALT=G[chr22:36782505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36816796	-	chr22	36817855	+	.	9	0	10882991_1	12.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=10882991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36816796(-)-22:36817855(-)__22_36799001_36824001D;SPAN=1059;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:0 DR:9 LR:-12.1 LO:18.81);ALT=[chr22:36817855[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	37143176	+	chr22	37147896	+	.	42	41	10883635_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGTAGCT;MAPQ=60;MATEID=10883635_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37142001_37167001_123C;SPAN=4720;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:21 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:41 DR:42 LR:-227.8 LO:227.8);ALT=T[chr22:37147896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
