chr9	29076010	+	chr9	29279559	+	.	17	0	5808682_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5808682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:29076010(+)-9:29279559(-)__9_29277501_29302501D;SPAN=203549;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:17 DP:10 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:17 LR:-49.51 LO:49.51);ALT=C[chr9:29279559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	29076945	+	chr9	29279560	+	TTTT	50	58	5808684_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;INSERTION=TTTT;MAPQ=60;MATEID=5808684_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_9_29277501_29302501_1C;SPAN=202615;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:11 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:58 DR:50 LR:-257.5 LO:257.5);ALT=A[chr9:29279560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	29505454	+	chr9	29507054	+	.	51	39	5809066_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5809066_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_29498001_29523001_218C;SPAN=1600;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:20 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:39 DR:51 LR:-208.0 LO:208.0);ALT=T[chr9:29507054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
