chr6	95193324	+	chr6	95194337	+	.	57	45	2947499_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=2947499_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_95182501_95207501_153C;SPAN=1013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:21 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:45 DR:57 LR:-247.6 LO:247.6);ALT=A[chr6:95194337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	96025514	+	chr6	96034277	+	.	5	6	2948798_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2948798_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_96015501_96040501_277C;SPAN=8763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:6 DR:5 LR:-5.818 LO:15.7);ALT=G[chr6:96034277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	96969811	+	chr6	96971018	+	.	10	0	2950889_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2950889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:96969811(+)-6:96971018(-)__6_96946501_96971501D;SPAN=1207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:0 DR:10 LR:-9.44 LO:20.03);ALT=C[chr6:96971018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
