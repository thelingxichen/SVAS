chr17	44249604	+	chr17	44270187	+	.	9	0	6411908_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6411908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:44249604(+)-17:44270187(-)__17_44247001_44272001D;SPAN=20583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=A[chr17:44270187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	44271105	+	chr17	44273732	+	.	0	28	6412104_1	77.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6412104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_44271501_44296501_179C;SPAN=2627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:55 GQ:54.5 PL:[77.6, 0.0, 54.5] SR:28 DR:0 LR:-77.71 LO:77.71);ALT=G[chr17:44273732[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
