chr12	24223450	+	chr12	24206281	+	.	47	36	7476535_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CTC;MAPQ=60;MATEID=7476535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_24206001_24231001_283C;SPAN=17169;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:73 DP:197 GQ:99 PL:[187.7, 0.0, 290.0] SR:36 DR:47 LR:-187.6 LO:188.8);ALT=]chr12:24223450]C;VARTYPE=BND:DUP-th;JOINTYPE=th
