chr1	229552128	+	chr1	231967699	-	.	28	0	857257_1	78.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=857257_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:229552128(+)-1:231967699(+)__1_231966001_231991001D;SPAN=2415571;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:51 GQ:42.5 PL:[78.8, 0.0, 42.5] SR:0 DR:28 LR:-79.1 LO:79.1);ALT=T]chr1:231967699];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	229552761	-	chr1	231967021	+	.	10	0	857259_1	23.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=857259_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:229552761(-)-1:231967021(-)__1_231966001_231991001D;SPAN=2414260;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=[chr1:231967021[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
