chrX	143406976	+	chrX	143409979	+	TAC	34	23	7545516_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=TAC;MAPQ=60;MATEID=7545516_2;MATENM=4;NM=1;NUMPARTS=3;REPSEQ=AGAAGA;SCTG=c_23_143398501_143423501_249C;SPAN=3003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:23 GQ:13.1 PL:[114.4, 13.1, 0.0] SR:23 DR:34 LR:-114.4 LO:114.4);ALT=A[chrX:143409979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	143406976	+	chrX	143410375	+	TACGCACTATTTGGATGCAATTTTTGGGACTTAATATGTGTTATACACTTTTATTTTAAAATATTTATTTACTTGAAATTCAACTTTAACTTGGTGTCCTATATTTTATCTGGCAATTCTATTGCTATAAGATGGGGCATCTGTTAAAGAATTGTATCTTAGCTCATGAGAGGCTGCCAAGCCACCTGAATTATTCCTTACGTCACCCCCCTGAGGCACACAATCCTTATTCACCATGGGCTCTACAATAAGCAGTTTATTCGATACACATCTACATAAACTTACTTCTGTAAGTACTAAGTACT	2	56	7545517_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;INSERTION=TACGCACTATTTGGATGCAATTTTTGGGACTTAATATGTGTTATACACTTTTATTTTAAAATATTTATTTACTTGAAATTCAACTTTAACTTGGTGTCCTATATTTTATCTGGCAATTCTATTGCTATAAGATGGGGCATCTGTTAAAGAATTGTATCTTAGCTCATGAGAGGCTGCCAAGCCACCTGAATTATTCCTTACGTCACCCCCCTGAGGCACACAATCCTTATTCACCATGGGCTCTACAATAAGCAGTTTATTCGATACACATCTACATAAACTTACTTCTGTAAGTACTAAGTACT;MAPQ=60;MATEID=7545517_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_23_143398501_143423501_249C;SPAN=3399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:14 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:56 DR:2 LR:-171.6 LO:171.6);ALT=A[chrX:143410375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
