chr3	103191898	+	chr3	103193053	-	.	8	0	2210044_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2210044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:103191898(+)-3:103193053(+)__3_103169501_103194501D;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:157 GQ:16 PL:[0.0, 16.0, 412.6] SR:0 DR:8 LR:16.13 LO:13.08);ALT=G]chr3:103193053];VARTYPE=BND:INV-hh;JOINTYPE=hh
