chr4	128474248	+	chr4	128430569	+	AAGAT	16	13	2906431_1	66.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAGAT;MAPQ=60;MATEID=2906431_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_128429001_128454001_3C;SPAN=43679;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:26 DP:70 GQ:66.8 PL:[66.8, 0.0, 103.1] SR:13 DR:16 LR:-66.86 LO:67.28);ALT=]chr4:128474248]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	128443510	-	chrX	124724260	+	.	6	5	11373344_1	26.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=11373344_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_124705001_124730001_207C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:5 DR:6 LR:-26.24 LO:26.3);ALT=[chrX:124724260[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	128456129	+	chr4	128465497	+	AA	5	6	2906231_1	0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=AA;MAPQ=60;MATEID=2906231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_128453501_128478501_341C;SPAN=9368;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:166 GQ:11.8 PL:[0.0, 11.8, 425.8] SR:6 DR:5 LR:11.96 LO:17.1);ALT=T[chr4:128465497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
