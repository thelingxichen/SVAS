chr11	28119463	+	chr11	28129610	+	.	9	0	4803033_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4803033_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:28119463(+)-11:28129610(-)__11_28126001_28151001D;SPAN=10147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=T[chr11:28129610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
