chr6	64131099	-	chr6	64132185	+	.	8	0	4245206_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4245206_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:64131099(-)-6:64132185(-)__6_64116501_64141501D;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:174 GQ:20.5 PL:[0.0, 20.5, 462.1] SR:0 DR:8 LR:20.73 LO:12.72);ALT=[chr6:64132185[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
