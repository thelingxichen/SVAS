chr17	67524784	-	chr17	67525866	+	.	5	2	6480992_1	0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=TGGTCTCGATCTCCTGACCTC;MAPQ=0;MATEID=6480992_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_67522001_67547001_300C;SPAN=1082;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:78 GQ:1.2 PL:[0.0, 1.2, 191.4] SR:2 DR:5 LR:1.326 LO:10.92);ALT=[chr17:67525866[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	68455097	+	chr17	68461177	+	.	68	23	6483779_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAGATTTTGTG;MAPQ=60;MATEID=6483779_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_68453001_68478001_89C;SPAN=6080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:402 GQ:99 PL:[162.0, 0.0, 812.3] SR:23 DR:68 LR:-161.8 LO:186.6);ALT=G[chr17:68461177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
