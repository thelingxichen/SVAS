chr9	69513477	+	chr2	95406469	+	.	8	0	5877061_1	10.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=5877061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:95406469(-)-9:69513477(+)__9_69506501_69531501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=]chr9:69513477]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	68411489	+	chr9	68414114	+	CTTGCTGCCTGGCTCAT	56	40	5874421_1	99.0	.	DISC_MAPQ=11;EVDNC=ASDIS;INSERTION=CTTGCTGCCTGGCTCAT;MAPQ=49;MATEID=5874421_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_9_68404001_68429001_439C;SPAN=2625;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:84 DP:358 GQ:99 PL:[180.4, 0.0, 688.7] SR:40 DR:56 LR:-180.3 LO:197.0);ALT=C[chr9:68414114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	68514095	+	chr9	69002875	-	.	8	0	5875314_1	10.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=5875314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:68514095(+)-9:69002875(+)__9_68992001_69017001D;SPAN=488780;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=G]chr9:69002875];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	69986659	+	chr9	69985437	+	.	8	0	5878703_1	2.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=5878703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:69985437(-)-9:69986659(+)__9_69972001_69997001D;SPAN=1222;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=]chr9:69986659]T;VARTYPE=BND:DUP-th;JOINTYPE=th
