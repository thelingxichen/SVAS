chr15	36826996	+	chr15	36828426	-	.	8	0	8850910_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=8850910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:36826996(+)-15:36828426(+)__15_36823501_36848501D;SPAN=1430;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:139 GQ:11.1 PL:[0.0, 11.1, 359.7] SR:0 DR:8 LR:11.25 LO:13.52);ALT=A]chr15:36828426];VARTYPE=BND:INV-hh;JOINTYPE=hh
