chr2	87545606	+	chr2	112300777	+	.	5	4	1258607_1	8.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGGCACAGTGGC;MAPQ=60;MATEID=1258607_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_112283501_112308501_338C;SPAN=24755171;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:4 DR:5 LR:-8.035 LO:17.94);ALT=C[chr2:112300777[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	87588026	+	chr2	87586943	+	.	31	0	1149421_1	35.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=1149421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:87586943(-)-2:87588026(+)__2_87563001_87588001D;SPAN=1083;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:246 GQ:35.8 PL:[35.8, 0.0, 560.6] SR:0 DR:31 LR:-35.68 LO:63.42);ALT=]chr2:87588026]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	111983099	+	chr2	111982009	+	.	44	0	1256203_1	74.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=1256203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:111982009(-)-2:111983099(+)__2_111965001_111990001D;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:263 GQ:74.2 PL:[74.2, 0.0, 562.7] SR:0 DR:44 LR:-73.99 LO:95.91);ALT=]chr2:111983099]T;VARTYPE=BND:DUP-th;JOINTYPE=th
