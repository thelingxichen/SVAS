chr7	146413149	+	chr7	146414636	+	A	56	39	5316448_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=5316448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_146412001_146437001_34C;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:19 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:39 DR:56 LR:-234.4 LO:234.4);ALT=T[chr7:146414636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	146413149	+	chr7	146415074	-	T	9	39	5316449_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=5316449_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_146412001_146437001_162C;SPAN=1925;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:47 DP:37 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:39 DR:9 LR:-138.6 LO:138.6);ALT=T]chr7:146415074];VARTYPE=BND:INV-hh;JOINTYPE=hh
