chrX	62652372	+	chrX	62780710	+	.	0	19	7434321_1	53.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=7434321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_62769001_62794001_6C;SPAN=128338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:34 GQ:27.2 PL:[53.6, 0.0, 27.2] SR:19 DR:0 LR:-53.9 LO:53.9);ALT=C[chrX:62780710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
