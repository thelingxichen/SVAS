chr8	580472	+	chr8	579162	+	.	23	0	5365959_1	57.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5365959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:579162(-)-8:580472(+)__8_563501_588501D;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:67 GQ:57.8 PL:[57.8, 0.0, 104.0] SR:0 DR:23 LR:-57.77 LO:58.52);ALT=]chr8:580472]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	594397	+	chr8	599415	+	CAA	59	45	5365843_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CAA;MAPQ=60;MATEID=5365843_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_588001_613001_185C;SPAN=5018;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:18 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:45 DR:59 LR:-250.9 LO:250.9);ALT=G[chr8:599415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	1409564	+	chr8	1410705	+	.	40	0	5367707_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=5367707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:1409564(+)-8:1410705(-)__8_1396501_1421501D;SPAN=1141;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:40 DP:26 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:40 LR:-118.8 LO:118.8);ALT=G[chr8:1410705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	2284948	+	chr8	2329100	-	.	15	0	5369469_1	43.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5369469_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:2284948(+)-8:2329100(+)__8_2327501_2352501D;SPAN=44152;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:22 GQ:7.4 PL:[43.7, 0.0, 7.4] SR:0 DR:15 LR:-44.75 LO:44.75);ALT=G]chr8:2329100];VARTYPE=BND:INV-hh;JOINTYPE=hh
