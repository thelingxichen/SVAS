chr4	21161002	+	chr4	21167098	+	.	52	39	2651539_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAAATTATACTAAA;MAPQ=60;MATEID=2651539_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_21143501_21168501_217C;SPAN=6096;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:22 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:39 DR:52 LR:-208.0 LO:208.0);ALT=A[chr4:21167098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
