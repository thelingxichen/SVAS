chr18	59672786	+	chr18	59674185	+	.	52	9	6647277_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCACAACATGGGGGAATTCTGGGAGATACAATTCAAGTTGAGATTTGGGTGGGGACACAGC;MAPQ=60;MATEID=6647277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_59657501_59682501_179C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:35 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:9 DR:52 LR:-178.2 LO:178.2);ALT=C[chr18:59674185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	60247770	+	chr18	60249068	+	.	8	0	6648694_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6648694_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:60247770(+)-18:60249068(-)__18_60245501_60270501D;SPAN=1298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:126 GQ:7.5 PL:[0.0, 7.5, 320.1] SR:0 DR:8 LR:7.729 LO:13.87);ALT=A[chr18:60249068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	61027027	+	chr18	61034242	+	CATTTCGTGCAACCAGAGTTATAAAAGCTCCTTGTTTATAGCACTCGATAGCAATGCACTTCCCGATGCCACTGGAACCTCCTGTA	0	11	6650777_1	24.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=CATTTCGTGCAACCAGAGTTATAAAAGCTCCTTGTTTATAGCACTCGATAGCAATGCACTTCCCGATGCCACTGGAACCTCCTGTA;MAPQ=60;MATEID=6650777_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_61005001_61030001_338C;SPAN=7215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:44 GQ:24.5 PL:[24.5, 0.0, 80.6] SR:11 DR:0 LR:-24.39 LO:26.15);ALT=T[chr18:61034242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	61077679	+	chr18	61089466	+	ATTTAACGACATGAAGAAAATACTGCACAGCATGCTGATAGAGCTGAAGGGCTTCTTCGTAGTTCCCAGCCTTGTCTTCTTGCGCTGCTTTGCTAGCCAGATCTATCGCTTT	0	23	6650846_1	66.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATTTAACGACATGAAGAAAATACTGCACAGCATGCTGATAGAGCTGAAGGGCTTCTTCGTAGTTCCCAGCCTTGTCTTCTTGCGCTGCTTTGCTAGCCAGATCTATCGCTTT;MAPQ=60;MATEID=6650846_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_61054001_61079001_20C;SPAN=11787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:36 GQ:20 PL:[66.2, 0.0, 20.0] SR:23 DR:0 LR:-67.45 LO:67.45);ALT=T[chr18:61089466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	61078814	+	chr18	61089466	+	.	0	19	6650930_1	41.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6650930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_61078501_61103501_148C;SPAN=10652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:78 GQ:41.6 PL:[41.6, 0.0, 147.2] SR:19 DR:0 LR:-41.59 LO:44.92);ALT=G[chr18:61089466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
