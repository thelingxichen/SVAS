chr6	68101533	+	chr6	68112167	+	.	87	32	2888076_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2888076_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_6_68110001_68135001_266C;SPAN=10634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:50 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:32 DR:87 LR:-303.7 LO:303.7);ALT=T[chr6:68112167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
