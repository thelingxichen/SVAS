chr2	196522128	+	chr2	196544764	+	.	8	0	1146883_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1146883_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:196522128(+)-2:196544764(-)__2_196514501_196539501D;SPAN=22636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=G[chr2:196544764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	197002453	+	chr2	197004343	+	.	13	8	1148298_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1148298_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_197004501_197029501_35C;SPAN=1890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:0 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:8 DR:13 LR:-52.81 LO:52.81);ALT=C[chr2:197004343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	197004524	+	chr2	197008284	+	ACATATCTGTTGCTGTGGTAATGGGATCATAGTTCAGGATTTCTGGAG	7	15	1148300_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ACATATCTGTTGCTGTGGTAATGGGATCATAGTTCAGGATTTCTGGAG;MAPQ=60;MATEID=1148300_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_197004501_197029501_102C;SPAN=3760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:74 GQ:36.2 PL:[36.2, 0.0, 141.8] SR:15 DR:7 LR:-36.07 LO:39.69);ALT=C[chr2:197008284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	197010779	+	chr2	197021163	+	.	5	6	1148317_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1148317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_197004501_197029501_28C;SPAN=10384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:82 GQ:7.7 PL:[7.7, 0.0, 189.2] SR:6 DR:5 LR:-7.493 LO:17.84);ALT=A[chr2:197021163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	197021371	+	chr2	197027986	+	ACCT	3	5	1148350_1	1.0	.	DISC_MAPQ=40;EVDNC=ASDIS;INSERTION=ACCT;MAPQ=60;MATEID=1148350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_197004501_197029501_99C;SPAN=6615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:80 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:5 DR:3 LR:-1.433 LO:13.15);ALT=T[chr2:197027986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	197028152	+	chr2	197036055	+	.	29	41	1148368_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1148368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_197004501_197029501_57C;SPAN=7903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:53 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:41 DR:29 LR:-168.3 LO:168.3);ALT=C[chr2:197036055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
