chr20	7964505	+	chr20	7967933	+	.	4	9	6910942_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=6910942_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_20_7962501_7987501_24C;SPAN=3428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:103 GQ:8.6 PL:[8.6, 0.0, 239.6] SR:9 DR:4 LR:-8.406 LO:21.66);ALT=C[chr20:7967933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	7968037	+	chr20	7980378	+	CATATCTTGCCAGAGATGCTAAAAAGACCAGCCATTCCAGACAT	0	13	6910955_1	15.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATATCTTGCCAGAGATGCTAAAAAGACCAGCCATTCCAGACAT;MAPQ=60;MATEID=6910955_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_7962501_7987501_327C;SPAN=12341;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:13 DR:0 LR:-15.01 LO:26.61);ALT=C[chr20:7980378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	7990962	+	chr20	8000085	+	.	0	10	6911204_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6911204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_7987001_8012001_42C;SPAN=9123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:122 GQ:0.2 PL:[0.2, 0.0, 293.9] SR:10 DR:0 LR:0.04279 LO:18.48);ALT=A[chr20:8000085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
