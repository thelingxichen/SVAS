chr17	55255300	+	chr22	22249853	-	.	14	0	10849324_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10849324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55255300(+)-22:22249853(+)__22_22246001_22271001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:31 GQ:34.7 PL:[38.0, 0.0, 34.7] SR:0 DR:14 LR:-37.82 LO:37.82);ALT=A]chr22:22249853];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr17	55687811	+	chr17	55689915	+	.	171	100	9725777_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=9725777_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_17_55664001_55689001_271C;SPAN=2104;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:217 DP:19 GQ:58.6 PL:[643.6, 58.6, 0.0] SR:100 DR:171 LR:-643.7 LO:643.7);ALT=T[chr17:55689915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	56336685	+	chr17	56343665	+	.	58	47	9728620_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTGC;MAPQ=60;MATEID=9728620_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_56325501_56350501_305C;SPAN=6980;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:92 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:47 DR:58 LR:-270.7 LO:270.7);ALT=C[chr17:56343665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
