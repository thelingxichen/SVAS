chr2	35976021	+	chr2	35997157	+	.	30	0	750772_1	89.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=750772_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:35976021(+)-2:35997157(-)__2_35990501_36015501D;SPAN=21136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:31 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=A[chr2:35997157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	36806008	+	chr2	36808432	+	.	0	12	752652_1	16.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=752652_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_36799001_36824001_332C;SPAN=2424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:87 GQ:16.1 PL:[16.1, 0.0, 194.3] SR:12 DR:0 LR:-16.04 LO:25.06);ALT=C[chr2:36808432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37311762	+	chr2	37316782	+	.	10	0	754140_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=754140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:37311762(+)-2:37316782(-)__2_37313501_37338501D;SPAN=5020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:0 DR:10 LR:-22.44 LO:23.91);ALT=A[chr2:37316782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37375006	+	chr2	37384048	+	.	11	0	754262_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=754262_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:37375006(+)-2:37384048(-)__2_37362501_37387501D;SPAN=9042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:0 DR:11 LR:-13.82 LO:22.76);ALT=A[chr2:37384048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37376319	+	chr2	37384050	+	.	12	0	754266_1	14.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=754266_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:37376319(+)-2:37384050(-)__2_37362501_37387501D;SPAN=7731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:94 GQ:14.3 PL:[14.3, 0.0, 212.3] SR:0 DR:12 LR:-14.15 LO:24.62);ALT=T[chr2:37384050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37426962	+	chr2	37428783	+	TCCAAGATGAAGGGATATTTCTTGCTCATTGTTTGCCTGAAAT	34	48	754441_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TCCAAGATGAAGGGATATTTCTTGCTCATTGTTTGCCTGAAAT;MAPQ=60;MATEID=754441_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_37411501_37436501_234C;SPAN=1821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:88 GQ:35.6 PL:[177.5, 0.0, 35.6] SR:48 DR:34 LR:-182.8 LO:182.8);ALT=G[chr2:37428783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37428869	+	chr2	37431447	+	.	0	12	754448_1	17.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=754448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_37411501_37436501_173C;SPAN=2578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:80 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:12 DR:0 LR:-17.94 LO:25.53);ALT=T[chr2:37431447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37456181	+	chr2	37458555	+	.	0	14	754608_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=754608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_37436001_37461001_249C;SPAN=2374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:103 GQ:18.5 PL:[18.5, 0.0, 229.7] SR:14 DR:0 LR:-18.31 LO:29.14);ALT=T[chr2:37458555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	37614007	-	chr2	37615746	+	.	8	0	755030_1	4.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=755030_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:37614007(-)-2:37615746(-)__2_37607501_37632501D;SPAN=1739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=[chr2:37615746[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	37873966	+	chr2	37898567	+	.	0	15	755669_1	37.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=755669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_37877001_37902001_49C;SPAN=24601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:45 GQ:37.4 PL:[37.4, 0.0, 70.4] SR:15 DR:0 LR:-37.32 LO:37.92);ALT=C[chr2:37898567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	38570658	+	chr2	38604283	+	.	9	4	757378_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTAG;MAPQ=60;MATEID=757378_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_38563001_38588001_249C;SPAN=33625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:38 GQ:22.7 PL:[22.7, 0.0, 68.9] SR:4 DR:9 LR:-22.72 LO:24.04);ALT=G[chr2:38604283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	38976895	+	chr2	38978440	+	.	13	0	758714_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=758714_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:38976895(+)-2:38978440(-)__2_38955001_38980001D;SPAN=1545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:131 GQ:7.7 PL:[7.7, 0.0, 308.0] SR:0 DR:13 LR:-7.422 LO:25.16);ALT=G[chr2:38978440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	38977338	+	chr2	38978371	+	.	0	25	758717_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=758717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_38955001_38980001_20C;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:112 GQ:52.4 PL:[52.4, 0.0, 217.4] SR:25 DR:0 LR:-52.18 LO:58.02);ALT=T[chr2:38978371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39005453	+	chr2	39008658	+	.	9	0	758933_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=758933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:39005453(+)-2:39008658(-)__2_39004001_39029001D;SPAN=3205;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=T[chr2:39008658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39006260	+	chr2	39008659	+	.	0	10	758936_1	8.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=758936_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_39004001_39029001_41C;SPAN=2399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:91 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:10 DR:0 LR:-8.356 LO:19.82);ALT=A[chr2:39008659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39103251	+	chr2	39107740	+	CTTCAGAAGTGTATAAGATCAGCTTTATCTTTCCAAATGGAGACAAGTAT	0	7	759326_1	1.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTTCAGAAGTGTATAAGATCAGCTTTATCTTTCCAAATGGAGACAAGTAT;MAPQ=60;MATEID=759326_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_39102001_39127001_349C;SPAN=4489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:7 DR:0 LR:-0.8912 LO:13.07);ALT=A[chr2:39107740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39103251	+	chr2	39107320	+	.	3	6	759325_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=759325_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_2_39102001_39127001_349C;SPAN=4069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:6 DR:3 LR:1.055 LO:10.95);ALT=A[chr2:39107320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39664663	+	chr2	39680977	+	.	9	0	760931_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=760931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:39664663(+)-2:39680977(-)__2_39665501_39690501D;SPAN=16314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:0 DR:9 LR:-22.12 LO:22.58);ALT=G[chr2:39680977[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	39664680	+	chr2	39681434	+	.	12	0	760932_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=760932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:39664680(+)-2:39681434(-)__2_39665501_39690501D;SPAN=16754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:0 DR:12 LR:-30.67 LO:30.91);ALT=T[chr2:39681434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
