chr3	174858271	+	chr3	175028421	+	.	77	56	2501666_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=2501666_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_175028001_175053001_313C;SPAN=170150;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:32 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:56 DR:77 LR:-307.0 LO:307.0);ALT=C[chr3:175028421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	175158865	+	chr3	175225978	+	.	103	70	2502168_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=2502168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_175224001_175249001_100C;SPAN=67113;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:135 DP:54 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:70 DR:103 LR:-399.4 LO:399.4);ALT=T[chr3:175225978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
