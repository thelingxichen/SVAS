chr3	80062866	+	chr3	80065278	-	TA	10	28	2133324_1	96.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TA;MAPQ=60;MATEID=2133324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_80041501_80066501_176C;SPAN=2412;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:71 GQ:73.4 PL:[96.5, 0.0, 73.4] SR:28 DR:10 LR:-96.43 LO:96.43);ALT=A]chr3:80065278];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	80590176	+	chr9	12556845	+	.	5	21	5783260_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTC;MAPQ=60;MATEID=5783260_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_12544001_12569001_7C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:34 GQ:17.3 PL:[63.5, 0.0, 17.3] SR:21 DR:5 LR:-64.73 LO:64.73);ALT=C[chr9:12556845[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	108936730	+	chr3	80590920	+	.	15	12	8316828_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AAACAAACAAACAAACAAA;MAPQ=45;MATEID=8316828_2;MATENM=0;NM=2;NUMPARTS=3;REPSEQ=AACAAACAAACAAACA;SCTG=c_13_108927001_108952001_509C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:18 DP:110 GQ:3.2 PL:[0.0, 3.2, 86.9] SR:12 DR:15 LR:4.639 LO:5.802);ALT=]chr13:108936730]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	80925314	+	chr3	80926605	+	.	0	91	2137393_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TTT;MAPQ=60;MATEID=2137393_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_80923501_80948501_407C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:70 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:91 DR:0 LR:-267.4 LO:267.4);ALT=T[chr3:80926605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	12556849	+	chr9	12559647	+	.	61	33	5783286_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CAATACAATACTTTTC;MAPQ=60;MATEID=5783286_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_12544001_12569001_233C;SPAN=2798;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:58 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:33 DR:61 LR:-254.2 LO:254.2);ALT=C[chr9:12559647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
