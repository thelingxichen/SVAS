chr11	104267751	+	chr11	104273230	+	.	72	53	4986586_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATA;MAPQ=60;MATEID=4986586_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_104247501_104272501_21C;SPAN=5479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:11 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:53 DR:72 LR:-280.6 LO:280.6);ALT=A[chr11:104273230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104813701	+	chr11	104815474	+	.	0	23	4987765_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4987765_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_104811001_104836001_40C;SPAN=1773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:86 GQ:52.7 PL:[52.7, 0.0, 155.0] SR:23 DR:0 LR:-52.62 LO:55.48);ALT=C[chr11:104815474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104815580	+	chr11	104817807	+	.	0	44	4987775_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=4987775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_104811001_104836001_32C;SPAN=2227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:91 GQ:97.7 PL:[120.8, 0.0, 97.7] SR:44 DR:0 LR:-120.7 LO:120.7);ALT=T[chr11:104817807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104822734	+	chr11	104825474	+	.	0	8	4987797_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4987797_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_104811001_104836001_89C;SPAN=2740;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:8 DR:0 LR:-3.65 LO:15.33);ALT=T[chr11:104825474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104825714	+	chr11	104839244	+	.	45	0	4987821_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4987821_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:104825714(+)-11:104839244(-)__11_104835501_104860501D;SPAN=13530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:53 GQ:7.5 PL:[141.9, 7.5, 0.0] SR:0 DR:45 LR:-144.0 LO:144.0);ALT=T[chr11:104839244[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104897085	+	chr11	104899851	+	TGCGGAAAATTTCCTCCACATCACAGGAACAGGCATATTCTTGCATATGTTCAATGAGTCTTCCAATAAAAACAGAGCCCATTGTGGGATGTCTCCAAGAAACATTAT	6	32	4988286_1	96.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGCGGAAAATTTCCTCCACATCACAGGAACAGGCATATTCTTGCATATGTTCAATGAGTCTTCCAATAAAAACAGAGCCCATTGTGGGATGTCTCCAAGAAACATTAT;MAPQ=60;MATEID=4988286_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_104884501_104909501_141C;SPAN=2766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:83 GQ:96.5 PL:[96.5, 0.0, 103.1] SR:32 DR:6 LR:-96.35 LO:96.37);ALT=T[chr11:104899851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104897680	+	chr11	104899851	+	.	3	4	4988289_1	2.0	.	DISC_MAPQ=52;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4988289_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_11_104884501_104909501_141C;SPAN=2171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:4 DR:3 LR:-2.246 LO:13.27);ALT=T[chr11:104899851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104902010	+	chr11	104903791	+	.	0	8	4988295_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4988295_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_104884501_104909501_230C;SPAN=1781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:8 DR:0 LR:-5.818 LO:15.7);ALT=G[chr11:104903791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104912449	+	chr11	104914210	+	.	0	19	4987995_1	38.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4987995_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_104909001_104934001_202C;SPAN=1761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:92 GQ:38 PL:[38.0, 0.0, 183.2] SR:19 DR:0 LR:-37.79 LO:43.36);ALT=G[chr11:104914210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	104912450	+	chr11	104915119	+	.	4	34	4987996_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGC;MAPQ=60;MATEID=4987996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_104909001_104934001_256C;SPAN=2669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:98 GQ:89 PL:[89.0, 0.0, 148.4] SR:34 DR:4 LR:-88.99 LO:89.81);ALT=C[chr11:104915119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
