chr13	43443321	+	chr13	51747959	-	.	17	0	8033197_1	43.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=8033197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:43443321(+)-13:51747959(+)__13_43438501_43463501D;SPAN=8304638;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:48 GQ:43.1 PL:[43.1, 0.0, 72.8] SR:0 DR:17 LR:-43.11 LO:43.54);ALT=G]chr13:51747959];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	51069350	+	chr13	51075079	+	.	165	115	8065430_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCTC;MAPQ=60;MATEID=8065430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_51058001_51083001_200C;SPAN=5729;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:229 DP:42 GQ:61.9 PL:[679.9, 61.9, 0.0] SR:115 DR:165 LR:-680.0 LO:680.0);ALT=C[chr13:51075079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
