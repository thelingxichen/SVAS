chr4	151688777	-	chr4	151690129	+	.	8	0	2992889_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2992889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:151688777(-)-4:151690129(-)__4_151679501_151704501D;SPAN=1352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:122 GQ:6.3 PL:[0.0, 6.3, 306.9] SR:0 DR:8 LR:6.645 LO:13.98);ALT=[chr4:151690129[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	152219332	-	chr4	152220656	+	.	9	0	2995490_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=2995490_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:152219332(-)-4:152220656(-)__4_152218501_152243501D;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:124 GQ:3.6 PL:[0.0, 3.6, 306.9] SR:0 DR:9 LR:3.886 LO:16.14);ALT=[chr4:152220656[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	152990314	+	chr4	152993952	+	C	82	46	2998505_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=2998505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_152978001_153003001_320C;SPAN=3638;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:101 DP:93 GQ:27 PL:[297.0, 27.0, 0.0] SR:46 DR:82 LR:-297.1 LO:297.1);ALT=T[chr4:152993952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	153458637	+	chr4	153474507	+	.	51	42	3000274_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=3000274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_153468001_153493001_22C;SPAN=15870;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:35 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:42 DR:51 LR:-224.5 LO:224.5);ALT=T[chr4:153474507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	154074599	+	chr4	153875835	+	.	10	0	3002872_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3002872_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:153875835(-)-4:154074599(+)__4_154056001_154081001D;SPAN=198764;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.75 LO:21.78);ALT=]chr4:154074599]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	20255414	+	chr4	153979395	+	.	2	33	8370641_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=CTTCCTTCCTTCCTTCCTTCCTTCCTTC;MAPQ=60;MATEID=8370641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_20237001_20262001_347C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:34 DP:48 GQ:16.7 PL:[99.2, 0.0, 16.7] SR:33 DR:2 LR:-102.5 LO:102.5);ALT=]chr14:20255414]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	125191874	+	chr5	125485938	-	.	21	0	3735454_1	59.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=3735454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:125191874(+)-5:125485938(+)__5_125170501_125195501D;SPAN=294064;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:35 GQ:23.6 PL:[59.9, 0.0, 23.6] SR:0 DR:21 LR:-60.61 LO:60.61);ALT=A]chr5:125485938];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	125498526	+	chr5	125496416	+	.	63	0	3736437_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3736437_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:125496416(-)-5:125498526(+)__5_125489001_125514001D;SPAN=2110;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:141 GQ:99 PL:[170.0, 0.0, 170.0] SR:0 DR:63 LR:-169.8 LO:169.8);ALT=]chr5:125498526]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	125496712	+	chr5	125498729	+	.	31	0	3736440_1	65.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3736440_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:125496712(+)-5:125498729(-)__5_125489001_125514001D;SPAN=2017;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:135 GQ:65.9 PL:[65.9, 0.0, 260.6] SR:0 DR:31 LR:-65.76 LO:72.38);ALT=G[chr5:125498729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	126065136	+	chr14	20777471	+	G	6	35	8373677_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=8373677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_20776001_20801001_421C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:63 GQ:49.1 PL:[101.9, 0.0, 49.1] SR:35 DR:6 LR:-102.7 LO:102.7);ALT=C[chr14:20777471[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
