chr8	115788620	+	chr1	99679031	+	.	21	0	5635216_1	50.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=5635216_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:99679031(-)-8:115788620(+)__8_115787001_115812001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:69 GQ:50.6 PL:[50.6, 0.0, 116.6] SR:0 DR:21 LR:-50.63 LO:52.07);ALT=]chr8:115788620]T;VARTYPE=BND:TRX-th;JOINTYPE=th
