chr3	192875332	+	chr3	192885406	+	.	157	107	2576974_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TCT;MAPQ=60;MATEID=2576974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_192864001_192889001_269C;SPAN=10074;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:210 DP:38 GQ:56.8 PL:[623.8, 56.8, 0.0] SR:107 DR:157 LR:-623.9 LO:623.9);ALT=T[chr3:192885406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
