chr11	127533450	+	chr11	127534511	+	.	0	63	7269743_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7269743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_127522501_127547501_198C;SPAN=1061;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:139 GQ:99 PL:[170.3, 0.0, 167.0] SR:63 DR:0 LR:-170.3 LO:170.3);ALT=T[chr11:127534511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
