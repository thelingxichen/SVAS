chr5	103854288	+	chr5	103860327	+	.	49	23	2545031_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AATAAAATTATTAA;MAPQ=60;MATEID=2545031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_103855501_103880501_168C;SPAN=6039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:15 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:23 DR:49 LR:-171.6 LO:171.6);ALT=A[chr5:103860327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
