chr6	125597393	+	chr6	125613973	+	TGTGGAATCATAGAAGTCTTGCAGTCTCCCAGGTTTGTGTTCAAGGTCTTCATATTCAGATGCTTGAAGAATCATTTCACATTGGTCTAGCTGCTTCACAAATTTGGCTTCTGCACTAGATTGGGTCTCGTACT	0	20	3015921_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGTGGAATCATAGAAGTCTTGCAGTCTCCCAGGTTTGTGTTCAAGGTCTTCATATTCAGATGCTTGAAGAATCATTTCACATTGGTCTAGCTGCTTCACAAATTTGGCTTCTGCACTAGATTGGGTCTCGTACT;MAPQ=60;MATEID=3015921_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_125587001_125612001_7C;SPAN=16580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:34 GQ:23.9 PL:[56.9, 0.0, 23.9] SR:20 DR:0 LR:-57.44 LO:57.44);ALT=C[chr6:125613973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	125598387	+	chr6	125613973	+	.	2	8	3015951_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=3015951_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TATATA;SCTG=c_6_125611501_125636501_57C;SPAN=15586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:29 GQ:18.2 PL:[18.2, 0.0, 33.8] SR:8 DR:2 LR:-18.16 LO:18.48);ALT=C[chr6:125613973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	125614100	+	chr6	125623007	+	.	12	0	3015960_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3015960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:125614100(+)-6:125623007(-)__6_125611501_125636501D;SPAN=8907;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:0 DR:12 LR:-17.4 LO:25.39);ALT=C[chr6:125623007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	125620015	+	chr6	125623030	+	.	8	0	3015972_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3015972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:125620015(+)-6:125623030(-)__6_125611501_125636501D;SPAN=3015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=T[chr6:125623030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	125621807	+	chr6	125622995	+	.	41	14	3015977_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3015977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_125611501_125636501_117C;SPAN=1188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:84 GQ:79.7 PL:[122.6, 0.0, 79.7] SR:14 DR:41 LR:-122.9 LO:122.9);ALT=T[chr6:125622995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	125708765	+	chr6	125711353	+	.	51	36	3016421_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGCTATGTATATTTTA;MAPQ=60;MATEID=3016421_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_125709501_125734501_34C;SPAN=2588;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:22 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:36 DR:51 LR:-204.7 LO:204.7);ALT=A[chr6:125711353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	126240577	+	chr6	126242087	+	.	7	4	3017366_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3017366_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_126224001_126249001_210C;SPAN=1510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:4 DR:7 LR:-5.276 LO:15.61);ALT=G[chr6:126242087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	126240583	+	chr6	126243825	+	.	8	0	3017367_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3017367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:126240583(+)-6:126243825(-)__6_126224001_126249001D;SPAN=3242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:0 DR:8 LR:-4.192 LO:15.42);ALT=T[chr6:126243825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	126661547	+	chr6	126667350	+	.	0	23	3018448_1	64.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=3018448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_126640501_126665501_91C;SPAN=5803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:42 GQ:35 PL:[64.7, 0.0, 35.0] SR:23 DR:0 LR:-64.93 LO:64.93);ALT=T[chr6:126667350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	126667468	+	chr6	126669610	+	.	0	30	3018362_1	78.0	.	EVDNC=ASSMB;HOMSEQ=AGGTAA;MAPQ=60;MATEID=3018362_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_126665001_126690001_42C;SPAN=2142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:77 GQ:78.2 PL:[78.2, 0.0, 107.9] SR:30 DR:0 LR:-78.17 LO:78.44);ALT=A[chr6:126669610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	127637649	+	chr6	127651952	+	CTGGAGTTCCTAGTGATTTCACAGCATTCAGATCAGATCCTGAAGAGAAAGTATTTTTTGCCCCACGGACAATGAGGCCTTTCCCCTCTGTCCAATTTTCCAATTCAATTACTTTTTCCAGAAGTTGTAGCATCATAAC	2	21	3020336_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=CTGGAGTTCCTAGTGATTTCACAGCATTCAGATCAGATCCTGAAGAGAAAGTATTTTTTGCCCCACGGACAATGAGGCCTTTCCCCTCTGTCCAATTTTCCAATTCAATTACTTTTTCCAGAAGTTGTAGCATCATAAC;MAPQ=60;MATEID=3020336_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_127645001_127670001_38C;SPAN=14303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:37 GQ:26.3 PL:[62.6, 0.0, 26.3] SR:21 DR:2 LR:-63.36 LO:63.36);ALT=T[chr6:127651952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	127648337	+	chr6	127652006	+	.	13	0	3020339_1	18.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3020339_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:127648337(+)-6:127652006(-)__6_127645001_127670001D;SPAN=3669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=A[chr6:127652006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	127652176	+	chr6	127664481	+	.	4	11	3020344_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3020344_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_127645001_127670001_58C;SPAN=12305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:88 GQ:22.4 PL:[22.4, 0.0, 190.7] SR:11 DR:4 LR:-22.37 LO:30.18);ALT=C[chr6:127664481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
