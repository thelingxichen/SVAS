chr2	66505594	+	chr2	66507554	+	.	75	42	829012_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TATAT;MAPQ=60;MATEID=829012_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_66493001_66518001_235C;SPAN=1960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:50 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:42 DR:75 LR:-283.9 LO:283.9);ALT=T[chr2:66507554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	66663000	+	chr2	66664868	+	.	27	27	829863_1	99.0	.	DISC_MAPQ=20;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=829863_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_66640001_66665001_219C;SPAN=1868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:97 GQ:89.3 PL:[145.4, 0.0, 89.3] SR:27 DR:27 LR:-146.1 LO:146.1);ALT=G[chr2:66664868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
