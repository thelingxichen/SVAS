chr1	109876083	+	chr1	109035476	+	.	65	0	453344_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=453344_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109035476(-)-1:109876083(+)__1_109858001_109883001D;SPAN=840607;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:39 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=]chr1:109876083]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	155531857	+	chr1	110191216	+	.	21	0	2425703_1	61.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2425703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110191216(-)-3:155531857(+)__3_155526001_155551001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:29 GQ:8.6 PL:[61.4, 0.0, 8.6] SR:0 DR:21 LR:-63.72 LO:63.72);ALT=]chr3:155531857]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	223760191	+	chr2	223762672	+	.	124	71	1712352_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TACTTTGTTCTTT;MAPQ=60;MATEID=1712352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_223758501_223783501_374C;SPAN=2481;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:172 DP:31 GQ:46.3 PL:[508.3, 46.3, 0.0] SR:71 DR:124 LR:-508.3 LO:508.3);ALT=T[chr2:223762672[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	1069522	+	chr2	223906780	+	.	10	31	1712899_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TTCCTTCCTTCCTTCCTTCCTTCCT;MAPQ=28;MATEID=1712899_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_2_223905501_223930501_6C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:31 DR:10 LR:-115.5 LO:115.5);ALT=]chr3:1069522]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	224039700	+	chr9	109426677	+	.	42	37	1713500_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1713500_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_224028001_224053001_383C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:39 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:37 DR:42 LR:-184.8 LO:184.8);ALT=T[chr9:109426677[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	109426854	+	chr2	224039705	+	AAATTTTAAAATTTAAAATATAAAG	33	43	1713501_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAATTTTAAAATTTAAAATATAAAG;MAPQ=60;MATEID=1713501_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_224028001_224053001_249C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:60 DP:40 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:43 DR:33 LR:-178.2 LO:178.2);ALT=]chr9:109426854]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	224731130	-	chr2	224732162	+	.	6	2	1716634_1	0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AAGAAAGAA;MAPQ=60;MATEID=1716634_2;MATENM=0;NM=22;NUMPARTS=2;SCTG=c_2_224714001_224739001_294C;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:136 GQ:16.8 PL:[0.0, 16.8, 363.0] SR:2 DR:6 LR:17.04 LO:9.431);ALT=[chr2:224732162[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	92696684	+	chr2	225020292	+	.	102	63	11312443_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=11312443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_92683501_92708501_465C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:142 DP:76 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:63 DR:102 LR:-419.2 LO:419.2);ALT=]chrX:92696684]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	1200564	-	chr3	154949022	+	.	2	41	1798373_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=ATATATA;MAPQ=60;MATEID=1798373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_1200501_1225501_264C;SPAN=153748458;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:42 DP:30 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:41 DR:2 LR:-122.1 LO:122.1);ALT=[chr3:154949022[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	156054148	+	chr3	47248229	+	.	17	61	2427273_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAGTGAGACTCTGTA;MAPQ=60;MATEID=2427273_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_156040501_156065501_307C;SPAN=108805919;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:82 GQ:2.1 PL:[201.3, 2.1, 0.0] SR:61 DR:17 LR:-211.3 LO:211.3);ALT=]chr3:156054148]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	47490669	+	chr3	47493441	+	.	0	120	1994839_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GC;MAPQ=60;MATEID=1994839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47481001_47506001_276C;SPAN=2772;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:120 DP:44 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:120 DR:0 LR:-356.5 LO:356.5);ALT=C[chr3:47493441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101730109	+	chr3	155027219	+	.	25	48	2423134_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2423134_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_155011501_155036501_189C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:31 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:48 DR:25 LR:-208.0 LO:208.0);ALT=]chr8:101730109]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	101717282	+	chr4	39974878	+	.	12	0	5581249_1	20.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5581249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:39974878(-)-8:101717282(+)__8_101699501_101724501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:0 DR:12 LR:-20.92 LO:26.38);ALT=]chr8:101717282]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	112272693	-	chr7	113309202	+	.	53	40	5141632_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=5141632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_113288001_113313001_828C;SPAN=1036509;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:91 DP:170 GQ:99 PL:[254.3, 0.0, 158.6] SR:40 DR:53 LR:-255.5 LO:255.5);ALT=[chr7:113309202[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	113278356	-	chr7	113308981	+	.	115	58	5141634_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=5141634_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_113288001_113313001_786C;SPAN=30625;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:155 DP:109 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:58 DR:115 LR:-458.8 LO:458.8);ALT=[chr7:113308981[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	113304906	+	chr7	113310352	+	.	121	0	5141880_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5141880_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:113304906(+)-7:113310352(-)__7_113288001_113313001D;SPAN=5446;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:121 DP:175 GQ:71.6 PL:[352.1, 0.0, 71.6] SR:0 DR:121 LR:-362.4 LO:362.4);ALT=A[chr7:113310352[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	113309208	+	chr7	119449935	+	AGTGTTATTTATAATTT	39	23	5234034_1	65.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AGTGTTATTTATAATTT;MAPQ=60;MATEID=5234034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119437501_119462501_476C;SPAN=6140727;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:429 GQ:65.4 PL:[65.4, 0.0, 976.4] SR:23 DR:39 LR:-65.33 LO:113.0);ALT=A[chr7:119449935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	93794269	+	chr7	114156676	+	.	34	39	5155610_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5155610_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_114145501_114170501_5C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:72 DP:237 GQ:99 PL:[173.5, 0.0, 401.3] SR:39 DR:34 LR:-173.5 LO:178.5);ALT=]chrX:93794269]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	118511939	+	chr7	114553649	+	.	42	28	5162378_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;MAPQ=60;MATEID=5162378_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_114537501_114562501_458C;SPAN=3958290;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:232 GQ:99 PL:[142.0, 0.0, 419.3] SR:28 DR:42 LR:-141.8 LO:149.5);ALT=]chr7:118511939]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	73783717	+	chr7	115123696	+	.	39	27	5174231_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5174231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_115101001_115126001_8C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:58 DP:243 GQ:99 PL:[125.8, 0.0, 462.5] SR:27 DR:39 LR:-125.6 LO:136.5);ALT=]chr8:73783717]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	115420825	+	chr7	115419623	+	.	10	0	5180801_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5180801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:115419623(-)-7:115420825(+)__7_115419501_115444501D;SPAN=1202;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:569 GQ:99 PL:[0.0, 121.0, 1624.0] SR:0 DR:10 LR:121.1 LO:11.72);ALT=]chr7:115420825]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	115692348	-	chr7	118423829	+	GAATAGT	186	75	5216336_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GAATAGT;MAPQ=60;MATEID=5216336_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_118408501_118433501_804C;SPAN=2731481;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:236 DP:425 GQ:99 PL:[664.0, 0.0, 367.0] SR:75 DR:186 LR:-668.5 LO:668.5);ALT=[chr7:118423829[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	115957391	-	chr7	119974386	+	.	40	18	5247531_1	10.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5247531_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119952001_119977001_630C;SPAN=4016995;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:561 GQ:10.1 PL:[10.1, 0.0, 1350.0] SR:18 DR:40 LR:-9.76 LO:91.99);ALT=[chr7:119974386[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	115997416	+	chr7	118752504	+	.	46	7	5224681_1	48.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=5224681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118751501_118776501_1023C;SPAN=2755088;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:419 GQ:48.3 PL:[48.3, 0.0, 969.2] SR:7 DR:46 LR:-48.23 LO:98.55);ALT=T[chr7:118752504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	116476385	+	chr7	118784002	-	.	33	12	5225811_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=5225811_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_118776001_118801001_672C;SPAN=2307617;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:41 DP:548 GQ:12.9 PL:[0.0, 12.9, 1357.0] SR:12 DR:33 LR:13.13 LO:74.1);ALT=A]chr7:118784002];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	116905059	-	chr15	70823811	+	.	14	12	8964487_1	75.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGGGAGGGAGGGAGGGAGGGAGGGAAGGAAGGAA;MAPQ=50;MATEID=8964487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_70805001_70830001_110C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:26 DP:19 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:12 DR:14 LR:-75.92 LO:75.92);ALT=[chr15:70823811[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	116933097	+	chr7	116934197	-	.	6	2	5190396_1	0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CTCAAGTGATCCTC;MAPQ=60;MATEID=5190396_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_116914001_116939001_382C;SPAN=1100;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:968 GQ:99 PL:[0.0, 235.6, 2822.0] SR:2 DR:6 LR:235.8 LO:6.835);ALT=G]chr7:116934197];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	119135589	+	chr7	116972812	+	.	41	18	5189617_1	54.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=5189617_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_116963001_116988001_1182C;SPAN=2162777;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:48 DP:383 GQ:54.9 PL:[54.9, 0.0, 873.5] SR:18 DR:41 LR:-54.68 LO:98.08);ALT=]chr7:119135589]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	117121237	+	chr7	118488083	+	CGTTGTGT	36	18	5217509_1	10.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CGTTGTGT;MAPQ=60;MATEID=5217509_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118482001_118507001_184C;SPAN=1366846;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:42 DP:475 GQ:10.1 PL:[10.1, 0.0, 1142.0] SR:18 DR:36 LR:-9.953 LO:79.08);ALT=G[chr7:118488083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	117142799	+	chr7	120330482	+	.	70	25	5191579_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAAA;MAPQ=60;MATEID=5191579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_117134501_117159501_410C;SPAN=3187683;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:87 DP:285 GQ:99 PL:[210.1, 0.0, 480.8] SR:25 DR:70 LR:-210.0 LO:215.9);ALT=A[chr7:120330482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	117689710	+	chr7	121705300	-	.	116	38	5204853_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5204853_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_117673501_117698501_122C;SPAN=4015590;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:135 DP:274 GQ:99 PL:[371.6, 0.0, 292.3] SR:38 DR:116 LR:-371.9 LO:371.9);ALT=G]chr7:121705300];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	118121523	-	chr7	118981037	+	TAAAC	49	18	5229842_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TAAAC;MAPQ=60;MATEID=5229842_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_118972001_118997001_502C;SPAN=859514;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:60 DP:342 GQ:99 PL:[105.6, 0.0, 722.9] SR:18 DR:49 LR:-105.4 LO:132.2);ALT=[chr7:118981037[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	118443664	+	chr7	118170911	+	C	106	42	5216903_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=5216903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118433001_118458001_412C;SPAN=272753;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:128 DP:463 GQ:99 PL:[297.3, 0.0, 825.4] SR:42 DR:106 LR:-297.1 LO:310.9);ALT=]chr7:118443664]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	118176721	+	chr7	118444821	+	.	106	36	5216907_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTAC;MAPQ=60;MATEID=5216907_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118433001_118458001_346C;SPAN=268100;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:127 DP:410 GQ:99 PL:[308.2, 0.0, 687.7] SR:36 DR:106 LR:-308.2 LO:316.1);ALT=C[chr7:118444821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	118177975	-	chr7	118430105	+	.	111	49	5216339_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=5216339_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118408501_118433501_893C;SPAN=252130;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:146 DP:334 GQ:99 PL:[391.6, 0.0, 418.0] SR:49 DR:111 LR:-391.5 LO:391.5);ALT=[chr7:118430105[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	118726893	+	chr7	119450134	+	.	7	42	5234035_1	17.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTCCTC;MAPQ=60;MATEID=5234035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119437501_119462501_232C;SPAN=723241;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:49 DP:533 GQ:17.6 PL:[17.6, 0.0, 1275.0] SR:42 DR:7 LR:-17.35 LO:93.13);ALT=C[chr7:119450134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	118731607	+	chr7	119394262	-	.	106	52	5233426_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTC;MAPQ=60;MATEID=5233426_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119388501_119413501_902C;SPAN=662655;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:146 DP:517 GQ:99 PL:[342.0, 0.0, 913.0] SR:52 DR:106 LR:-341.9 LO:356.3);ALT=A]chr7:119394262];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	118776423	-	chr7	118793834	+	.	39	43	5225823_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5225823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118776001_118801001_700C;SPAN=17411;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:82 DP:894 GQ:28.8 PL:[28.8, 0.0, 2141.0] SR:43 DR:39 LR:-28.48 LO:155.8);ALT=[chr7:118793834[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	118831248	+	chr7	118834755	+	CAAATAAGTGA	218	114	5225441_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CAAATAAGTGA;MAPQ=60;MATEID=5225441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118825001_118850001_770C;SPAN=3507;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:338 DP:238 GQ:91.4 PL:[1003.0, 91.4, 0.0] SR:114 DR:218 LR:-1003.0 LO:1003.0);ALT=T[chr7:118834755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	118851011	+	chr7	119000648	+	.	39	20	5227095_1	59.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=5227095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_118849501_118874501_257C;SPAN=149637;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:404 GQ:59.1 PL:[59.1, 0.0, 920.6] SR:20 DR:39 LR:-58.9 LO:104.4);ALT=A[chr7:119000648[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	119003138	+	chr7	119004403	-	.	21	0	5230569_1	0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=5230569_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:119003138(+)-7:119004403(+)__7_118996501_119021501D;SPAN=1265;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:21 DP:766 GQ:99 PL:[0.0, 137.9, 2136.0] SR:0 DR:21 LR:138.2 LO:28.64);ALT=C]chr7:119004403];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	93798174	+	chr7	119100295	+	.	45	63	5232959_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=5232959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119094501_119119501_1051C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:128 DP:472 GQ:99 PL:[294.9, 0.0, 849.4] SR:63 DR:45 LR:-294.7 LO:309.7);ALT=]chrX:93798174]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chrX	93798218	+	chr7	119100546	+	.	12	0	5232965_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5232965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:119100546(-)-23:93798218(+)__7_119094501_119119501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:12 DP:492 GQ:93.3 PL:[0.0, 93.3, 1380.0] SR:0 DR:12 LR:93.68 LO:15.76);ALT=]chrX:93798218]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	119709219	-	chr7	121689822	+	.	38	17	5241469_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=5241469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119707001_119732001_144C;SPAN=1980603;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:50 DP:742 GQ:35.6 PL:[0.0, 35.6, 1872.0] SR:17 DR:38 LR:35.98 LO:88.01);ALT=[chr7:121689822[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	119853025	+	chr7	120317208	+	.	23	8	5245703_1	0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=5245703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_119829501_119854501_718C;SPAN=464183;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:29 DP:505 GQ:40.8 PL:[0.0, 40.8, 1307.0] SR:8 DR:23 LR:41.09 LO:48.97);ALT=A[chr7:120317208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	120034884	+	chr7	120521380	+	.	19	14	5249472_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5249472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_120025501_120050501_867C;SPAN=486496;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:37 DP:651 GQ:53.8 PL:[0.0, 53.8, 1687.0] SR:14 DR:19 LR:54.24 LO:62.31);ALT=C[chr7:120521380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	120454918	+	chr7	120125628	+	.	43	15	5250527_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5250527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_120123501_120148501_290C;SPAN=329290;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:572 GQ:10.4 PL:[10.4, 0.0, 1377.0] SR:15 DR:43 LR:-10.08 LO:93.88);ALT=]chr7:120454918]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	120604730	-	chrX	92560525	+	.	102	46	11310524_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=11310524_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_92536501_92561501_112C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:132 DP:103 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:46 DR:102 LR:-389.5 LO:389.5);ALT=[chrX:92560525[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	122106295	+	chr7	122104868	+	.	29	0	5267380_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5267380_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:122104868(-)-7:122106295(+)__7_122083501_122108501D;SPAN=1427;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:29 DP:1016 GQ:99 PL:[0.0, 179.2, 2825.0] SR:0 DR:29 LR:179.5 LO:40.06);ALT=]chr7:122106295]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	122675155	-	chr7	122676417	+	.	9	0	5266541_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5266541_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:122675155(-)-7:122676417(-)__7_122671501_122696501D;SPAN=1262;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:133 GQ:6 PL:[0.0, 6.0, 333.3] SR:0 DR:9 LR:6.324 LO:15.86);ALT=[chr7:122676417[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	101730011	-	chr13	25670814	+	.	7	37	7958869_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGAATGCTCCTAAATG;MAPQ=40;MATEID=7958869_2;MATENM=43;NM=4;NUMPARTS=2;SCTG=c_13_25651501_25676501_53C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:43 DP:78 GQ:68 PL:[120.8, 0.0, 68.0] SR:37 DR:7 LR:-121.6 LO:121.6);ALT=[chr13:25670814[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	110033444	+	chr9	110035449	+	A	50	31	5956671_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=5956671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_110029501_110054501_130C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:56 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:31 DR:50 LR:-201.3 LO:201.3);ALT=T[chr9:110035449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110537535	+	chr9	110540596	+	.	83	38	5957710_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TAAAAATATTTTGTA;MAPQ=60;MATEID=5957710_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_110519501_110544501_72C;SPAN=3061;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:16 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:38 DR:83 LR:-303.7 LO:303.7);ALT=A[chr9:110540596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	71594663	+	chr15	71597706	+	.	105	50	8967760_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=8967760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_71589001_71614001_102C;SPAN=3043;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:127 DP:107 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:50 DR:105 LR:-376.3 LO:376.3);ALT=A[chr15:71597706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72385978	+	chr15	72388159	+	.	132	102	8971959_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GCCTGTAATCCCA;MAPQ=60;MATEID=8971959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72373001_72398001_8C;SPAN=2181;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:207 DP:66 GQ:55.9 PL:[613.9, 55.9, 0.0] SR:102 DR:132 LR:-614.0 LO:614.0);ALT=A[chr15:72388159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	90409454	+	chrX	93186830	+	.	46	0	11316141_1	99.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=11316141_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:90409454(+)-23:93186830(-)__23_93173501_93198501D;SPAN=2777376;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:46 DP:141 GQ:99 PL:[113.9, 0.0, 226.1] SR:0 DR:46 LR:-113.6 LO:115.8);ALT=A[chrX:93186830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	92621882	+	chrX	92696965	+	.	127	54	11312499_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTTT;MAPQ=60;MATEID=11312499_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_92683501_92708501_621C;SPAN=75083;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:160 DP:116 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:54 DR:127 LR:-475.3 LO:475.3);ALT=T[chrX:92696965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	92740536	+	chrX	93275162	-	.	118	58	11314551_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=11314551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_93271501_93296501_342C;SPAN=534626;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:162 DP:136 GQ:43.6 PL:[478.6, 43.6, 0.0] SR:58 DR:118 LR:-478.6 LO:478.6);ALT=T]chrX:93275162];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	92796299	+	chrX	92801505	+	.	138	106	11311788_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAT;MAPQ=60;MATEID=11311788_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_92781501_92806501_371C;SPAN=5206;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:192 DP:107 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:106 DR:138 LR:-567.7 LO:567.7);ALT=T[chrX:92801505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	93486122	+	chrX	93453708	+	.	73	25	11317020_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ATG;MAPQ=60;MATEID=11317020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_93467501_93492501_131C;SPAN=32414;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:89 DP:117 GQ:21.2 PL:[262.1, 0.0, 21.2] SR:25 DR:73 LR:-274.1 LO:274.1);ALT=]chrX:93486122]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	93604956	-	chrX	93780434	+	.	70	38	11318738_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=11318738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_93761501_93786501_55C;SPAN=175478;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:91 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:38 DR:70 LR:-303.7 LO:303.7);ALT=[chrX:93780434[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
