chr5	174130029	+	chr5	174131988	+	.	59	0	3943170_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=3943170_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:174130029(+)-5:174131988(-)__5_174121501_174146501D;SPAN=1959;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:59 DP:106 GQ:90.2 PL:[166.1, 0.0, 90.2] SR:0 DR:59 LR:-167.2 LO:167.2);ALT=A[chr5:174131988[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
