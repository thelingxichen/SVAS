chr12	118941242	+	chr13	100082612	+	.	18	40	7856640_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TATCCAT;MAPQ=60;MATEID=7856640_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_118923001_118948001_204C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:102 GQ:99 PL:[117.8, 0.0, 127.7] SR:40 DR:18 LR:-117.6 LO:117.6);ALT=T[chr13:100082612[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	99254189	+	chr13	99257489	-	.	21	29	8263750_1	88.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GCAGTGAG;MAPQ=9;MATEID=8263750_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_99249501_99274501_521C;SPAN=3300;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:41 DP:173 GQ:88.7 PL:[88.7, 0.0, 329.6] SR:29 DR:21 LR:-88.47 LO:96.37);ALT=C]chr13:99257489];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	99257406	-	chr13	99258525	+	TATA	15	53	8263771_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;INSERTION=TATA;MAPQ=38;MATEID=8263771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_99249501_99274501_309C;SPAN=1119;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:111 GQ:92.3 PL:[174.8, 0.0, 92.3] SR:53 DR:15 LR:-175.9 LO:175.9);ALT=[chr13:99258525[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
