chr5	106484529	+	chr5	94409552	-	.	20	25	5563801_1	99.0	.	BX=CATCTTAGTGAGGGTT-1_1,TGAAAGACAACTCATG-1_1,TCGCGTTCAATTAAGG-1_1,GCATCTCGTACGTCGC-1_1,GTTCATTAGAAAGCTT-1_1,TTAGGCAAGTCCGGTC-1_1,ACACTCCCACATGCGC-1_3,GCTGAATAGGTGTAGC-1_1,TAGCGTAGTGCTCGAC-1_2,AATCGTGTCCACTGCT-1_1,TCAATCTCATATGTGC-1_1,TCTCATAAGAGTATGT-1_1,GACTTGACACGTGCGT-1_1,AAGACAACAGGAAGAA-1_1,AACAAGATCAAAGCGG-1_1,TGTGGTAGTCCTCCAT-1_1,CTCGGTTTCGGCGCAT-1_1,TTGTCCGTCTCCACAC-1_1,CCATGGGGTTACCAGT-1_1,CCTCCCTCATAACAAG-1_1,AACGATCGTATGTGTC-1_1,TACCTTAAGTGTGATA-1_1,TCGCGGATCCAAGTAC-1_1,TCTGCCACACGAGCTC-1_1,GTTTAGGGTCGATTGT-1_1,TGCGCAGTCGCTGACG-1_1,AGAGCTTCAATGGGAC-1_1,CAGGAGAGTCGTAGCC-1_1,CATGCCTCAACATAGA-1_1,AGGCGAATCTCTGCTG-1_1,CAACCAATCTACACCC-1_1;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5563801_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_106477001_106502001_8C;SPAN=12074977;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:20 GQ:5.4 PL:[0.0, 5.4, 59.4] SR:0 DR:0 LR:5.619 LO:0.0),OC001T.bam(GT:1/1 AD:37 DP:36 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:25 DR:20 LR:-112.2 LO:112.2);ALT=c]chr5:106484529];VARTYPE=BND:INV-tt;JOINTYPE=tt	.
chr5	94411322	-	chr5	106482726	+	.	47	39	5563802_1	99.0	.	BX=CCTAAAGCATCGTTAG-1_1,TACGGGCAGATGCGAC-1_1,GACCAATCATGTTGCA-1_1,CGTCCATCACGAAAGC-1_1,GCAGCCATCCCTTCGA-1_2,ACGCTAAAGGACTTAA-1_1,TTGTCCGTCGAATGCT-1_1,CGCTATCTCATGTGGT-1_1,CCTTCCCAGGAAACAG-1_1,AGGGAGTGTTATCGGT-1_1,AGCGCCAGTTAAAGAC-1_3,CATATTCCACACCGAC-1_1,TATCTACGTTCAAGGG-1_4,GGGAGATCAGGTGAAC-1_1,CAAGCGCAGTAGTATG-1_1,TTTACTGGTGTTCAAC-1_1,TATCAGGGTTTAAGCC-1_1,AGGGAACTCGACCCTT-1_1,GACACGCTCCGAACGC-1_1,AGATGGGTCTAATGGC-1_2,ATACGCAAGATTCAAG-1_1,GGACATTAGTTAGGGC-1_1,TACTTGTGTGTTGTTG-1_1,GCGCAACTCGAATGCT-1_2,AGCATTGCACTTAAGC-1_3,TCTCACGTCTGCACTC-1_1,GGAAGCAGTGTTAAGA-1_1,TAGCAGTGTGAACCTT-1_2,CACGTAACATCGATGT-1_1,CCTAAAGGTCCGCAGT-1_3,GCCAAATCATGGGAAC-1_1,GTTCATTAGTGCGATG-1_2,CAAAGCTTCTGGCCGA-1_1,ATCACTTCATTCCGTC-1_1,TTGGCTCTCGTAGATC-1_3,GCCTATCTCATCTTTG-1_1,ACCCAGGCATCGGGCT-1_1,GTTGAACCAAACAACA-1_1,TTAGGCAGTACCAACT-1_2,CATTACTGTACAACGG-1_1,ACGATCAAGCGACCAA-1_1,TGCGCGATCCGTCTAC-1_1;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAG;MAPQ=60;MATEID=5563802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_106477001_106502001_367C;SPAN=12071404;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:17 GQ:4.5 PL:[0.0, 4.5, 49.5] SR:0 DR:0 LR:4.776 LO:0.0),OC001T.bam(GT:1/1 AD:66 DP:36 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:47 LR:-201.3 LO:201.3);ALT=[chr5:106482726[T;VARTYPE=BND:INV-hh;JOINTYPE=hh	.
chr5	94411322	-	chr5	106482726	+	.	47	39	5563802_1	99.0	.	BX=CCTAAAGCATCGTTAG-1_1,TACGGGCAGATGCGAC-1_1,GACCAATCATGTTGCA-1_1,CGTCCATCACGAAAGC-1_1,GCAGCCATCCCTTCGA-1_2,ACGCTAAAGGACTTAA-1_1,TTGTCCGTCGAATGCT-1_1,CGCTATCTCATGTGGT-1_1,CCTTCCCAGGAAACAG-1_1,AGGGAGTGTTATCGGT-1_1,AGCGCCAGTTAAAGAC-1_3,CATATTCCACACCGAC-1_1,TATCTACGTTCAAGGG-1_4,GGGAGATCAGGTGAAC-1_1,CAAGCGCAGTAGTATG-1_1,TTTACTGGTGTTCAAC-1_1,TATCAGGGTTTAAGCC-1_1,AGGGAACTCGACCCTT-1_1,GACACGCTCCGAACGC-1_1,AGATGGGTCTAATGGC-1_2,ATACGCAAGATTCAAG-1_1,GGACATTAGTTAGGGC-1_1,TACTTGTGTGTTGTTG-1_1,GCGCAACTCGAATGCT-1_2,AGCATTGCACTTAAGC-1_3,TCTCACGTCTGCACTC-1_1,GGAAGCAGTGTTAAGA-1_1,TAGCAGTGTGAACCTT-1_2,CACGTAACATCGATGT-1_1,CCTAAAGGTCCGCAGT-1_3,GCCAAATCATGGGAAC-1_1,GTTCATTAGTGCGATG-1_2,CAAAGCTTCTGGCCGA-1_1,ATCACTTCATTCCGTC-1_1,TTGGCTCTCGTAGATC-1_3,GCCTATCTCATCTTTG-1_1,ACCCAGGCATCGGGCT-1_1,GTTGAACCAAACAACA-1_1,TTAGGCAGTACCAACT-1_2,CATTACTGTACAACGG-1_1,ACGATCAAGCGACCAA-1_1,TGCGCGATCCGTCTAC-1_1;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAG;MAPQ=60;MATEID=5563802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_106477001_106502001_367C;SPAN=12071404;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:17 GQ:4.5 PL:[0.0, 4.5, 49.5] SR:0 DR:0 LR:4.776 LO:0.0),OC001T.bam(GT:1/1 AD:66 DP:36 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:47 LR:-201.3 LO:201.3);ALT=[chr5:106482726[T;VARTYPE=BND:INV-hh;JOINTYPE=hh	.
chr5	106484529	+	chr5	94409552	-	.	20	25	5563801_1	99.0	.	BX=CATCTTAGTGAGGGTT-1_1,TGAAAGACAACTCATG-1_1,TCGCGTTCAATTAAGG-1_1,GCATCTCGTACGTCGC-1_1,GTTCATTAGAAAGCTT-1_1,TTAGGCAAGTCCGGTC-1_1,ACACTCCCACATGCGC-1_3,GCTGAATAGGTGTAGC-1_1,TAGCGTAGTGCTCGAC-1_2,AATCGTGTCCACTGCT-1_1,TCAATCTCATATGTGC-1_1,TCTCATAAGAGTATGT-1_1,GACTTGACACGTGCGT-1_1,AAGACAACAGGAAGAA-1_1,AACAAGATCAAAGCGG-1_1,TGTGGTAGTCCTCCAT-1_1,CTCGGTTTCGGCGCAT-1_1,TTGTCCGTCTCCACAC-1_1,CCATGGGGTTACCAGT-1_1,CCTCCCTCATAACAAG-1_1,AACGATCGTATGTGTC-1_1,TACCTTAAGTGTGATA-1_1,TCGCGGATCCAAGTAC-1_1,TCTGCCACACGAGCTC-1_1,GTTTAGGGTCGATTGT-1_1,TGCGCAGTCGCTGACG-1_1,AGAGCTTCAATGGGAC-1_1,CAGGAGAGTCGTAGCC-1_1,CATGCCTCAACATAGA-1_1,AGGCGAATCTCTGCTG-1_1,CAACCAATCTACACCC-1_1;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5563801_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_106477001_106502001_8C;SPAN=12074977;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:20 GQ:5.4 PL:[0.0, 5.4, 59.4] SR:0 DR:0 LR:5.619 LO:0.0),OC001T.bam(GT:1/1 AD:37 DP:36 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:25 DR:20 LR:-112.2 LO:112.2);ALT=c]chr5:106484529];VARTYPE=BND:INV-tt;JOINTYPE=tt	.
