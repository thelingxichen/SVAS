chrX	37639395	+	chrX	37641340	+	.	9	0	7400046_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7400046_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:37639395(+)-23:37641340(-)__23_37632001_37657001D;SPAN=1945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=A[chrX:37641340[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	37639404	+	chrX	37642741	+	.	22	0	7400047_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7400047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:37639404(+)-23:37642741(-)__23_37632001_37657001D;SPAN=3337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:56 GQ:57.5 PL:[57.5, 0.0, 77.3] SR:0 DR:22 LR:-57.45 LO:57.63);ALT=A[chrX:37642741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	37641436	+	chrX	37642742	+	.	0	22	7400049_1	53.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=7400049_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GGG;SCTG=c_23_37632001_37657001_101C;SPAN=1306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:69 GQ:53.9 PL:[53.9, 0.0, 113.3] SR:22 DR:0 LR:-53.93 LO:55.09);ALT=G[chrX:37642742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	37641436	+	chrX	37652917	+	TCAGCACTGGCACTGGCCAGGGCCCCTGCAGCCTGCCTGAATTTCAACTGCATGCTGATTCTCTTGCCAGTCTGTCGAAATCTGCTGTCCTTCCTCAGGGGTTCCAGTGCGTGCTGCTCAACAAGAGTTCGAAGACAACTGGACAGGAATCTCACCTTTCATAAAATGGTGGCATGGATGATTGCACTTCACTCT	0	26	7400050_1	68.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TCAGCACTGGCACTGGCCAGGGCCCCTGCAGCCTGCCTGAATTTCAACTGCATGCTGATTCTCTTGCCAGTCTGTCGAAATCTGCTGTCCTTCCTCAGGGGTTCCAGTGCGTGCTGCTCAACAAGAGTTCGAAGACAACTGGACAGGAATCTCACCTTTCATAAAATGGTGGCATGGATGATTGCACTTCACTCT;MAPQ=60;MATEID=7400050_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_37632001_37657001_101C;SPAN=11481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:65 GQ:68.3 PL:[68.3, 0.0, 88.1] SR:26 DR:0 LR:-68.22 LO:68.38);ALT=G[chrX:37652917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	37664421	+	chrX	37665638	+	.	3	2	7400024_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7400024_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_37656501_37681501_180C;SPAN=1217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:58 GQ:2.4 PL:[0.0, 2.4, 145.2] SR:2 DR:3 LR:2.51 LO:7.082);ALT=G[chrX:37665638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	37701182	+	chrX	37706731	+	.	8	0	7400210_1	19.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7400210_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:37701182(+)-23:37706731(-)__23_37705501_37730501D;SPAN=5549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:0 DR:8 LR:-19.36 LO:19.88);ALT=A[chrX:37706731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
