chr3	140544408	+	chr3	140547043	+	.	0	117	2364309_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCACT;MAPQ=60;MATEID=2364309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_140532001_140557001_145C;SPAN=2635;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:46 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:117 DR:0 LR:-346.6 LO:346.6);ALT=T[chr3:140547043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
