chr16	17830105	+	chr16	18003312	+	.	26	0	9187896_1	85.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=9187896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:17830105(+)-16:18003312(-)__16_17983001_18008001D;SPAN=173207;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:26 DP:29 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:26 LR:-85.54 LO:85.54);ALT=A[chr16:18003312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18832544	+	chr16	18838377	+	.	88	77	9194040_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GAGATATTTAGTATGTTTCT;MAPQ=60;MATEID=9194040_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_16_18816001_18841001_133C;SPAN=5833;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:141 DP:41 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:77 DR:88 LR:-415.9 LO:415.9);ALT=T[chr16:18838377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	19449758	-	chr22	46045011	+	.	8	41	9197974_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=AGAAAGAAAGAAAGAAAGAAAGAAA;MAPQ=60;MATEID=9197974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_19428501_19453501_256C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:41 DR:8 LR:-138.6 LO:138.6);ALT=[chr22:46045011[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr22	45687732	+	chr22	45686343	+	.	11	0	10905135_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10905135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:45686343(-)-22:45687732(+)__22_45668001_45693001D;SPAN=1389;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:135 GQ:0 PL:[0.0, 0.0, 326.7] SR:0 DR:11 LR:0.2638 LO:20.3);ALT=]chr22:45687732]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	45746447	+	chr22	45745440	+	.	40	6	10905246_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTCCTGACCTTGTGATCTGCCTGCCTCGGCCTCCCATAGTGCTGGGATTACAGGCGTGAGCCACCG;MAPQ=60;MATEID=10905246_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_22_45741501_45766501_188C;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:63 GQ:19.4 PL:[131.6, 0.0, 19.4] SR:6 DR:40 LR:-136.0 LO:136.0);ALT=]chr22:45746447]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	46014091	+	chr22	47986745	-	.	29	0	10910562_1	85.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=10910562_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:46014091(+)-22:47986745(+)__22_47971001_47996001D;SPAN=1972654;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:29 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=A]chr22:47986745];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr22	46964004	+	chr22	46962499	+	.	29	0	10907815_1	74.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=10907815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:46962499(-)-22:46964004(+)__22_46942001_46967001D;SPAN=1505;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:81 GQ:74 PL:[74.0, 0.0, 120.2] SR:0 DR:29 LR:-73.78 LO:74.45);ALT=]chr22:46964004]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	47231680	+	chr22	46968633	+	CAA	55	45	10909353_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CAA;MAPQ=60;MATEID=10909353_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_47211501_47236501_206C;SPAN=263047;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:46 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:45 DR:55 LR:-237.7 LO:237.7);ALT=]chr22:47231680]C;VARTYPE=BND:DUP-th;JOINTYPE=th
