chr3	32046583	+	chr3	31824042	+	.	78	0	1927331_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1927331_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:31824042(-)-3:32046583(+)__3_32021501_32046501D;SPAN=222541;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:6 GQ:21 PL:[231.0, 21.0, 0.0] SR:0 DR:78 LR:-231.1 LO:231.1);ALT=]chr3:32046583]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	32046937	+	chr3	31824043	+	.	81	43	1927467_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGACT;MAPQ=60;MATEID=1927467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32046001_32071001_421C;SPAN=222894;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:81 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:43 DR:81 LR:-323.5 LO:323.5);ALT=]chr3:32046937]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	32102052	+	chr3	32107884	+	.	179	120	1928273_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1928273_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_32095001_32120001_270C;SPAN=5832;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:240 DP:47 GQ:64.9 PL:[712.9, 64.9, 0.0] SR:120 DR:179 LR:-713.0 LO:713.0);ALT=C[chr3:32107884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32806763	+	chr3	32808062	+	.	62	17	1931521_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=TTGCAGTGAGCCAAGAT;MAPQ=44;MATEID=1931521_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32805501_32830501_381C;SPAN=1299;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:70 DP:98 GQ:32.9 PL:[204.5, 0.0, 32.9] SR:17 DR:62 LR:-211.6 LO:211.6);ALT=T[chr3:32808062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
