chr3	90377321	-	chr3	90380426	+	ACAAGAAGATGA	32	35	2171919_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCACAGG;INSERTION=ACAAGAAGATGA;MAPQ=60;MATEID=2171919_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CACA;SCTG=c_3_90380501_90405501_3C;SPAN=3105;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:12 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:35 DR:32 LR:-194.7 LO:194.7);ALT=[chr3:90380426[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	90421075	-	chr3	90423187	+	.	11	0	2171575_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2171575_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:90421075(-)-3:90423187(-)__3_90405001_90430001D;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:162 GQ:7.3 PL:[0.0, 7.3, 405.9] SR:0 DR:11 LR:7.579 LO:19.4);ALT=[chr3:90423187[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
