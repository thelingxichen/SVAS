chr7	149305824	+	chr7	149282148	+	.	19	0	5322395_1	55.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=5322395_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:149282148(-)-7:149305824(+)__7_149303001_149328001D;SPAN=23676;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:26 GQ:6.2 PL:[55.7, 0.0, 6.2] SR:0 DR:19 LR:-57.8 LO:57.8);ALT=]chr7:149305824]G;VARTYPE=BND:DUP-th;JOINTYPE=th
