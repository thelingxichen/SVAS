chr2	20233042	+	chr2	20234078	+	.	5	5	709046_1	7.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=709046_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_20212501_20237501_148C;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:5 DR:5 LR:-7.222 LO:17.79);ALT=T[chr2:20234078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	20234823	+	chr2	20237077	+	.	2	7	709065_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=709065_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_20237001_20262001_47C;SPAN=2254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:7 DR:2 LR:-16.93 LO:18.66);ALT=G[chr2:20237077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	20240773	+	chr2	20251168	+	.	0	38	709084_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TACC;MAPQ=60;MATEID=709084_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_20237001_20262001_99C;SPAN=10395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:94 GQ:99 PL:[100.1, 0.0, 126.5] SR:38 DR:0 LR:-99.97 LO:100.2);ALT=C[chr2:20251168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	20840941	+	chr2	20845098	+	.	0	8	710692_1	6.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=710692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_20825001_20850001_31C;SPAN=4157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:8 DR:0 LR:-6.36 LO:15.8);ALT=C[chr2:20845098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	20845248	+	chr2	20850788	+	.	8	0	710719_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=710719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:20845248(+)-2:20850788(-)__2_20849501_20874501D;SPAN=5540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=T[chr2:20850788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	21348353	+	chr2	21347270	+	.	18	0	711769_1	32.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=711769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:21347270(-)-2:21348353(+)__2_21339501_21364501D;SPAN=1083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:0 DR:18 LR:-32.87 LO:40.05);ALT=]chr2:21348353]C;VARTYPE=BND:DUP-th;JOINTYPE=th
