chr6	96387601	+	chr6	96389422	+	AA	62	62	4329224_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=AA;MAPQ=60;MATEID=4329224_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_96383001_96408001_16C;SPAN=1821;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:21 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:62 DR:62 LR:-300.4 LO:300.4);ALT=G[chr6:96389422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
