chr6	56758355	+	chr6	56760945	+	.	106	0	2864590_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=2864590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:56758355(+)-6:56760945(-)__6_56742001_56767001D;SPAN=2590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:323 GQ:99 PL:[262.6, 0.0, 520.1] SR:0 DR:106 LR:-262.4 LO:267.1);ALT=T[chr6:56760945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	57183397	+	chr6	57185255	+	.	0	9	2866143_1	4.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2866143_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_57183001_57208001_181C;SPAN=1858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:9 DR:0 LR:-3.971 LO:17.23);ALT=T[chr6:57185255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	57284911	+	chr6	57289366	+	TTACAGCTTCG	93	62	2866607_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TTACAGCTTCG;MAPQ=60;MATEID=2866607_2;MATENM=0;NM=40;NUMPARTS=2;SCTG=c_6_57281001_57306001_65C;SPAN=4455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:127 DP:163 GQ:18.7 PL:[375.2, 0.0, 18.7] SR:62 DR:93 LR:-394.1 LO:394.1);ALT=T[chr6:57289366[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	57746319	-	chr6	58353250	+	.	2	2	2870174_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTGACCAAAT;MAPQ=38;MATEID=2870174_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_58334501_58359501_281C;SPAN=606931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:59 GQ:2.7 PL:[0.0, 2.7, 148.5] SR:2 DR:2 LR:2.781 LO:7.052);ALT=[chr6:58353250[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
