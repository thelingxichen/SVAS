chr2	33224462	+	chr2	33227293	+	.	68	51	956849_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=956849_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_33222001_33247001_44C;SPAN=2831;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:101 DP:19 GQ:27 PL:[297.0, 27.0, 0.0] SR:51 DR:68 LR:-297.1 LO:297.1);ALT=A[chr2:33227293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
