chr2	127630610	+	chr2	127490057	+	.	79	15	1324598_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ATTG;MAPQ=60;MATEID=1324598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_127620501_127645501_424C;SPAN=140553;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:69 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:15 DR:79 LR:-241.0 LO:241.0);ALT=]chr2:127630610]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	127674758	+	chr2	127677273	+	.	131	107	1324378_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=1324378_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_127669501_127694501_130C;SPAN=2515;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:188 DP:34 GQ:50.8 PL:[557.8, 50.8, 0.0] SR:107 DR:131 LR:-557.8 LO:557.8);ALT=C[chr2:127677273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
