chr16	62544333	+	chr16	62550669	+	AAGGT	134	41	9360644_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AAGGT;MAPQ=60;MATEID=9360644_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_62548501_62573501_174C;SPAN=6336;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:144 DP:17 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:41 DR:134 LR:-425.8 LO:425.8);ALT=A[chr16:62550669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	63362844	+	chr16	63350361	+	.	0	62	9363841_1	99.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=9363841_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_63332501_63357501_232C;SPAN=12483;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:62 DP:74 GQ:6.6 PL:[191.4, 6.6, 0.0] SR:62 DR:0 LR:-197.4 LO:197.4);ALT=]chr16:63362844]A;VARTYPE=BND:DUP-th;JOINTYPE=th
