chr7	29860045	+	chr7	29519649	+	.	6	4	4661075_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=4661075_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_29841001_29866001_408C;SPAN=340396;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:160 GQ:16.9 PL:[0.0, 16.9, 422.5] SR:4 DR:6 LR:16.94 LO:13.02);ALT=]chr7:29860045]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	29881662	+	chr7	29682913	+	.	50	23	4661293_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4661293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_29865501_29890501_62C;SPAN=198749;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:59 DP:113 GQ:99 PL:[164.3, 0.0, 108.2] SR:23 DR:50 LR:-164.7 LO:164.7);ALT=]chr7:29881662]C;VARTYPE=BND:DUP-th;JOINTYPE=th
