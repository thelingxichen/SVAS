chr18	76494764	-	chr18	76498681	+	.	12	0	10092132_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10092132_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:76494764(-)-18:76498681(-)__18_76489001_76514001D;SPAN=3917;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:12 DP:595 GQ:99 PL:[0.0, 121.3, 1687.0] SR:0 DR:12 LR:121.6 LO:14.77);ALT=[chr18:76498681[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	76728685	+	chr22	50933872	+	.	15	0	10917142_1	46.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=10917142_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:76728685(+)-22:50933872(-)__22_50911001_50936001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:18 GQ:1.5 PL:[46.2, 1.5, 0.0] SR:0 DR:15 LR:-47.65 LO:47.65);ALT=G[chr22:50933872[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr18	76797689	+	chr18	76796622	+	.	4	2	10094733_1	0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=TCCACCCAGGCATCCTGG;MAPQ=0;MATEID=10094733_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_18_76783001_76808001_196C;SECONDARY;SPAN=1067;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:161 GQ:26.8 PL:[0.0, 26.8, 442.3] SR:2 DR:4 LR:27.11 LO:7.09);ALT=]chr18:76797689]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	51119772	+	chr22	51117945	+	.	40	0	10917405_1	99.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=10917405_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:51117945(-)-22:51119772(+)__22_51107001_51132001D;SPAN=1827;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:0 DR:40 LR:-109.9 LO:109.9);ALT=]chr22:51119772]G;VARTYPE=BND:DUP-th;JOINTYPE=th
