chr20	10394581	+	chr20	10401172	+	.	0	29	6918972_1	69.0	.	EVDNC=ASSMB;HOMSEQ=TTACCT;MAPQ=60;MATEID=6918972_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_10388001_10413001_29C;SPAN=6591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:96 GQ:69.8 PL:[69.8, 0.0, 162.2] SR:29 DR:0 LR:-69.72 LO:71.79);ALT=T[chr20:10401172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	10401432	+	chr20	10414752	+	.	56	0	6919042_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6919042_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:10401432(+)-20:10414752(-)__20_10412501_10437501D;SPAN=13320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:55 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:56 LR:-165.0 LO:165.0);ALT=A[chr20:10414752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	11281584	-	chrX	81651235	+	TTTAATACT	19	28	6921816_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTTAATACT;MAPQ=60;MATEID=6921816_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_20_11270001_11295001_404C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:30 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:28 DR:19 LR:-112.2 LO:112.2);ALT=[chrX:81651235[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr20	11647434	+	chr20	11648671	+	.	41	35	6922888_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTCA;MAPQ=60;MATEID=6922888_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_20_11637501_11662501_342C;SPAN=1237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:67 GQ:18 PL:[198.0, 18.0, 0.0] SR:35 DR:41 LR:-198.0 LO:198.0);ALT=A[chr20:11648671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	80457705	+	chrX	80533828	+	.	11	0	7459595_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7459595_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:80457705(+)-23:80533828(-)__23_80433501_80458501D;SPAN=76123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:0 DR:11 LR:-18.43 LO:23.96);ALT=G[chrX:80533828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	80532669	+	chrX	80533829	+	.	4	46	7459697_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=7459697_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GGGG;SCTG=c_23_80531501_80556501_238C;SPAN=1160;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:81 GQ:60.8 PL:[133.4, 0.0, 60.8] SR:46 DR:4 LR:-134.5 LO:134.5);ALT=G[chrX:80533829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	80533911	+	chrX	80552692	+	.	3	17	7459704_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=7459704_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_23_80531501_80556501_238C;SPAN=18781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:64 GQ:48.8 PL:[48.8, 0.0, 104.9] SR:17 DR:3 LR:-48.68 LO:49.87);ALT=G[chrX:80552692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	81096653	+	chrX	81102693	+	.	49	35	7460460_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGGCAATTTGG;MAPQ=60;MATEID=7460460_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_23_81095001_81120001_102C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:25 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:35 DR:49 LR:-194.7 LO:194.7);ALT=G[chrX:81102693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
