chr5	97401563	+	chr5	97402761	+	.	0	51	3629386_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=3629386_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_97387501_97412501_54C;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:51 DP:102 GQ:99 PL:[140.9, 0.0, 104.6] SR:51 DR:0 LR:-141.0 LO:141.0);ALT=G[chr5:97402761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	97509883	+	chr5	97511060	-	.	8	0	3630002_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3630002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:97509883(+)-5:97511060(+)__5_97510001_97535001D;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:0 DR:8 LR:-8.798 LO:16.28);ALT=C]chr5:97511060];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	14394624	+	chr5	97869171	+	TGATGGGGTTGTTTGTTTTTTCTTGTAAATGTGT	4	134	9525557_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=TGATGGGGTTGTTTGTTTTTTCTTGTAAATGTGT;MAPQ=60;MATEID=9525557_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_17_14381501_14406501_229C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:138 DP:51 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:134 DR:4 LR:-409.3 LO:409.3);ALT=]chr17:14394624]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	97869240	+	chr17	14394623	+	GTTTAGGTTAAAGCATACATATCTTATCCATTAATTTAGGTGTTTTATGTTTCCTGTAGTTATTGTTATTGGAATGTTTTTTCTTAAACATTTTCTGAAAAGTTAATGATGCATAGAAAAATTTTTGCTTGTTGATATATCAATCTACTTTACTGAACCCTTATACTGGTCTAATAGTTTTTGGCTGAATCTCTTAAATGTGCTAGATAGATAATATTACCATTTGAAAATATTGTGAGTGTTTTCTCCTTTTTTCTTCAATATTTTAGATCTCTGTTTTTTCTTCTCAATGCATTGAC	2	132	9525558_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=GTTTAGGTTAAAGCATACATATCTTATCCATTAATTTAGGTGTTTTATGTTTCCTGTAGTTATTGTTATTGGAATGTTTTTTCTTAAACATTTTCTGAAAAGTTAATGATGCATAGAAAAATTTTTGCTTGTTGATATATCAATCTACTTTACTGAACCCTTATACTGGTCTAATAGTTTTTGGCTGAATCTCTTAAATGTGCTAGATAGATAATATTACCATTTGAAAATATTGTGAGTGTTTTCTCCTTTTTTCTTCAATATTTTAGATCTCTGTTTTTTCTTCTCAATGCATTGAC;MAPQ=60;MATEID=9525558_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_17_14381501_14406501_229C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:133 DP:49 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:132 DR:2 LR:-392.8 LO:392.8);ALT=T[chr17:14394623[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	98345117	+	chr5	98347483	+	AC	0	79	3633224_1	99.0	.	EVDNC=ASSMB;INSERTION=AC;MAPQ=60;MATEID=3633224_2;MATENM=1;NM=5;NUMPARTS=2;SCTG=c_5_98343001_98368001_226C;SPAN=2366;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:34 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:79 DR:0 LR:-234.4 LO:234.4);ALT=C[chr5:98347483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	14189911	+	chr17	14191556	+	.	131	84	9524211_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=9524211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_14185501_14210501_77C;SPAN=1645;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:179 DP:32 GQ:48.4 PL:[531.4, 48.4, 0.0] SR:84 DR:131 LR:-531.4 LO:531.4);ALT=A[chr17:14191556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	14746283	-	chr17	14747765	+	.	8	0	9526635_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=9526635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:14746283(-)-17:14747765(-)__17_14724501_14749501D;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:120 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.103 LO:14.04);ALT=[chr17:14747765[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	15595508	-	chr17	18593411	+	.	5	24	9531299_1	74.0	.	DISC_MAPQ=15;EVDNC=ASDIS;HOMSEQ=TCATAAAAAACAGTTTCAGTAAGAAATTACAAATTTTCTT;MAPQ=46;MATEID=9531299_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_15582001_15607001_14C;SPAN=2997903;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:77 GQ:74.9 PL:[74.9, 0.0, 111.2] SR:24 DR:5 LR:-74.87 LO:75.27);ALT=[chr17:18593411[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	18286842	+	chr17	74017600	-	.	9	0	9545879_1	8.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=9545879_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:18286842(+)-17:74017600(+)__17_18277001_18302001D;SPAN=55730758;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-7.764 LO:17.89);ALT=T]chr17:74017600];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	73985741	-	chr17	73986988	+	.	8	0	9816276_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9816276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73985741(-)-17:73986988(-)__17_73965501_73990501D;SPAN=1247;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:142 GQ:11.7 PL:[0.0, 11.7, 366.3] SR:0 DR:8 LR:12.06 LO:13.44);ALT=[chr17:73986988[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
