chr16	20571933	+	chr16	20475592	+	.	0	10	9202764_1	13.0	.	EVDNC=ASSMB;HOMSEQ=TCAGGTAT;MAPQ=57;MATEID=9202764_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_20457501_20482501_323C;SPAN=96341;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:10 DR:0 LR:-13.5 LO:20.92);ALT=]chr16:20571933]T;VARTYPE=BND:DUP-th;JOINTYPE=th
