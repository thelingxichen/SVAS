chr2	170641518	+	chr2	170643952	+	.	103	80	1497538_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=TCATTATTTTC;MAPQ=0;MATEID=1497538_2;MATENM=6;NM=1;NUMPARTS=2;SCTG=c_2_170618001_170643001_339C;SPAN=2434;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:149 DP:27 GQ:40.3 PL:[442.3, 40.3, 0.0] SR:80 DR:103 LR:-442.3 LO:442.3);ALT=C[chr2:170643952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	171510865	+	chr2	171512056	-	.	8	0	1500844_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1500844_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:171510865(+)-2:171512056(+)__2_171500001_171525001D;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:143 GQ:12 PL:[0.0, 12.0, 369.6] SR:0 DR:8 LR:12.33 LO:13.42);ALT=A]chr2:171512056];VARTYPE=BND:INV-hh;JOINTYPE=hh
