chr5	127407443	+	chr5	127410917	+	.	67	59	3744323_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=3744323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_127400001_127425001_104C;SPAN=3474;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:98 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:59 DR:67 LR:-307.0 LO:307.0);ALT=G[chr5:127410917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
