chr10	53651436	+	chr10	53761867	+	.	62	50	6268614_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=6268614_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_53630501_53655501_147C;SPAN=110431;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:42 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:50 DR:62 LR:-267.4 LO:267.4);ALT=T[chr10:53761867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
