chr8	121437607	+	chr8	121444270	+	.	0	18	4048668_1	35.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4048668_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_121422001_121447001_25C;SPAN=6663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:87 GQ:35.9 PL:[35.9, 0.0, 174.5] SR:18 DR:0 LR:-35.85 LO:41.09);ALT=C[chr8:121444270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	121444363	+	chr8	121455423	+	.	0	22	4048745_1	58.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=4048745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_121446501_121471501_15C;SPAN=11060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:54 GQ:58.1 PL:[58.1, 0.0, 71.3] SR:22 DR:0 LR:-57.99 LO:58.09);ALT=C[chr8:121455423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	121444411	+	chr8	121457307	+	.	24	0	4048746_1	66.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4048746_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:121444411(+)-8:121457307(-)__8_121446501_121471501D;SPAN=12896;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:48 GQ:49.7 PL:[66.2, 0.0, 49.7] SR:0 DR:24 LR:-66.34 LO:66.34);ALT=A[chr8:121457307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	121455563	+	chr8	121457307	+	.	18	0	4048760_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4048760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:121455563(+)-8:121457307(-)__8_121446501_121471501D;SPAN=1744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:95 GQ:33.8 PL:[33.8, 0.0, 195.5] SR:0 DR:18 LR:-33.68 LO:40.32);ALT=A[chr8:121457307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	121551209	+	chr8	121554050	+	.	3	2	4048981_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4048981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_121544501_121569501_109C;SPAN=2841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:87 GQ:6.9 PL:[0.0, 6.9, 224.4] SR:2 DR:3 LR:7.065 LO:8.445);ALT=G[chr8:121554050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
