chr2	242506103	+	chr2	242507335	+	ATT	133	95	1790602_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=ATT;MAPQ=27;MATEID=1790602_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_242501001_242526001_249C;SPAN=1232;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:203 DP:34 GQ:54.7 PL:[600.7, 54.7, 0.0] SR:95 DR:133 LR:-600.7 LO:600.7);ALT=A[chr2:242507335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	242854838	+	chr2	242867435	+	CTGCAATACCTGC	61	62	1791927_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTGCAATACCTGC;MAPQ=60;MATEID=1791927_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_242844001_242869001_67C;SPAN=12597;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:101 DP:87 GQ:27 PL:[297.0, 27.0, 0.0] SR:62 DR:61 LR:-297.1 LO:297.1);ALT=C[chr2:242867435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
