chr2	48576644	-	chr2	48578157	+	.	10	0	988634_1	13.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=988634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:48576644(-)-2:48578157(-)__2_48559001_48584001D;SPAN=1513;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:0 DR:10 LR:-12.96 LO:20.79);ALT=[chr2:48578157[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
