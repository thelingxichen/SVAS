chr1	105255033	+	chr1	105256189	+	.	59	34	441726_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=441726_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_1_105252001_105277001_15C;SPAN=1156;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:14 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:34 DR:59 LR:-247.6 LO:247.6);ALT=C[chr1:105256189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
