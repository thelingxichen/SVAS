chr6	129319530	+	chr6	129325575	+	.	52	36	3024000_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGAAGTATGATGACA;MAPQ=60;MATEID=3024000_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_129311001_129336001_59C;SPAN=6045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:72 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:36 DR:52 LR:-211.3 LO:211.3);ALT=A[chr6:129325575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	129963165	+	chr6	130031169	+	.	12	8	3025238_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3025238_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_130021501_130046501_109C;SPAN=68004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:36 GQ:39.8 PL:[39.8, 0.0, 46.4] SR:8 DR:12 LR:-39.76 LO:39.8);ALT=T[chr6:130031169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
