chr9	21007163	+	chr9	21011587	+	.	8	0	4152192_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4152192_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:21007163(+)-9:21011587(-)__9_20996501_21021501D;SPAN=4424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=T[chr9:21011587[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21008147	+	chr9	21011588	+	.	12	15	4152196_1	64.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4152196_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_20996501_21021501_147C;SPAN=3441;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:67 GQ:64.4 PL:[64.4, 0.0, 97.4] SR:15 DR:12 LR:-64.37 LO:64.76);ALT=T[chr9:21011588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21008147	+	chr9	21015894	+	TCAGCAAGAACACACAAAGGATAAATTGGCATCCATAGTGTTTGACTGAGCCATGTCAAGACAGCATAGGATATTCCTATGACTGATAACATGCTATAAGTG	6	27	4152197_1	85.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TACCT;INSERTION=TCAGCAAGAACACACAAAGGATAAATTGGCATCCATAGTGTTTGACTGAGCCATGTCAAGACAGCATAGGATATTCCTATGACTGATAACATGCTATAAGTG;MAPQ=60;MATEID=4152197_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_20996501_21021501_147C;SPAN=7747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:63 GQ:65.6 PL:[85.4, 0.0, 65.6] SR:27 DR:6 LR:-85.37 LO:85.37);ALT=T[chr9:21015894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21011696	+	chr9	21015894	+	.	2	8	4152200_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TACCT;MAPQ=60;MATEID=4152200_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_20996501_21021501_147C;SPAN=4198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:8 DR:2 LR:-14.27 LO:19.37);ALT=T[chr9:21015894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21016011	+	chr9	21029294	+	GCAAAAACCTTGGGAGAAGATGGTTTGACTCAATGCCAACATATATGTGCAGCAGTTCCAGGAGAGATACGGATTGGCAAAGTCGCATCACAAGTCCAATAGCATAAAAAGTGTCAACCATTGAAT	4	122	4152376_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GCAAAAACCTTGGGAGAAGATGGTTTGACTCAATGCCAACATATATGTGCAGCAGTTCCAGGAGAGATACGGATTGGCAAAGTCGCATCACAAGTCCAATAGCATAAAAAGTGTCAACCATTGAAT;MAPQ=60;MATEID=4152376_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_21021001_21046001_7C;SPAN=13283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:44 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:122 DR:4 LR:-366.4 LO:366.4);ALT=T[chr9:21029294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21016011	+	chr9	21026595	+	.	0	35	4152375_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4152375_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_21021001_21046001_7C;SPAN=10584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:40 GQ:7.5 PL:[112.2, 7.5, 0.0] SR:35 DR:0 LR:-113.5 LO:113.5);ALT=T[chr9:21026595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21016056	+	chr9	21031550	+	.	8	0	4152209_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4152209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:21016056(+)-9:21031550(-)__9_20996501_21021501D;SPAN=15494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:22 GQ:20.6 PL:[20.6, 0.0, 30.5] SR:0 DR:8 LR:-20.45 LO:20.61);ALT=A[chr9:21031550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21026724	+	chr9	21029294	+	.	2	81	4152386_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4152386_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_9_21021001_21046001_7C;SPAN=2570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:87 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:81 DR:2 LR:-257.5 LO:257.5);ALT=T[chr9:21029294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21026773	+	chr9	21031548	+	.	105	0	4152387_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4152387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:21026773(+)-9:21031548(-)__9_21021001_21046001D;SPAN=4775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:44 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:0 DR:105 LR:-310.3 LO:310.3);ALT=T[chr9:21031548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21029455	+	chr9	21031557	+	.	46	0	4152391_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4152391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:21029455(+)-9:21031557(-)__9_21021001_21046001D;SPAN=2102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:49 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:46 LR:-145.2 LO:145.2);ALT=G[chr9:21031557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21968244	+	chr9	21970901	+	.	4	13	4153719_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4153719_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_21952001_21977001_193C;SPAN=2657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:78 GQ:31.7 PL:[31.7, 0.0, 157.1] SR:13 DR:4 LR:-31.68 LO:36.46);ALT=G[chr9:21970901[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21971154	+	chr9	21994542	+	.	8	0	4153723_1	13.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=4153723_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:21971154(+)-9:21994542(-)__9_21952001_21977001D;SPAN=23388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=C[chr9:21994542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	21971210	+	chr9	21994136	+	.	0	23	4153725_1	65.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=4153725_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_21952001_21977001_194C;SPAN=22926;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:39 GQ:29 PL:[65.3, 0.0, 29.0] SR:23 DR:0 LR:-66.1 LO:66.1);ALT=G[chr9:21994136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	104204434	+	chr9	22413928	+	.	0	29	4365703_1	92.0	.	EVDNC=ASSMB;HOMSEQ=GAAGAGGAAGAGGAA;MAPQ=60;MATEID=4365703_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_104198501_104223501_116C;SPAN=81790506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:34 GQ:5.7 PL:[92.4, 5.7, 0.0] SR:29 DR:0 LR:-93.0 LO:93.0);ALT=]chr9:104204434]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	22496527	+	chr9	22504345	+	T	41	40	4154205_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=4154205_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_22491001_22516001_131C;SPAN=7818;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:20 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:40 DR:41 LR:-194.7 LO:194.7);ALT=T[chr9:22504345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	104153135	+	chr9	104160783	+	.	13	6	4365341_1	16.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4365341_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_104149501_104174501_239C;SPAN=7648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:124 GQ:16.1 PL:[16.1, 0.0, 283.4] SR:6 DR:13 LR:-15.92 LO:30.4);ALT=G[chr9:104160783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
