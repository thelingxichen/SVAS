chr6	1842332	+	chr6	1786678	+	.	4	5	3984381_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3984381_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_1837501_1862501_252C;SPAN=55654;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:7 DP:71 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:5 DR:4 LR:-3.871 LO:13.53);ALT=]chr6:1842332]A;VARTYPE=BND:DUP-th;JOINTYPE=th
