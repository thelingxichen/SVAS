chr5	172430170	+	chr5	172438654	+	.	91	42	3935065_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=3935065_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_172406501_172431501_296C;SPAN=8484;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:119 DP:52 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:42 DR:91 LR:-353.2 LO:353.2);ALT=A[chr5:172438654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	172973014	+	chr5	172974751	+	.	64	46	3937371_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GGAG;MAPQ=60;MATEID=3937371_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_172970001_172995001_182C;SPAN=1737;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:95 GQ:12.3 PL:[254.1, 12.3, 0.0] SR:46 DR:64 LR:-259.7 LO:259.7);ALT=G[chr5:172974751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
