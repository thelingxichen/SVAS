chrX	7623882	+	chrX	7673883	+	.	57	39	7359430_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=7359430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_7668501_7693501_0C;SPAN=50001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:9 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:39 DR:57 LR:-217.9 LO:217.9);ALT=C[chrX:7673883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	7868859	+	chrX	7870030	+	.	0	13	7359632_1	26.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7359632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_7864501_7889501_199C;SPAN=1171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:62 GQ:26.3 PL:[26.3, 0.0, 122.0] SR:13 DR:0 LR:-26.12 LO:29.76);ALT=C[chrX:7870030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	7894174	+	chrX	7895327	+	.	8	2	7359739_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7359739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_7889001_7914001_48C;SPAN=1153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:2 DR:8 LR:-10.97 LO:16.77);ALT=C[chrX:7895327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
