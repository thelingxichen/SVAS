chr6	112408923	+	chr6	112418242	+	.	9	5	2987490_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2987490_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_112406001_112431001_241C;SPAN=9319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:5 DR:9 LR:-8.577 LO:18.05);ALT=G[chr6:112418242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
