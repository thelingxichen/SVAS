chr5	106019406	+	chr5	106239812	+	.	9	0	3663625_1	17.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=3663625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:106019406(+)-5:106239812(-)__5_106232001_106257001D;SPAN=220406;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=C[chr5:106239812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
