chr4	64513	+	chr4	67888	+	TGTTTTTTATTATAA	0	34	2607198_1	0	.	EVDNC=ASSMB;INSERTION=TGTTTTTTATTATAA;MAPQ=60;MATEID=2607198_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_49001_74001_895C;SPAN=3375;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:34 DP:624 GQ:56.5 PL:[0.0, 56.5, 1627.0] SR:34 DR:0 LR:56.82 LO:56.62);ALT=T[chr4:67888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	86017	+	chr4	367143	+	.	25	27	2605691_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTGGAGAGAAACCCTACAAATGTGAAAAATGTGGCAAAGC;MAPQ=60;MATEID=2605691_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_4_343001_368001_307C;SPAN=281126;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:50 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:27 DR:25 LR:-148.5 LO:148.5);ALT=C[chr4:367143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	752279	+	chr4	753747	+	.	33	32	2606627_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CTCTCCCGAG;MAPQ=60;MATEID=2606627_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_4_735001_760001_233C;SPAN=1468;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:25 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:32 DR:33 LR:-184.8 LO:184.8);ALT=G[chr4:753747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1088927	+	chr4	1090160	+	.	8	0	2607920_1	3.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2607920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1088927(+)-4:1090160(-)__4_1078001_1103001D;SPAN=1233;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:0 DR:8 LR:-3.379 LO:15.29);ALT=T[chr4:1090160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1651678	-	chr4	1653815	+	.	8	0	2609626_1	0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2609626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1651678(-)-4:1653815(-)__4_1641501_1666501D;SPAN=2137;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:180 GQ:22.3 PL:[0.0, 22.3, 481.9] SR:0 DR:8 LR:22.36 LO:12.6);ALT=[chr4:1653815[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
