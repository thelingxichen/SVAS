chr12	129230114	+	chr12	129233186	+	.	29	0	5390890_1	80.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5390890_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:129230114(+)-12:129233186(-)__12_129213001_129238001D;SPAN=3072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:57 GQ:57.2 PL:[80.3, 0.0, 57.2] SR:0 DR:29 LR:-80.48 LO:80.48);ALT=A[chr12:129233186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
