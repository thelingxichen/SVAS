chr16	50709834	+	chr16	50711308	+	.	0	10	6210277_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6210277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_50690501_50715501_181C;SPAN=1474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:10 DR:0 LR:-17.57 LO:22.03);ALT=T[chr16:50711308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	50711469	+	chr16	50715113	+	.	14	0	6210388_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6210388_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:50711469(+)-16:50715113(-)__16_50715001_50740001D;SPAN=3644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:27 GQ:25.7 PL:[38.9, 0.0, 25.7] SR:0 DR:14 LR:-39.02 LO:39.02);ALT=G[chr16:50715113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	50776150	+	chr16	50783481	+	.	13	0	6210448_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6210448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:50776150(+)-16:50783481(-)__16_50764001_50789001D;SPAN=7331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:46 GQ:30.5 PL:[30.5, 0.0, 80.0] SR:0 DR:13 LR:-30.45 LO:31.73);ALT=G[chr16:50783481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	50776752	+	chr16	50783483	+	.	2	3	6210450_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACAG;MAPQ=60;MATEID=6210450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_50764001_50789001_29C;SPAN=6731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:47 GQ:0.5 PL:[0.5, 0.0, 112.7] SR:3 DR:2 LR:-0.4706 LO:7.462);ALT=G[chr16:50783483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
