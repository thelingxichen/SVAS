chr5	158630670	+	chr5	158636236	+	.	8	0	2624870_1	11.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2624870_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:158630670(+)-5:158636236(-)__5_158613001_158638001D;SPAN=5566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=A[chr5:158636236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	158690400	+	chr5	158695873	+	.	9	0	2624884_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2624884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:158690400(+)-5:158695873(-)__5_158686501_158711501D;SPAN=5473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=C[chr5:158695873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	66982806	+	chr5	159349715	+	.	28	0	7439918_1	82.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7439918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:159349715(-)-23:66982806(+)__23_66958501_66983501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:27 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:0 DR:28 LR:-82.52 LO:82.52);ALT=]chrX:66982806]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	159436261	+	chr5	159437506	+	.	25	0	2626114_1	65.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2626114_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:159436261(+)-5:159437506(-)__5_159421501_159446501D;SPAN=1245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:62 GQ:65.9 PL:[65.9, 0.0, 82.4] SR:0 DR:25 LR:-65.73 LO:65.86);ALT=G[chr5:159437506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	159832142	+	chr5	159833475	+	.	0	9	2626807_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2626807_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_159813501_159838501_35C;SPAN=1333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:9 DR:0 LR:-12.1 LO:18.81);ALT=G[chr5:159833475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	159842348	+	chr5	159846028	+	.	13	0	2626834_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2626834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:159842348(+)-5:159846028(-)__5_159838001_159863001D;SPAN=3680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:73 GQ:23.3 PL:[23.3, 0.0, 152.0] SR:0 DR:13 LR:-23.14 LO:28.73);ALT=A[chr5:159846028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
