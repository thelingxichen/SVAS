chr1	21722529	-	chr1	21723634	+	.	9	0	114476_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=114476_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:21722529(-)-1:21723634(-)__1_21707001_21732001D;SPAN=1105;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:140 GQ:8.1 PL:[0.0, 8.1, 356.4] SR:0 DR:9 LR:8.221 LO:15.65);ALT=[chr1:21723634[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
