chr15	52122033	+	chr15	52155006	+	.	57	38	5951038_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5951038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_52111501_52136501_92C;SPAN=32973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:38 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:38 DR:57 LR:-208.0 LO:208.0);ALT=G[chr15:52155006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	52155207	+	chr15	52161412	+	.	3	11	5951070_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5951070_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_52160501_52185501_202C;SPAN=6205;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:37 GQ:32.9 PL:[32.9, 0.0, 56.0] SR:11 DR:3 LR:-32.89 LO:33.24);ALT=G[chr15:52161412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	52311575	+	chr15	52338027	+	.	19	16	5951456_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=5951456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_52307501_52332501_138C;SPAN=26452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:7 GQ:9 PL:[99.0, 9.0, 0.0] SR:16 DR:19 LR:-99.02 LO:99.02);ALT=T[chr15:52338027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	52446273	+	chr15	52471965	+	.	0	10	5951811_1	24.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5951811_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_52454501_52479501_284C;SPAN=25692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:30 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:10 DR:0 LR:-24.88 LO:25.28);ALT=A[chr15:52471965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
