chr4	12715773	+	chr13	34803277	+	ATG	4	16	7997949_1	59.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=ATG;MAPQ=53;MATEID=7997949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_34790001_34815001_265C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:20 DP:10 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:16 DR:4 LR:-59.41 LO:59.41);ALT=A[chr13:34803277[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	34135730	+	chr13	34144822	+	.	76	53	7995288_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=7995288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_34128501_34153501_129C;SPAN=9092;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:95 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:53 DR:76 LR:-287.2 LO:287.2);ALT=T[chr13:34144822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
