chr5	61602364	+	chr5	61642956	+	.	8	5	2484535_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2484535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_61593001_61618001_176C;SPAN=40592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:24 GQ:26.6 PL:[29.9, 0.0, 26.6] SR:5 DR:8 LR:-29.81 LO:29.81);ALT=G[chr5:61642956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	61602395	+	chr5	61643872	+	.	13	0	2484536_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2484536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:61602395(+)-5:61643872(-)__5_61593001_61618001D;SPAN=41477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:26 GQ:26 PL:[35.9, 0.0, 26.0] SR:0 DR:13 LR:-35.93 LO:35.93);ALT=T[chr5:61643872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	61643051	+	chr5	61648413	+	ATTGACCTGGAGAGCATCTTTTCACTTAACCCTGACCTTGTTCCTGATGAAGAAATTGAACCCAGTCCAGAAACACCTCCACCTCCAGCATCCTCAGCCAAAGTAAACAAAATTGTAAAGAATCGACGGACTGTAGCTTCTATTAAGAATGACCCTCCTTCAAGAGATAATAG	0	26	2484426_1	70.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATTGACCTGGAGAGCATCTTTTCACTTAACCCTGACCTTGTTCCTGATGAAGAAATTGAACCCAGTCCAGAAACACCTCCACCTCCAGCATCCTCAGCCAAAGTAAACAAAATTGTAAAGAATCGACGGACTGTAGCTTCTATTAAGAATGACCCTCCTTCAAGAGATAATAG;MAPQ=60;MATEID=2484426_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_61642001_61667001_241C;SPAN=5362;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:57 GQ:67.1 PL:[70.4, 0.0, 67.1] SR:26 DR:0 LR:-70.39 LO:70.39);ALT=G[chr5:61648413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
