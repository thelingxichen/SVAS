chr1	61060479	+	chr1	61062109	+	TTTTATAGGAGCCT	0	11	172902_1	14.0	.	EVDNC=ASSMB;INSERTION=TTTTATAGGAGCCT;MAPQ=60;MATEID=172902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_61054001_61079001_176C;SPAN=1630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:82 GQ:14.3 PL:[14.3, 0.0, 182.6] SR:11 DR:0 LR:-14.1 LO:22.83);ALT=T[chr1:61062109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	61062660	+	chr1	61060495	+	CCA	20	20	172903_1	87.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCA;MAPQ=60;MATEID=172903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_61054001_61079001_327C;SPAN=2165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:78 GQ:87.8 PL:[87.8, 0.0, 101.0] SR:20 DR:20 LR:-87.8 LO:87.86);ALT=]chr1:61062660]C;VARTYPE=BND:DUP-th;JOINTYPE=th
