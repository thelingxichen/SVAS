chr9	19116649	+	chr9	19118319	+	.	2	2	4149321_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4149321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_19110001_19135001_273C;SPAN=1670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:59 GQ:2.7 PL:[0.0, 2.7, 148.5] SR:2 DR:2 LR:2.781 LO:7.052);ALT=T[chr9:19118319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	19121166	+	chr9	19126112	+	AGTTGATGGCTGATTCAGAATAGGCAGTCTCTCCTCAATCCTGTCTAGCCCCTTACAGGCATAGGTATTGGCAACTGCAA	0	32	4149331_1	90.0	.	EVDNC=ASSMB;INSERTION=AGTTGATGGCTGATTCAGAATAGGCAGTCTCTCCTCAATCCTGTCTAGCCCCTTACAGGCATAGGTATTGGCAACTGCAA;MAPQ=60;MATEID=4149331_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_19110001_19135001_143C;SPAN=4946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:56 GQ:44.3 PL:[90.5, 0.0, 44.3] SR:32 DR:0 LR:-91.26 LO:91.26);ALT=G[chr9:19126112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	19126308	+	chr9	19127417	+	GGTTGTGGATCAACTGCAACGGATGCCATTTTTCTTCCTGGAGAAAGAAAT	61	21	4149345_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGTTGTGGATCAACTGCAACGGATGCCATTTTTCTTCCTGGAGAAAGAAAT;MAPQ=60;MATEID=4149345_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_19110001_19135001_53C;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:58 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:21 DR:61 LR:-208.0 LO:208.0);ALT=C[chr9:19127417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
