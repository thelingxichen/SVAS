chr4	71878019	-	chr4	71955678	+	.	14	6	2749835_1	59.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=AGGAGGCCTGCCTGCCTCTGTAGACTCCACCTCTGGGGGCAGGGCATAGCCGAACAAAAGGCA;MAPQ=60;MATEID=2749835_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_4_71932001_71957001_1C;SPAN=77659;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:20 DP:8 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:6 DR:14 LR:-59.41 LO:59.41);ALT=[chr4:71955678[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	71878175	+	chr4	71955601	-	.	12	29	2749454_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=GAGATCTGAGAACGGACA;MAPQ=19;MATEID=2749454_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_4_71858501_71883501_172C;SPAN=77426;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:53 GQ:22.1 PL:[104.6, 0.0, 22.1] SR:29 DR:12 LR:-107.3 LO:107.3);ALT=A]chr4:71955601];VARTYPE=BND:INV-hh;JOINTYPE=hh
