chr20	39657740	+	chr20	39690033	+	ATCGAAGCGGATTTCCGATTGAAT	0	30	7012314_1	81.0	.	EVDNC=ASSMB;INSERTION=ATCGAAGCGGATTTCCGATTGAAT;MAPQ=60;MATEID=7012314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_39690001_39715001_233C;SPAN=32293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:64 GQ:71.9 PL:[81.8, 0.0, 71.9] SR:30 DR:0 LR:-81.71 LO:81.71);ALT=G[chr20:39690033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	39690130	+	chr20	39704807	+	.	0	8	7012315_1	0	.	EVDNC=ASSMB;HOMSEQ=ACAG;MAPQ=60;MATEID=7012315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_39690001_39715001_186C;SPAN=14677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:8 DR:0 LR:5.561 LO:14.1);ALT=G[chr20:39704807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	39704936	+	chr20	39706220	+	.	2	12	7012374_1	12.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=7012374_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_39690001_39715001_253C;SPAN=1284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:99 GQ:12.8 PL:[12.8, 0.0, 227.3] SR:12 DR:2 LR:-12.79 LO:24.33);ALT=T[chr20:39706220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	39704936	+	chr20	39708722	+	TCGAGCCTCTGGGGATGCAAAAATAAAGAAGGAGAAGGAAAATGGCTTCTC	2	15	7012375_1	23.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TAG;INSERTION=TCGAGCCTCTGGGGATGCAAAAATAAAGAAGGAGAAGGAAAATGGCTTCTC;MAPQ=60;MATEID=7012375_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_39690001_39715001_253C;SPAN=3786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:96 GQ:23.6 PL:[23.6, 0.0, 208.4] SR:15 DR:2 LR:-23.51 LO:32.21);ALT=T[chr20:39708722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	40126868	+	chr20	40127932	+	.	0	4	7013696_1	0	.	EVDNC=ASSMB;HOMSEQ=AACCT;MAPQ=60;MATEID=7013696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_40106501_40131501_158C;SPAN=1064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:113 GQ:17.1 PL:[0.0, 17.1, 306.9] SR:4 DR:0 LR:17.41 LO:5.901);ALT=T[chr20:40127932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	40162248	+	chr20	40246978	+	.	9	0	7014075_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7014075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:40162248(+)-20:40246978(-)__20_40229001_40254001D;SPAN=84730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=T[chr20:40246978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	40559921	+	chr20	40561561	-	.	10	0	7015132_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7015132_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:40559921(+)-20:40561561(+)__20_40547501_40572501D;SPAN=1640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:102 GQ:5.6 PL:[5.6, 0.0, 239.9] SR:0 DR:10 LR:-5.376 LO:19.3);ALT=C]chr20:40561561];VARTYPE=BND:INV-hh;JOINTYPE=hh
