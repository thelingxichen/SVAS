chr8	128806981	+	chr8	128902835	+	.	7	7	4070696_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4070696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_128894501_128919501_311C;SPAN=95854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:35 GQ:30.2 PL:[30.2, 0.0, 53.3] SR:7 DR:7 LR:-30.13 LO:30.52);ALT=G[chr8:128902835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	129465168	+	chr8	129471267	+	.	56	24	4072858_1	0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAGCTTGTGTTTTT;MAPQ=60;MATEID=4072858_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_129458001_129483001_91C;SPAN=6099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:66 DP:1454 GQ:99 PL:[0.0, 175.6, 3882.0] SR:24 DR:56 LR:176.1 LO:104.6);ALT=T[chr8:129471267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
