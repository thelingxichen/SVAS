chr17	11948606	-	chr17	13091777	+	.	64	47	9519830_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=9519830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_13083001_13108001_23C;SPAN=1143171;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:99 DP:42 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:47 DR:64 LR:-293.8 LO:293.8);ALT=[chr17:13091777[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	11948774	+	chr17	11983182	-	.	73	18	9517484_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=9517484_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_11980501_12005501_11C;SPAN=34408;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:33 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:18 DR:73 LR:-244.3 LO:244.3);ALT=C]chr17:11983182];VARTYPE=BND:INV-hh;JOINTYPE=hh
