chr6	84569512	+	chr6	84573891	+	.	12	0	2924034_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2924034_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:84569512(+)-6:84573891(-)__6_84574001_84599001D;SPAN=4379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:0 GQ:3 PL:[33.0, 3.0, 0.0] SR:0 DR:12 LR:-33.01 LO:33.01);ALT=T[chr6:84573891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	84569579	+	chr6	84603239	+	CCTTTAAAACAGGGCAGAAGCCTTATGGATTGGATTCGACTGACCAAAAGTGGAAAGGATCTAACGGGATTAAAAGGCAGGTTAATTGAAGTAACTGAAGAAGAACTTAAGAAACACAACAAAAAAGATGATTGTTGGATATGCATAAG	3	23	2924023_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=CCTTTAAAACAGGGCAGAAGCCTTATGGATTGGATTCGACTGACCAAAAGTGGAAAGGATCTAACGGGATTAAAAGGCAGGTTAATTGAAGTAACTGAAGAAGAACTTAAGAAACACAACAAAAAAGATGATTGTTGGATATGCATAAG;MAPQ=60;MATEID=2924023_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_84549501_84574501_111C;SPAN=33660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:57 GQ:60.5 PL:[60.5, 0.0, 77.0] SR:23 DR:3 LR:-60.48 LO:60.6);ALT=A[chr6:84603239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	85318151	+	chr6	85324221	+	.	63	54	2925877_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAATGT;MAPQ=60;MATEID=2925877_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_85309001_85334001_46C;SPAN=6070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:50 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:54 DR:63 LR:-267.4 LO:267.4);ALT=T[chr6:85324221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	86079896	-	chr6	86080952	+	.	8	0	2927493_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2927493_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:86079896(-)-6:86080952(-)__6_86068501_86093501D;SPAN=1056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=[chr6:86080952[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	86708754	+	chr6	86714792	+	.	60	28	2929141_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=AAGAAAATGTGGCAC;MAPQ=60;MATEID=2929141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_86705501_86730501_180C;SPAN=6038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:20 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:28 DR:60 LR:-260.8 LO:260.8);ALT=T[chr6:86714792[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
