chr19	7118388	-	chr19	7119667	+	.	8	0	10136329_1	0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=10136329_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7118388(-)-19:7119667(-)__19_7105001_7130001D;SPAN=1279;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr19:7119667[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
