chr11	134104947	+	chr11	134109884	+	.	2	3	5059864_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5059864_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_134088501_134113501_241C;SPAN=4937;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:3 DR:2 LR:6.574 LO:6.671);ALT=G[chr11:134109884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	134119817	+	chr11	134122734	+	GTAGTTACGAACACCATCCCAGCATGTTGTCTGTTTGGGCTGTGCTTTGAGATCCTCAATGCTGAACTTCACATCTACACCTTTCTCTAGGCGGCTCTCTGGCTCTGACTTCATCAGCCAGTGGCTGCTTAGATTCTTCAAACAGTTTTTAGTGGCTGAAGTCTTCTGAGGGTTGGAGTCCTCCACTTTAGCTAATGCCTCACCTGAGTTCTCAGTTTTGGTGCGTTTTCCTGATAGTCCCTTGT	0	32	5060073_1	83.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GTAGTTACGAACACCATCCCAGCATGTTGTCTGTTTGGGCTGTGCTTTGAGATCCTCAATGCTGAACTTCACATCTACACCTTTCTCTAGGCGGCTCTCTGGCTCTGACTTCATCAGCCAGTGGCTGCTTAGATTCTTCAAACAGTTTTTAGTGGCTGAAGTCTTCTGAGGGTTGGAGTCCTCCACTTTAGCTAATGCCTCACCTGAGTTCTCAGTTTTGGTGCGTTTTCCTGATAGTCCCTTGT;MAPQ=60;MATEID=5060073_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_134113001_134138001_363C;SPAN=2917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:84 GQ:83 PL:[83.0, 0.0, 119.3] SR:32 DR:0 LR:-82.88 LO:83.27);ALT=G[chr11:134122734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	134121248	+	chr11	134123120	+	.	35	0	5060078_1	97.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5060078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:134121248(+)-11:134123120(-)__11_134113001_134138001D;SPAN=1872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:67 GQ:64.4 PL:[97.4, 0.0, 64.4] SR:0 DR:35 LR:-97.72 LO:97.72);ALT=A[chr11:134123120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
