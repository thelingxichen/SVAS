chr2	174977755	-	chr2	174978868	+	.	8	0	1517085_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1517085_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:174977755(-)-2:174978868(-)__2_174954501_174979501D;SPAN=1113;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:174 GQ:20.5 PL:[0.0, 20.5, 462.1] SR:0 DR:8 LR:20.73 LO:12.72);ALT=[chr2:174978868[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	175928550	+	chr6	103027994	-	.	19	40	1521079_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATAAAG;MAPQ=60;MATEID=1521079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_175910001_175935001_27C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:40 DR:19 LR:-118.8 LO:118.8);ALT=G]chr6:103027994];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	176346682	+	chr2	176352722	+	.	109	27	1522530_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAAAATAAATGTTT;MAPQ=60;MATEID=1522530_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_176326501_176351501_289C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:123 DP:21 GQ:33 PL:[363.0, 33.0, 0.0] SR:27 DR:109 LR:-363.1 LO:363.1);ALT=T[chr2:176352722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	177265645	+	chr2	177272041	+	.	145	100	1526084_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TATT;MAPQ=60;MATEID=1526084_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_177257501_177282501_316C;SPAN=6396;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:207 DP:55 GQ:55.9 PL:[613.9, 55.9, 0.0] SR:100 DR:145 LR:-614.0 LO:614.0);ALT=T[chr2:177272041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
