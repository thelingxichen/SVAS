chr6	161273060	+	chr6	161268824	+	.	12	0	4471785_1	21.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4471785_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:161268824(-)-6:161273060(+)__6_161259001_161284001D;SPAN=4236;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:0 DR:12 LR:-21.19 LO:26.47);ALT=]chr6:161273060]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	161273588	+	chr6	161271139	+	.	15	0	4471797_1	30.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4471797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:161271139(-)-6:161273588(+)__6_161259001_161284001D;SPAN=2449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:70 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:0 DR:15 LR:-30.55 LO:34.51);ALT=]chr6:161273588]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	161602303	-	chr6	161603388	+	.	8	0	4471993_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4471993_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:161602303(-)-6:161603388(-)__6_161577501_161602501D;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=[chr6:161603388[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	162222618	+	chr6	162506783	+	.	93	78	4473160_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4473160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_162484001_162509001_40C;SPAN=284165;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:141 DP:13 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:78 DR:93 LR:-415.9 LO:415.9);ALT=G[chr6:162506783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	162536770	+	chr6	162929715	+	.	77	51	4473220_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;MAPQ=60;MATEID=4473220_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_162925001_162950001_1C;SPAN=392945;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:8 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:51 DR:77 LR:-300.4 LO:300.4);ALT=G[chr6:162929715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	163814230	+	chr8	75185139	-	.	11	38	5508230_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5508230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_75166001_75191001_25C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:46 DP:37 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:38 DR:11 LR:-135.3 LO:135.3);ALT=C]chr8:75185139];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr15	86556627	+	chr6	163903710	+	.	16	0	9044293_1	38.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=9044293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:163903710(-)-15:86556627(+)__15_86534001_86559001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:53 GQ:38.6 PL:[38.6, 0.0, 88.1] SR:0 DR:16 LR:-38.46 LO:39.6);ALT=]chr15:86556627]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	75362871	+	chr8	75367000	+	CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA	68	77	5508627_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA;MAPQ=60;MATEID=5508627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_75362001_75387001_106C;SPAN=4129;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:42 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:77 DR:68 LR:-346.6 LO:346.6);ALT=A[chr8:75367000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47057588	+	chr11	47063712	+	AAAGTGGGATAGTGGAATGCAC	0	84	6787940_1	99.0	.	EVDNC=ASSMB;INSERTION=AAAGTGGGATAGTGGAATGCAC;MAPQ=60;MATEID=6787940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47040001_47065001_175C;SPAN=6124;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:70 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:84 DR:0 LR:-247.6 LO:247.6);ALT=A[chr11:47063712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47768676	-	chr11	47836656	+	.	85	32	6793095_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=6793095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47824001_47849001_265C;SPAN=67980;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:110 DP:96 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:32 DR:85 LR:-326.8 LO:326.8);ALT=[chr11:47836656[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	47836639	+	chr11	47863419	-	.	79	22	6792421_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGCTAATTTTTGTATTTTT;MAPQ=33;MATEID=6792421_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47848501_47873501_29C;SPAN=26780;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:106 GQ:25.2 PL:[306.9, 25.2, 0.0] SR:22 DR:79 LR:-307.1 LO:307.1);ALT=C]chr11:47863419];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	47939382	+	chr11	47942807	+	.	86	62	6792830_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CGCC;MAPQ=60;MATEID=6792830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47922001_47947001_37C;SPAN=3425;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:120 DP:115 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:62 DR:86 LR:-356.5 LO:356.5);ALT=C[chr11:47942807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	86535784	+	chr11	48528022	+	.	11	26	9044296_1	82.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=9044296_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_15_86534001_86559001_390C;SECONDARY;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:28 DP:24 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:26 DR:11 LR:-82.52 LO:82.52);ALT=]chr15:86535784]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	48600858	+	chr11	48604283	+	.	67	58	6796710_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=6796710_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_48583501_48608501_415C;SPAN=3425;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:93 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:58 DR:67 LR:-303.7 LO:303.7);ALT=C[chr11:48604283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	48714063	+	chr11	48715074	+	.	0	25	6797099_1	63.0	.	EVDNC=ASSMB;HOMSEQ=AAACCTTTCTTTTCATTC;MAPQ=60;MATEID=6797099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_48706001_48731001_360C;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:71 GQ:63.5 PL:[63.5, 0.0, 106.4] SR:25 DR:0 LR:-63.29 LO:63.95);ALT=C[chr11:48715074[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	49204268	+	chr11	49884340	-	.	11	0	6804431_1	15.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6804431_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:49204268(+)-11:49884340(+)__11_49882001_49907001D;SPAN=680072;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:0 DR:11 LR:-15.45 LO:23.15);ALT=T]chr11:49884340];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	49899242	+	chr11	55660127	+	.	9	0	6804517_1	20.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=6804517_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:49899242(+)-11:55660127(-)__11_49882001_49907001D;SPAN=5760885;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:36 GQ:20 PL:[20.0, 0.0, 66.2] SR:0 DR:9 LR:-19.96 LO:21.4);ALT=G[chr11:55660127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	55660265	+	chr11	49899540	+	.	8	0	6804518_1	11.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6804518_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:49899540(-)-11:55660265(+)__11_49882001_49907001D;SPAN=5760725;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=]chr11:55660265]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	50488876	+	chr11	50490669	-	.	13	0	6806791_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6806791_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:50488876(+)-11:50490669(+)__11_50470001_50495001D;SPAN=1793;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:128 GQ:8.3 PL:[8.3, 0.0, 302.0] SR:0 DR:13 LR:-8.235 LO:25.3);ALT=C]chr11:50490669];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	50566393	+	chr11	50568347	-	.	14	0	6806992_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6806992_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:50566393(+)-11:50568347(+)__11_50543501_50568501D;SPAN=1954;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:127 GQ:11.9 PL:[11.9, 0.0, 295.7] SR:0 DR:14 LR:-11.81 LO:27.77);ALT=T]chr11:50568347];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	51254707	-	chr11	51258715	+	.	9	0	6809225_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6809225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:51254707(-)-11:51258715(-)__11_51254001_51279001D;SPAN=4008;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:128 GQ:4.8 PL:[0.0, 4.8, 320.1] SR:0 DR:9 LR:4.969 LO:16.01);ALT=[chr11:51258715[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	55084821	+	chr11	55196633	+	.	10	0	6812454_1	17.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6812454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:55084821(+)-11:55196633(-)__11_55174001_55199001D;SPAN=111812;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=T[chr11:55196633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	55360089	-	chr11	55431551	+	G	16	105	6813199_1	99.0	.	DISC_MAPQ=19;EVDNC=TSI_L;INSERTION=G;MAPQ=19;MATEID=6813199_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_11_55345501_55370501_4C;SPAN=71462;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:84 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:105 DR:16 LR:-323.5 LO:323.5);ALT=[chr11:55431551[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	55364889	-	chr11	55431551	+	CAGCCAAATCTCATCTTGAATTGTAGCTCCAGTAATTCCTATGTGG	51	160	6813218_1	99.0	.	DISC_MAPQ=5;EVDNC=TSI_G;INSERTION=CAGCCAAATCTCATCTTGAATTGTAGCTCCAGTAATTCCTATGTGG;MAPQ=19;MATEID=6813218_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_55345501_55370501_4C;SPAN=66662;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:189 DP:11 GQ:51.1 PL:[561.1, 51.1, 0.0] SR:160 DR:51 LR:-561.1 LO:561.1);ALT=[chr11:55431551[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	55365428	+	chr11	55445868	-	.	101	52	6813703_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=TTTT;MAPQ=60;MATEID=6813703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_55443501_55468501_47C;SPAN=80440;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:145 DP:19 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:52 DR:101 LR:-429.1 LO:429.1);ALT=T]chr11:55445868];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	55444016	-	chr11	55457756	+	.	67	125	6813708_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGTTT;MAPQ=60;MATEID=6813708_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_55443501_55468501_21C;SECONDARY;SPAN=13740;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:178 DP:53 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:125 DR:67 LR:-528.1 LO:528.1);ALT=[chr11:55457756[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
