chr10	26999055	+	chr10	27002150	+	.	18	0	6156261_1	35.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6156261_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:26999055(+)-10:27002150(-)__10_26999001_27024001D;SPAN=3095;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:87 GQ:35.9 PL:[35.9, 0.0, 174.5] SR:0 DR:18 LR:-35.85 LO:41.09);ALT=C[chr10:27002150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27154695	+	chr10	27156504	-	.	8	0	6157187_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6157187_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:27154695(+)-10:27156504(+)__10_27146001_27171001D;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:165 GQ:18.1 PL:[0.0, 18.1, 435.7] SR:0 DR:8 LR:18.29 LO:12.91);ALT=T]chr10:27156504];VARTYPE=BND:INV-hh;JOINTYPE=hh
