chr12	25259494	-	chr12	25260554	+	CATATACATATATATATATATATATATAT	33	68	7483366_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=ATATATATATGCAGAGA;INSERTION=CATATACATATATATATATATATATATAT;MAPQ=60;MATEID=7483366_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_12_25259501_25284501_246C;SECONDARY;SPAN=1060;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:89 DP:133 GQ:63.2 PL:[257.9, 0.0, 63.2] SR:68 DR:33 LR:-264.2 LO:264.2);ALT=[chr12:25260554[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	25956194	-	chr12	104359693	+	.	5	6	7487212_1	0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CTGGCAG;MAPQ=0;MATEID=7487212_2;MATENM=0;NM=1;NUMPARTS=2;REPSEQ=GG;SCTG=c_12_25945501_25970501_15C;SECONDARY;SPAN=78403499;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:174 GQ:17.2 PL:[0.0, 17.2, 455.5] SR:6 DR:5 LR:17.43 LO:14.78);ALT=[chr12:104359693[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	104359630	-	chr12	125801148	+	.	52	59	7892669_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;MAPQ=60;MATEID=7892669_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_125783001_125808001_312C;SPAN=21441518;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:57 GQ:24 PL:[264.0, 24.0, 0.0] SR:59 DR:52 LR:-264.1 LO:264.1);ALT=[chr12:125801148[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	104359839	+	chr12	104373609	+	.	22	0	7816398_1	62.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7816398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104359839(+)-12:104373609(-)__12_104370001_104395001D;SPAN=13770;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:36 GQ:23.3 PL:[62.9, 0.0, 23.3] SR:0 DR:22 LR:-63.79 LO:63.79);ALT=G[chr12:104373609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104378707	+	chr12	104380723	+	.	18	0	7816430_1	38.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=7816430_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104378707(+)-12:104380723(-)__12_104370001_104395001D;SPAN=2016;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:77 GQ:38.6 PL:[38.6, 0.0, 147.5] SR:0 DR:18 LR:-38.56 LO:42.19);ALT=C[chr12:104380723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104379506	+	chr12	104380726	+	.	32	48	7816433_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;MAPQ=26;MATEID=7816433_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_104370001_104395001_171C;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:62 DP:86 GQ:26.3 PL:[181.4, 0.0, 26.3] SR:48 DR:32 LR:-187.9 LO:187.9);ALT=A[chr12:104380726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
