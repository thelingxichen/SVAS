chr4	67122068	+	chr4	67123492	+	AGACCATCC	28	50	2740584_1	99.0	.	DISC_MAPQ=20;EVDNC=ASDIS;INSERTION=AGACCATCC;MAPQ=0;MATEID=2740584_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_67105501_67130501_344C;SECONDARY;SPAN=1424;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:26 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:50 DR:28 LR:-211.3 LO:211.3);ALT=G[chr4:67123492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
