chr5	109274627	+	chr5	109617414	+	.	40	50	3675752_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TT;MAPQ=60;MATEID=3675752_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_109613001_109638001_269C;SPAN=342787;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:53 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:50 DR:40 LR:-217.9 LO:217.9);ALT=T[chr5:109617414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
