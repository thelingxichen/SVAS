chr12	74014499	+	chr7	125264207	+	AATTGTTCAAAAAAAAAA	0	63	7745212_1	99.0	.	EVDNC=ASSMB;INSERTION=AATTGTTCAAAAAAAAAA;MAPQ=60;MATEID=7745212_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_73990001_74015001_307C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:63 DP:115 GQ:99 PL:[176.9, 0.0, 101.0] SR:63 DR:0 LR:-177.9 LO:177.9);ALT=]chr12:74014499]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	125264220	+	chr12	74014367	+	ATTATA	38	53	7745214_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTATA;MAPQ=60;MATEID=7745214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_73990001_74015001_493C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:102 GQ:25.4 PL:[220.1, 0.0, 25.4] SR:53 DR:38 LR:-228.6 LO:228.6);ALT=C[chr12:74014367[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	126045889	+	chr7	126051448	+	.	52	45	5274118_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=5274118_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_126028001_126053001_1C;SPAN=5559;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:16 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:45 DR:52 LR:-250.9 LO:250.9);ALT=C[chr7:126051448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	72189159	+	chr12	72190574	+	.	201	140	7729846_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7729846_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_12_72177001_72202001_32C;SPAN=1415;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:320 DP:71 GQ:86.6 PL:[950.6, 86.6, 0.0] SR:140 DR:201 LR:-950.6 LO:950.6);ALT=G[chr12:72190574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	72987377	-	chr12	72988957	+	.	8	0	7737051_1	0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=7737051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:72987377(-)-12:72988957(-)__12_72985501_73010501D;SPAN=1580;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:229 GQ:35.5 PL:[0.0, 35.5, 627.1] SR:0 DR:8 LR:35.63 LO:11.76);ALT=[chr12:72988957[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	73771177	+	chr12	73772793	+	.	51	35	7743571_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAA;MAPQ=60;MATEID=7743571_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_73769501_73794501_164C;SPAN=1616;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:69 DP:192 GQ:99 PL:[176.0, 0.0, 288.2] SR:35 DR:51 LR:-175.8 LO:177.3);ALT=A[chr12:73772793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
