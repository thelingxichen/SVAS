chr16	113799	+	chr16	345781	+	.	0	45	9115662_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=9115662_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_16_343001_368001_4C;SPAN=231982;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:45 DP:8 GQ:12 PL:[132.0, 12.0, 0.0] SR:45 DR:0 LR:-132.0 LO:132.0);ALT=C[chr16:345781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
