chr7	56021011	+	chr7	56022600	+	.	0	13	3320868_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3320868_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_56007001_56032001_374C;SPAN=1589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:13 DR:0 LR:-19.34 LO:27.64);ALT=G[chr7:56022600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56032395	+	chr7	56045818	+	.	22	5	3320922_1	60.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3320922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_56031501_56056501_50C;SPAN=13423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:70 GQ:60.2 PL:[60.2, 0.0, 109.7] SR:5 DR:22 LR:-60.26 LO:61.05);ALT=G[chr7:56045818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56045958	+	chr7	56049165	+	TTCACAATGTTAAACCGGAATGCCTAGAAGCATACAACAAAATTT	0	17	3320996_1	28.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTCACAATGTTAAACCGGAATGCCTAGAAGCATACAACAAAATTT;MAPQ=60;MATEID=3320996_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_56031501_56056501_298C;SPAN=3207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:102 GQ:28.7 PL:[28.7, 0.0, 216.8] SR:17 DR:0 LR:-28.48 LO:37.03);ALT=T[chr7:56049165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56119609	+	chr7	56122059	+	.	16	0	3321286_1	23.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3321286_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:56119609(+)-7:56122059(-)__7_56105001_56130001D;SPAN=2450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:108 GQ:23.6 PL:[23.6, 0.0, 238.1] SR:0 DR:16 LR:-23.56 LO:33.95);ALT=A[chr7:56122059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56122197	+	chr7	56123317	+	.	0	8	3321300_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=51;MATEID=3321300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_56105001_56130001_273C;SPAN=1120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:8 DR:0 LR:0.6845 LO:14.7);ALT=G[chr7:56123317[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56132072	+	chr7	56136173	+	.	50	7	3321369_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3321369_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_56129501_56154501_146C;SPAN=4101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:123 GQ:99 PL:[135.2, 0.0, 161.6] SR:7 DR:50 LR:-135.0 LO:135.2);ALT=G[chr7:56136173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56132098	+	chr7	56140687	+	.	19	0	3321370_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3321370_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:56132098(+)-7:56140687(-)__7_56129501_56154501D;SPAN=8589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:122 GQ:29.9 PL:[29.9, 0.0, 264.2] SR:0 DR:19 LR:-29.67 LO:40.77);ALT=G[chr7:56140687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56136332	+	chr7	56140688	+	.	0	35	3321393_1	89.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3321393_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_56129501_56154501_247C;SPAN=4356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:96 GQ:89.6 PL:[89.6, 0.0, 142.4] SR:35 DR:0 LR:-89.53 LO:90.21);ALT=G[chr7:56140688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56146202	+	chr7	56147218	+	.	4	4	3321462_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3321462_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_56129501_56154501_209C;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:121 GQ:12.6 PL:[0.0, 12.6, 316.8] SR:4 DR:4 LR:12.98 LO:9.741);ALT=G[chr7:56147218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56172181	+	chr7	56174069	+	.	131	0	3321888_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=3321888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:56172181(+)-7:56174069(-)__7_56154001_56179001D;SPAN=1888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:131 DP:148 GQ:33.4 PL:[425.8, 33.4, 0.0] SR:0 DR:131 LR:-427.5 LO:427.5);ALT=A[chr7:56174069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	56217755	+	chr7	56220248	+	.	26	0	3322089_1	73.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=3322089_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:56217755(+)-7:56220248(-)__7_56203001_56228001D;SPAN=2493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:47 GQ:40.1 PL:[73.1, 0.0, 40.1] SR:0 DR:26 LR:-73.58 LO:73.58);ALT=T[chr7:56220248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
