chr3	162213707	+	chr3	162235597	+	.	130	96	2451710_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2451710_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_162190001_162215001_329C;SPAN=21890;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:182 DP:17 GQ:49 PL:[538.0, 49.0, 0.0] SR:96 DR:130 LR:-538.0 LO:538.0);ALT=T[chr3:162235597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	162512134	+	chr3	162626351	+	AAATACTGTCTTCCC	0	48	2453055_1	99.0	.	EVDNC=ASSMB;INSERTION=AAATACTGTCTTCCC;MAPQ=60;MATEID=2453055_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_162606501_162631501_254C;SPAN=114217;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:35 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:48 DR:0 LR:-141.9 LO:141.9);ALT=C[chr3:162626351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	162545363	-	chr3	162547659	+	G	67	65	2452507_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=2452507_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_162533001_162558001_61C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:114 DP:28 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:65 DR:67 LR:-336.7 LO:336.7);ALT=[chr3:162547659[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	162764902	+	chr3	162769085	+	.	117	79	2453235_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=2453235_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_162753501_162778501_325C;SPAN=4183;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:152 DP:37 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:79 DR:117 LR:-448.9 LO:448.9);ALT=A[chr3:162769085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
