chr12	101799783	+	chr12	101801469	+	.	8	0	5311832_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5311832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:101799783(+)-12:101801469(-)__12_101797501_101822501D;SPAN=1686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=C[chr12:101801469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	102183836	+	chr12	102190454	+	.	0	7	5312958_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5312958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_102165001_102190001_325C;SPAN=6618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:33 GQ:14.3 PL:[14.3, 0.0, 63.8] SR:7 DR:0 LR:-14.17 LO:16.07);ALT=C[chr12:102190454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	102190542	+	chr12	102224334	+	.	0	14	5313173_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CACCT;MAPQ=60;MATEID=5313173_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_102214001_102239001_4C;SPAN=33792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:34 GQ:37.1 PL:[37.1, 0.0, 43.7] SR:14 DR:0 LR:-37.0 LO:37.05);ALT=T[chr12:102224334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	102506012	+	chr12	102512140	+	.	0	11	5313889_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5313889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_102508001_102533001_174C;SPAN=6128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:11 DR:0 LR:-24.12 LO:26.03);ALT=T[chr12:102512140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
