chrX	30819816	+	chrX	30813668	+	.	16	63	11053572_1	99.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=TGTGCCTTGCCTT;MAPQ=0;MATEID=11053572_2;MATENM=0;NM=1;NUMPARTS=2;REPSEQ=CCC;SCTG=c_23_30796501_30821501_343C;SECONDARY;SPAN=6148;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:77 DP:340 GQ:99 PL:[162.1, 0.0, 663.8] SR:63 DR:16 LR:-162.1 LO:179.2);ALT=]chrX:30819816]T;VARTYPE=BND:DUP-th;JOINTYPE=th
