chr3	71008542	+	chr3	71015040	+	.	0	7	1475292_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1475292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_71001001_71026001_180C;SPAN=6498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:105 GQ:5.1 PL:[0.0, 5.1, 264.0] SR:7 DR:0 LR:5.34 LO:12.29);ALT=C[chr3:71015040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71247545	+	chr3	71348969	+	.	0	13	1476587_1	29.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=1476587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_71344001_71369001_180C;SPAN=101424;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:13 DR:0 LR:-28.83 LO:30.91);ALT=T[chr3:71348969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71247588	+	chr3	71355108	+	.	15	0	1476588_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1476588_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:71247588(+)-3:71355108(-)__3_71344001_71369001D;SPAN=107520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:0 DR:15 LR:-34.89 LO:36.48);ALT=A[chr3:71355108[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71349032	+	chr3	71355028	+	.	10	12	1476614_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1476614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_71344001_71369001_209C;SPAN=5996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:106 GQ:37.4 PL:[37.4, 0.0, 218.9] SR:12 DR:10 LR:-37.3 LO:44.76);ALT=C[chr3:71355028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71542707	+	chr3	71630700	+	.	10	6	1477574_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1477574_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_71613501_71638501_168C;SPAN=87993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:53 GQ:38.6 PL:[38.6, 0.0, 88.1] SR:6 DR:10 LR:-38.46 LO:39.6);ALT=C[chr3:71630700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71630895	+	chr3	71632721	+	.	16	0	1477632_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1477632_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:71630895(+)-3:71632721(-)__3_71613501_71638501D;SPAN=1826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:120 GQ:20.3 PL:[20.3, 0.0, 271.1] SR:0 DR:16 LR:-20.31 LO:33.16);ALT=T[chr3:71632721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	71830744	+	chr3	71834107	+	.	47	46	1478576_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1478576_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_71834001_71859001_242C;SPAN=3363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:57 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:46 DR:47 LR:-194.7 LO:194.7);ALT=C[chr3:71834107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
