chr5	37379658	+	chr5	37381703	+	.	0	9	2454493_1	13.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=27;MATEID=2454493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_37362501_37387501_27C;SPAN=2045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:62 GQ:13.1 PL:[13.1, 0.0, 135.2] SR:9 DR:0 LR:-12.91 LO:19.01);ALT=T[chr5:37381703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
