chr5	174058021	+	chrX	126744483	-	.	10	0	7521283_1	26.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7521283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:174058021(+)-23:126744483(+)__23_126738501_126763501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:26 GQ:26 PL:[26.0, 0.0, 35.9] SR:0 DR:10 LR:-25.97 LO:26.07);ALT=A]chrX:126744483];VARTYPE=BND:TRX-hh;JOINTYPE=hh
