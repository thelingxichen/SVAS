chr2	172906237	+	chr2	172910236	+	.	39	49	1508077_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAATTAGCCGGGCGTGGTGG;MAPQ=60;MATEID=1508077_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_172896501_172921501_199C;SPAN=3999;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:80 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:49 DR:39 LR:-241.0 LO:241.0);ALT=G[chr2:172910236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	173004263	+	chr2	173007481	+	.	58	30	1508452_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTAGAGATGGGGTTT;MAPQ=60;MATEID=1508452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172994501_173019501_329C;SPAN=3218;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:77 DP:80 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:30 DR:58 LR:-237.7 LO:237.7);ALT=T[chr2:173007481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	173179996	+	chr2	173186105	+	.	54	30	1510758_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=AGAATCTTTTCTTTGTC;MAPQ=60;MATEID=1510758_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_2_173166001_173191001_31C;SPAN=6109;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:70 DP:102 GQ:41.9 PL:[203.6, 0.0, 41.9] SR:30 DR:54 LR:-209.2 LO:209.2);ALT=C[chr2:173186105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
