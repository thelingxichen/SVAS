chr7	141786241	+	chr7	141759848	+	.	30	0	5307106_1	89.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5307106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:141759848(-)-7:141786241(+)__7_141781501_141806501D;SPAN=26393;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:30 DP:11 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=]chr7:141786241]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	141760577	+	chr7	141786875	+	.	36	0	5307107_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5307107_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:141760577(+)-7:141786875(-)__7_141781501_141806501D;SPAN=26298;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:36 DP:12 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=T[chr7:141786875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142359260	-	chr7	142362014	+	.	14	46	5307846_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=AAG;MAPQ=60;MATEID=5307846_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_7_142345001_142370001_212C;SPAN=2754;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:51 DP:45 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:46 DR:14 LR:-148.5 LO:148.5);ALT=[chr7:142362014[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	142359543	+	chr7	142360546	-	.	9	0	5307849_1	19.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5307849_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:142359543(+)-7:142360546(+)__7_142345001_142370001D;SPAN=1003;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=A]chr7:142360546];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	142360600	+	chr7	142362013	+	.	41	0	5307853_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5307853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:142360600(+)-7:142362013(-)__7_142345001_142370001D;SPAN=1413;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:8 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=A[chr7:142362013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
