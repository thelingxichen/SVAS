chr10	71281030	+	chr10	71291093	+	.	182	81	6340581_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=60;MATEID=6340581_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_71270501_71295501_95C;SPAN=10063;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:237 DP:63 GQ:64 PL:[703.0, 64.0, 0.0] SR:81 DR:182 LR:-703.1 LO:703.1);ALT=C[chr10:71291093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	71731235	+	chr13	91986528	-	.	3	9	6342391_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6342391_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_71711501_71736501_212C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:9 DR:3 LR:-15.67 LO:21.47);ALT=T]chr13:91986528];VARTYPE=BND:TRX-hh;JOINTYPE=hh
