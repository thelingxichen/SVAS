chr11	92869804	+	chr11	92875914	+	ATACATAAC	72	47	4962300_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=ATACATAAC;MAPQ=60;MATEID=4962300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_92855001_92880001_198C;SPAN=6110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:34 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:47 DR:72 LR:-307.0 LO:307.0);ALT=T[chr11:92875914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93471718	+	chr11	93474582	+	.	17	0	4963314_1	30.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4963314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:93471718(+)-11:93474582(-)__11_93467501_93492501D;SPAN=2864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:96 GQ:30.2 PL:[30.2, 0.0, 201.8] SR:0 DR:17 LR:-30.11 LO:37.52);ALT=C[chr11:93474582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93472499	+	chr11	93474488	+	.	0	68	4963316_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4963316_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_93467501_93492501_361C;SPAN=1989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:105 GQ:57.5 PL:[196.1, 0.0, 57.5] SR:68 DR:0 LR:-200.1 LO:200.1);ALT=T[chr11:93474488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93474939	+	chr11	93483509	+	.	8	0	4963324_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4963324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:93474939(+)-11:93483509(-)__11_93467501_93492501D;SPAN=8570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:0 DR:8 LR:-8.527 LO:16.22);ALT=A[chr11:93483509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93480614	+	chr11	93483510	+	.	0	8	4963338_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4963338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_93467501_93492501_51C;SPAN=2896;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:8 DR:0 LR:-9.611 LO:16.46);ALT=G[chr11:93483510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	93679244	+	chr11	93681424	+	.	67	42	4964104_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCCTGTTGGATTCTT;MAPQ=60;MATEID=4964104_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_11_93663501_93688501_142C;SPAN=2180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:38 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:42 DR:67 LR:-260.8 LO:260.8);ALT=T[chr11:93681424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94224131	+	chr11	94226850	+	AGTGCATCTGCAGTACTCATTTTTATGGTCAGTCAAGCTCCTCTGGGACCAGGTTCTTCTCCAAGAACCCCTGGGTACTGTACTCAAATGTCAGAAAATGCACTCGATTCCAAATTCTAGAAATT	0	17	4965091_1	37.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGTGCATCTGCAGTACTCATTTTTATGGTCAGTCAAGCTCCTCTGGGACCAGGTTCTTCTCCAAGAACCCCTGGGTACTGTACTCAAATGTCAGAAAATGCACTCGATTCCAAATTCTAGAAATT;MAPQ=60;MATEID=4965091_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_94202501_94227501_12C;SPAN=2719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:70 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:17 DR:0 LR:-37.15 LO:40.17);ALT=A[chr11:94226850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94696681	+	chr11	94699458	+	.	0	26	4966369_1	63.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4966369_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_94692501_94717501_53C;SPAN=2777;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:83 GQ:63.5 PL:[63.5, 0.0, 136.1] SR:26 DR:0 LR:-63.34 LO:64.87);ALT=T[chr11:94699458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94699579	+	chr11	94704140	+	TCCTGGCCTGCTCTTCAGCTCTTTCTTTTTTAATTTTTTCCAGTTCTGCAAGAAGAGCTGCAGTATCATCATCATCACTTTCTTCTTCAAAATCTTCATCTTCCT	0	14	4966381_1	27.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCCTGGCCTGCTCTTCAGCTCTTTCTTTTTTAATTTTTTCCAGTTCTGCAAGAAGAGCTGCAGTATCATCATCATCACTTTCTTCTTCAAAATCTTCATCTTCCT;MAPQ=60;MATEID=4966381_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_11_94692501_94717501_141C;SPAN=4561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:14 DR:0 LR:-27.52 LO:31.83);ALT=T[chr11:94704140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94699579	+	chr11	94703152	+	.	2	6	4966380_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=4966380_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CC;SCTG=c_11_94692501_94717501_141C;SPAN=3573;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:6 DR:2 LR:-8.527 LO:16.22);ALT=T[chr11:94703152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94704280	+	chr11	94706660	+	.	10	0	4966395_1	8.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4966395_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:94704280(+)-11:94706660(-)__11_94692501_94717501D;SPAN=2380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=T[chr11:94706660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94704702	+	chr11	94706660	+	.	23	0	4966398_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4966398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:94704702(+)-11:94706660(-)__11_94692501_94717501D;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:97 GQ:49.7 PL:[49.7, 0.0, 185.0] SR:0 DR:23 LR:-49.64 LO:54.07);ALT=A[chr11:94706660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	94705386	+	chr11	94706660	+	.	35	0	4966399_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4966399_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:94705386(+)-11:94706660(-)__11_94692501_94717501D;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:0 DR:35 LR:-91.97 LO:92.16);ALT=T[chr11:94706660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	95523907	+	chr11	95532395	+	.	0	12	4968249_1	28.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4968249_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_95525501_95550501_81C;SPAN=8488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:40 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:12 DR:0 LR:-28.78 LO:29.66);ALT=G[chr11:95532395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
