chr8	133769583	+	chr8	133772721	+	.	9	0	4084471_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4084471_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:133769583(+)-8:133772721(-)__8_133770001_133795001D;SPAN=3138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=A[chr8:133772721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	133771163	+	chr8	133772722	+	.	14	9	4084474_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4084474_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TCTC;SCTG=c_8_133770001_133795001_222C;SPAN=1559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:93 GQ:27.8 PL:[27.8, 0.0, 196.1] SR:9 DR:14 LR:-27.62 LO:35.09);ALT=T[chr8:133772722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
