chr5	67160818	+	chr5	66936736	+	A	5	7	3494322_1	8.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=A;MAPQ=5;MATEID=3494322_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_67154501_67179501_231C;SPAN=224082;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:7 DR:5 LR:-8.035 LO:17.94);ALT=]chr5:67160818]G;VARTYPE=BND:DUP-th;JOINTYPE=th
