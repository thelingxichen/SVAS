chr12	37991228	+	chr12	37994618	+	.	50	37	5153842_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=AGAGCAGTTTTGAAACACT;MAPQ=60;MATEID=5153842_2;MATENM=1;NM=1;NUMPARTS=3;SCTG=c_12_37975001_38000001_51C;SPAN=3390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:20 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:37 DR:50 LR:-221.2 LO:221.2);ALT=T[chr12:37994618[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	38010175	+	chr12	38018062	+	.	49	0	5153882_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=5153882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:38010175(+)-12:38018062(-)__12_37999501_38024501D;SPAN=7887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:9 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:49 LR:-145.2 LO:145.2);ALT=A[chr12:38018062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
