chr2	30473684	-	chr2	30474809	+	.	8	0	950787_1	9.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=950787_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:30473684(-)-2:30474809(-)__2_30453501_30478501D;SPAN=1125;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=[chr2:30474809[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
