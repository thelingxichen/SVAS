chrX	56756022	+	chrX	56843751	+	TCTTTGAGTGATTGCAGTATGACTCCATTTCCCTGGTGCATTCATATAATAGTTCACCTGGTGAAAACAATGAAGATTATTTACAATGCTACCCTGCTTTTTCTGGTGTCCTGAACCTGGAAGTTGTGCTTTTTA	7	51	7430930_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TCTTTGAGTGATTGCAGTATGACTCCATTTCCCTGGTGCATTCATATAATAGTTCACCTGGTGAAAACAATGAAGATTATTTACAATGCTACCCTGCTTTTTCTGGTGTCCTGAACCTGGAAGTTGTGCTTTTTA;MAPQ=60;MATEID=7430930_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_56840001_56865001_229C;SPAN=87729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:40 GQ:15 PL:[165.0, 15.0, 0.0] SR:51 DR:7 LR:-165.0 LO:165.0);ALT=G[chrX:56843751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	56756022	+	chrX	56758493	+	.	9	25	7430748_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=7430748_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_56742001_56767001_244C;SPAN=2471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:59 GQ:53.3 PL:[89.6, 0.0, 53.3] SR:25 DR:9 LR:-90.14 LO:90.14);ALT=G[chrX:56758493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	56758632	+	chrX	56843751	+	.	7	30	7430931_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=7430931_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_56840001_56865001_229C;SPAN=85119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:30 DR:7 LR:-118.8 LO:118.8);ALT=G[chrX:56843751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
