chr11	56731202	-	chr11	56732499	+	.	5	3	6818439_1	0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=ATCTGATCTTTGACAAACCTGA;MAPQ=24;MATEID=6818439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_56717501_56742501_203C;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:116 GQ:4.8 PL:[0.0, 4.8, 290.4] SR:3 DR:5 LR:5.019 LO:14.16);ALT=[chr11:56732499[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
