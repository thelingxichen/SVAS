chr5	142780464	+	chr5	142783970	+	.	14	0	2601618_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2601618_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:142780464(+)-5:142783970(-)__5_142761501_142786501D;SPAN=3506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:48 GQ:33.2 PL:[33.2, 0.0, 82.7] SR:0 DR:14 LR:-33.21 LO:34.4);ALT=A[chr5:142783970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	143545168	+	chr5	143549410	+	.	0	7	2602562_1	17.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2602562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_143545501_143570501_99C;SPAN=4242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:22 GQ:17.3 PL:[17.3, 0.0, 33.8] SR:7 DR:0 LR:-17.15 LO:17.52);ALT=T[chr5:143549410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
