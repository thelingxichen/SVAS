chr9	9058751	+	chr15	25855251	+	.	7	40	5905740_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=GAG;MAPQ=41;MATEID=5905740_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_25847501_25872501_67C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:21 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:40 DR:7 LR:-128.7 LO:128.7);ALT=G[chr15:25855251[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
