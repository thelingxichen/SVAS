chr2	50814528	+	chr2	50816643	-	.	32	0	790092_1	86.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=790092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:50814528(+)-2:50816643(+)__2_50813001_50838001D;SPAN=2115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:73 GQ:86 PL:[86.0, 0.0, 89.3] SR:0 DR:32 LR:-85.86 LO:85.87);ALT=A]chr2:50816643];VARTYPE=BND:INV-hh;JOINTYPE=hh
