chrX	78620055	+	chrX	78577497	+	.	8	7	11262494_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=11262494_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_78596001_78621001_140C;SPAN=42558;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:64 GQ:19.1 PL:[19.1, 0.0, 134.6] SR:7 DR:8 LR:-18.97 LO:24.12);ALT=]chrX:78620055]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	78680098	+	chrX	78682204	+	GA	12	6	11262926_1	11.0	.	DISC_MAPQ=40;EVDNC=ASDIS;INSERTION=GA;MAPQ=60;MATEID=11262926_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_78669501_78694501_234C;SPAN=2106;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:141 GQ:11.6 PL:[11.6, 0.0, 328.4] SR:6 DR:12 LR:-11.31 LO:29.51);ALT=T[chrX:78682204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	78921889	+	chrX	78923365	-	.	35	59	11263759_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GA;MAPQ=60;MATEID=11263759_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_78914501_78939501_161C;SPAN=1476;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:97 GQ:6.3 PL:[247.5, 6.3, 0.0] SR:59 DR:35 LR:-257.5 LO:257.5);ALT=A]chrX:78923365];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	78921938	+	chrX	78926076	+	.	23	0	11263760_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=11263760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:78921938(+)-23:78926076(-)__23_78914501_78939501D;SPAN=4138;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:65 GQ:58.4 PL:[58.4, 0.0, 98.0] SR:0 DR:23 LR:-58.31 LO:58.9);ALT=T[chrX:78926076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	78923226	-	chrX	78926077	+	.	30	68	11263761_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CAT;MAPQ=60;MATEID=11263761_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_23_78914501_78939501_178C;SPAN=2851;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:78 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:68 DR:30 LR:-254.2 LO:254.2);ALT=[chrX:78926077[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
