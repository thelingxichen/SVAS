chr2	214874705	+	chr2	214876214	+	.	17	12	1192543_1	62.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=1192543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_214865001_214890001_320C;SPAN=1509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:60 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:12 DR:17 LR:-62.97 LO:63.12);ALT=G[chr2:214876214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
