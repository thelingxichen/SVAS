chr11	107923528	+	chr11	107925373	+	.	0	7	4994911_1	4.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4994911_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_107922501_107947501_284C;SPAN=1845;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:69 GQ:4.4 PL:[4.4, 0.0, 162.8] SR:7 DR:0 LR:-4.413 LO:13.62);ALT=G[chr11:107925373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	107992406	+	chr11	108002631	+	.	5	6	4995514_1	12.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=4995514_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_107971501_107996501_199C;SPAN=10225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:6 DR:5 LR:-12.54 LO:15.5);ALT=G[chr11:108002631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	107992406	+	chr11	108004545	+	AAATAAGATATGTGGAACGGAGTTATGTATCAAAACCCACTTTGA	31	24	4995515_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAATAAGATATGTGGAACGGAGTTATGTATCAAAACCCACTTTGA;MAPQ=60;MATEID=4995515_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_107971501_107996501_199C;SPAN=12139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:24 DR:31 LR:-115.5 LO:115.5);ALT=G[chr11:108004545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	108361896	+	chr11	108368890	+	.	4	3	4996062_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4996062_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_108339001_108364001_66C;SPAN=6994;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:33 GQ:7.7 PL:[7.7, 0.0, 70.4] SR:3 DR:4 LR:-7.565 LO:10.66);ALT=T[chr11:108368890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
