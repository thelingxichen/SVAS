chr12	19503508	-	chr12	19506199	+	.	10	0	7447921_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=7447921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:19503508(-)-12:19506199(-)__12_19502001_19527001D;SPAN=2691;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:239 GQ:31.6 PL:[0.0, 31.6, 643.6] SR:0 DR:10 LR:31.74 LO:15.49);ALT=[chr12:19506199[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
