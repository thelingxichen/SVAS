chr6	75950132	+	chr6	75953433	+	.	90	0	2905707_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2905707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:75950132(+)-6:75953433(-)__6_75950001_75975001D;SPAN=3301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:81 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:0 DR:90 LR:-267.4 LO:267.4);ALT=A[chr6:75953433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	75951030	+	chr6	75953435	+	.	55	0	2905711_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=2905711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:75951030(+)-6:75953435(-)__6_75950001_75975001D;SPAN=2405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:94 GQ:70.4 PL:[156.2, 0.0, 70.4] SR:0 DR:55 LR:-157.8 LO:157.8);ALT=A[chr6:75953435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	76489702	-	chr6	76490792	+	.	8	0	2907154_1	4.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=2907154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:76489702(-)-6:76490792(-)__6_76489001_76514001D;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:0 DR:8 LR:-4.192 LO:15.42);ALT=[chr6:76490792[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	77097496	+	chr6	77102642	+	.	77	47	2908364_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTAT;MAPQ=60;MATEID=2908364_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_6_77077001_77102001_158C;SPAN=5146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:11 GQ:27 PL:[297.0, 27.0, 0.0] SR:47 DR:77 LR:-297.1 LO:297.1);ALT=T[chr6:77102642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	77437200	+	chr6	77459050	+	.	12	0	2909027_1	36.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=2909027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:77437200(+)-6:77459050(-)__6_77444501_77469501D;SPAN=21850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:15 GQ:0.6 PL:[36.3, 0.6, 0.0] SR:0 DR:12 LR:-37.56 LO:37.56);ALT=G[chr6:77459050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
