chr19	27933683	+	chr19	27930485	+	.	10	0	10232854_1	15.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=10232854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:27930485(-)-19:27933683(+)__19_27905501_27930501D;SPAN=3198;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:65 GQ:15.5 PL:[15.5, 0.0, 140.9] SR:0 DR:10 LR:-15.4 LO:21.4);ALT=]chr19:27933683]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	27957073	+	chr19	27960383	+	.	33	35	10233085_1	99.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=CCAAACACCACAT;MAPQ=33;MATEID=10233085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_27954501_27979501_256C;SPAN=3310;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:99 GQ:82.1 PL:[158.0, 0.0, 82.1] SR:35 DR:33 LR:-159.3 LO:159.3);ALT=T[chr19:27960383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	27961383	+	chr19	27963247	+	.	58	45	10233092_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTTTTACACCATAGGCCTCA;MAPQ=60;MATEID=10233092_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_27954501_27979501_44C;SPAN=1864;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:104 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:45 DR:58 LR:-307.0 LO:307.0);ALT=A[chr19:27963247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
