chr10	109449439	+	chr10	109462254	+	.	9	0	4686052_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4686052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:109449439(+)-10:109462254(-)__10_109441501_109466501D;SPAN=12815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:0 DR:9 LR:-17.25 LO:20.3);ALT=T[chr10:109462254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
