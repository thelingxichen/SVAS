chr7	158062156	+	chr7	158073629	+	.	70	40	5359707_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=5359707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_158074001_158099001_182C;SPAN=11473;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:0 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:40 DR:70 LR:-247.6 LO:247.6);ALT=C[chr7:158073629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
