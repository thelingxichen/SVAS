chr1	93291056	+	chr1	93292095	-	.	10	0	420915_1	13.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=420915_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93291056(+)-1:93292095(+)__1_93271501_93296501D;SPAN=1039;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:0 DR:10 LR:-13.5 LO:20.92);ALT=G]chr1:93292095];VARTYPE=BND:INV-hh;JOINTYPE=hh
