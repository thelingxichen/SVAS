chr11	134732900	+	chr11	134734113	+	.	198	173	7313627_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=7313627_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_134725501_134750501_240C;SPAN=1213;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:298 DP:67 GQ:80.6 PL:[884.6, 80.6, 0.0] SR:173 DR:198 LR:-884.6 LO:884.6);ALT=T[chr11:134734113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
