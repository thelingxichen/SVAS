chr10	85598460	+	chr10	85601788	-	.	17	44	6403939_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCCAGCACTTTGGGAGGCCGAGGTGGGCGG;MAPQ=49;MATEID=6403939_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_10_85578501_85603501_304C;SPAN=3328;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:131 GQ:99 PL:[129.8, 0.0, 185.9] SR:44 DR:17 LR:-129.6 LO:130.2);ALT=G]chr10:85601788];VARTYPE=BND:INV-hh;JOINTYPE=hh
