chr21	43547905	+	chr21	43549822	+	.	11	0	7186549_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7186549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:43547905(+)-21:43549822(-)__21_43536501_43561501D;SPAN=1917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:90 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:0 DR:11 LR:-11.93 LO:22.35);ALT=C[chr21:43549822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	43547950	+	chr21	43557517	+	.	9	0	7186550_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7186550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:43547950(+)-21:43557517(-)__21_43536501_43561501D;SPAN=9567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:82 GQ:7.7 PL:[7.7, 0.0, 189.2] SR:0 DR:9 LR:-7.493 LO:17.84);ALT=T[chr21:43557517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	43549912	+	chr21	43557547	+	.	0	11	7186557_1	16.0	.	EVDNC=ASSMB;HOMSEQ=AGGTGAG;MAPQ=60;MATEID=7186557_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_43536501_43561501_268C;SPAN=7635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:11 DR:0 LR:-16.26 LO:23.36);ALT=G[chr21:43557547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	43639351	+	chr21	43645783	+	.	8	0	7186724_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7186724_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:43639351(+)-21:43645783(-)__21_43634501_43659501D;SPAN=6432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=C[chr21:43645783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	43934087	+	chr21	43938384	+	.	17	0	7187637_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7187637_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:43934087(+)-21:43938384(-)__21_43928501_43953501D;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.57 LO:43.16);ALT=G[chr21:43938384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	43938622	+	chr21	43945885	+	.	0	7	7187649_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7187649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_43928501_43953501_321C;SPAN=7263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:7 DR:0 LR:1.005 LO:12.81);ALT=T[chr21:43945885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44050100	+	chr21	44048681	+	.	25	0	7188010_1	61.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=7188010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:44048681(-)-21:44050100(+)__21_44026501_44051501D;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:78 GQ:61.4 PL:[61.4, 0.0, 127.4] SR:0 DR:25 LR:-61.39 LO:62.68);ALT=]chr21:44050100]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	44313491	+	chr21	44317035	+	.	11	2	7189273_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7189273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_44296001_44321001_436C;SPAN=3544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:67 GQ:18.2 PL:[18.2, 0.0, 143.6] SR:2 DR:11 LR:-18.16 LO:23.88);ALT=G[chr21:44317035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44313511	+	chr21	44328971	+	.	13	0	7189274_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7189274_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:44313511(+)-21:44328971(-)__21_44296001_44321001D;SPAN=15460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:28 GQ:32 PL:[35.3, 0.0, 32.0] SR:0 DR:13 LR:-35.33 LO:35.33);ALT=G[chr21:44328971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44313515	+	chr21	44323291	+	.	9	0	7189275_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7189275_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:44313515(+)-21:44323291(-)__21_44296001_44321001D;SPAN=9776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:0 DR:9 LR:-22.12 LO:22.58);ALT=T[chr21:44323291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44317157	+	chr21	44328974	+	.	0	20	7189287_1	54.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7189287_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_44296001_44321001_471C;SPAN=11817;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:42 GQ:44.9 PL:[54.8, 0.0, 44.9] SR:20 DR:0 LR:-54.67 LO:54.67);ALT=A[chr21:44328974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44515902	+	chr21	44527559	+	.	20	0	7189692_1	56.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=7189692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:44515902(+)-21:44527559(-)__21_44516501_44541501D;SPAN=11657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:36 GQ:29.9 PL:[56.3, 0.0, 29.9] SR:0 DR:20 LR:-56.66 LO:56.66);ALT=C[chr21:44527559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44521545	+	chr21	44524425	+	.	0	45	7189713_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7189713_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_44516501_44541501_70C;SPAN=2880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:113 GQ:99 PL:[118.1, 0.0, 154.4] SR:45 DR:0 LR:-117.9 LO:118.2);ALT=G[chr21:44524425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44521594	+	chr21	44527565	+	.	26	0	7189715_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7189715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:44521594(+)-21:44527565(-)__21_44516501_44541501D;SPAN=5971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:96 GQ:59.9 PL:[59.9, 0.0, 172.1] SR:0 DR:26 LR:-59.82 LO:62.88);ALT=A[chr21:44527565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44524512	+	chr21	44527561	+	.	35	22	7189720_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;MAPQ=52;MATEID=7189720_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_44516501_44541501_116C;SPAN=3049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:84 GQ:83 PL:[119.3, 0.0, 83.0] SR:22 DR:35 LR:-119.5 LO:119.5);ALT=T[chr21:44527561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	44970368	+	chr21	44973301	+	.	64	33	7190723_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GAGA;MAPQ=60;MATEID=7190723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_44957501_44982501_159C;SPAN=2933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:46 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:33 DR:64 LR:-247.6 LO:247.6);ALT=A[chr21:44973301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45079676	+	chr21	45089762	+	.	0	7	7191128_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=7191128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45080001_45105001_16C;SPAN=10086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:7 DR:0 LR:-12.54 LO:15.5);ALT=G[chr21:45089762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45194642	+	chr21	45196082	+	.	167	27	7191517_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=7191517_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45178001_45203001_96C;SPAN=1440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:77 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:27 DR:167 LR:-514.9 LO:514.9);ALT=T[chr21:45196082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45422724	+	chr21	45423854	-	.	5	2	7192226_1	4.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TGCCTGGCCTT;MAPQ=60;MATEID=7192226_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45423001_45448001_207C;SPAN=1130;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:45 GQ:4.4 PL:[4.4, 0.0, 103.4] SR:2 DR:5 LR:-4.313 LO:9.938);ALT=A]chr21:45423854];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr21	45553662	+	chr21	45555940	+	.	45	0	7192623_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7192623_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:45553662(+)-21:45555940(-)__21_45545501_45570501D;SPAN=2278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:102 GQ:99 PL:[121.1, 0.0, 124.4] SR:0 DR:45 LR:-120.9 LO:120.9);ALT=C[chr21:45555940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45556056	+	chr21	45557056	+	.	3	12	7192632_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=7192632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45545501_45570501_247C;SPAN=1000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:76 GQ:29 PL:[29.0, 0.0, 154.4] SR:12 DR:3 LR:-28.92 LO:33.9);ALT=G[chr21:45557056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45560224	+	chr21	45563086	+	.	9	8	7192645_1	23.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7192645_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45545501_45570501_355C;SPAN=2862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:72 GQ:23.6 PL:[23.6, 0.0, 149.0] SR:8 DR:9 LR:-23.41 LO:28.82);ALT=G[chr21:45563086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45619169	+	chr21	45620717	+	GGGAGGCTGAGGCAGAAGAACCACT	51	54	7193032_1	99.0	.	DISC_MAPQ=49;EVDNC=TSI_G;HOMSEQ=TGAAC;INSERTION=GGGAGGCTGAGGCAGAAGAACCACT;MAPQ=60;MATEID=7193032_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_21_45594501_45619501_142C;SPAN=1548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:12 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:54 DR:51 LR:-293.8 LO:293.8);ALT=C[chr21:45620717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45720057	+	chr21	45731986	+	.	16	0	7192908_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7192908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:45720057(+)-21:45731986(-)__21_45717001_45742001D;SPAN=11929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:46 GQ:40.4 PL:[40.4, 0.0, 70.1] SR:0 DR:16 LR:-40.35 LO:40.82);ALT=C[chr21:45731986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45720074	+	chr21	45730887	+	CATGAACGCTGCTGTCCGGGCTGTGACGCGCATGGGCATTTATGTGGGTGCCAAAGTCTTCCTCATCTACG	27	45	7192910_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CATGAACGCTGCTGTCCGGGCTGTGACGCGCATGGGCATTTATGTGGGTGCCAAAGTCTTCCTCATCTACG;MAPQ=60;MATEID=7192910_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_45717001_45742001_30C;SPAN=10813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:66 GQ:4.5 PL:[168.3, 4.5, 0.0] SR:45 DR:27 LR:-174.7 LO:174.7);ALT=G[chr21:45730887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45720074	+	chr21	45726562	+	.	27	10	7192909_1	75.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=7192909_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_21_45717001_45742001_30C;SPAN=6488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:52 GQ:48.8 PL:[75.2, 0.0, 48.8] SR:10 DR:27 LR:-75.28 LO:75.28);ALT=G[chr21:45726562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	45730967	+	chr21	45731987	+	.	0	20	7192934_1	43.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=7192934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_45717001_45742001_286C;SPAN=1020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:83 GQ:43.7 PL:[43.7, 0.0, 155.9] SR:20 DR:0 LR:-43.53 LO:47.18);ALT=G[chr21:45731987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46191407	+	chr21	46193462	+	.	3	3	7194392_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7194392_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46182501_46207501_359C;SPAN=2055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:91 GQ:11.1 PL:[0.0, 11.1, 240.9] SR:3 DR:3 LR:11.45 LO:6.281);ALT=G[chr21:46193462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46197381	+	chr21	46221630	+	.	18	0	7194458_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7194458_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46197381(+)-21:46221630(-)__21_46207001_46232001D;SPAN=24249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:30 GQ:21.5 PL:[51.2, 0.0, 21.5] SR:0 DR:18 LR:-51.95 LO:51.95);ALT=C[chr21:46221630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46208073	+	chr21	46221630	+	.	11	0	7194463_1	19.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7194463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46208073(+)-21:46221630(-)__21_46207001_46232001D;SPAN=13557;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:0 DR:11 LR:-19.51 LO:24.29);ALT=A[chr21:46221630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46226959	+	chr21	46233890	+	GCTGGAGTGTCAGTTTCATTGATTGGCTGCCCGTCGAACCTGAATCTGATCTGCCTCATTGACAAGC	0	96	7194530_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=GCTGGAGTGTCAGTTTCATTGATTGGCTGCCCGTCGAACCTGAATCTGATCTGCCTCATTGACAAGC;MAPQ=60;MATEID=7194530_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_46231501_46256501_68C;SPAN=6931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:47 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:96 DR:0 LR:-283.9 LO:283.9);ALT=T[chr21:46233890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46227000	+	chr21	46237906	+	.	13	0	7194531_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7194531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46227000(+)-21:46237906(-)__21_46231501_46256501D;SPAN=10906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:39 GQ:32.3 PL:[32.3, 0.0, 62.0] SR:0 DR:13 LR:-32.35 LO:32.87);ALT=T[chr21:46237906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46229036	+	chr21	46233890	+	.	3	68	7194532_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=7194532_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_21_46231501_46256501_68C;SPAN=4854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:47 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:68 DR:3 LR:-204.7 LO:204.7);ALT=G[chr21:46233890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46229086	+	chr21	46237861	+	.	43	0	7194533_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7194533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46229086(+)-21:46237861(-)__21_46231501_46256501D;SPAN=8775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:16 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=A[chr21:46237861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46234021	+	chr21	46237862	+	.	102	34	7194539_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7194539_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46231501_46256501_164C;SPAN=3841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:53 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:34 DR:102 LR:-326.8 LO:326.8);ALT=T[chr21:46237862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46276280	+	chr21	46281078	+	.	15	27	7194879_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7194879_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46256001_46281001_373C;SPAN=4798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:44 GQ:1.4 PL:[103.7, 0.0, 1.4] SR:27 DR:15 LR:-109.4 LO:109.4);ALT=C[chr21:46281078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46281238	+	chr21	46293471	+	.	22	0	7194607_1	49.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7194607_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46281238(+)-21:46293471(-)__21_46280501_46305501D;SPAN=12233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:86 GQ:49.4 PL:[49.4, 0.0, 158.3] SR:0 DR:22 LR:-49.32 LO:52.57);ALT=A[chr21:46293471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46285418	+	chr21	46293470	+	.	17	0	7194620_1	34.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7194620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46285418(+)-21:46293470(-)__21_46280501_46305501D;SPAN=8052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:81 GQ:34.4 PL:[34.4, 0.0, 159.8] SR:0 DR:17 LR:-34.17 LO:38.93);ALT=T[chr21:46293470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46306819	+	chr21	46308608	+	.	16	9	7194990_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7194990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_241C;SPAN=1789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:100 GQ:42.2 PL:[42.2, 0.0, 200.6] SR:9 DR:16 LR:-42.23 LO:48.1);ALT=T[chr21:46308608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46310140	+	chr21	46311721	+	.	10	10	7194999_1	39.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CACCTG;MAPQ=60;MATEID=7194999_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_21_46305001_46330001_204C;SPAN=1581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:75 GQ:39.2 PL:[39.2, 0.0, 141.5] SR:10 DR:10 LR:-39.1 LO:42.43);ALT=G[chr21:46311721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46311912	+	chr21	46313319	+	.	7	6	7195004_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7195004_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_21_46305001_46330001_204C;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:6 DR:7 LR:-9.982 LO:20.14);ALT=C[chr21:46313319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46313459	+	chr21	46314886	+	.	2	4	7195010_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=7195010_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_75C;SPAN=1427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:54 GQ:2 PL:[2.0, 0.0, 127.4] SR:4 DR:2 LR:-1.875 LO:9.519);ALT=T[chr21:46314886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46314977	+	chr21	46318982	+	.	2	3	7195014_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7195014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_79C;SPAN=4005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:62 GQ:0 PL:[0.0, 0.0, 148.5] SR:3 DR:2 LR:0.2923 LO:9.206);ALT=T[chr21:46318982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46320391	+	chr21	46321406	+	.	16	12	7195033_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=7195033_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_354C;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:60 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:12 DR:16 LR:-62.97 LO:63.12);ALT=C[chr21:46321406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46321649	+	chr21	46323279	+	.	13	8	7195037_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=7195037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_371C;SPAN=1630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:101 GQ:32.3 PL:[32.3, 0.0, 210.5] SR:8 DR:13 LR:-32.05 LO:39.78);ALT=C[chr21:46323279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46323453	+	chr21	46326829	+	.	0	9	7195045_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=7195045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46305001_46330001_181C;SPAN=3376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:9 DR:0 LR:-6.951 LO:17.74);ALT=G[chr21:46326829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46327011	+	chr21	46330199	+	.	0	98	7194690_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7194690_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46329501_46354501_357C;SPAN=3188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:77 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:98 DR:0 LR:-290.5 LO:290.5);ALT=C[chr21:46330199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46327062	+	chr21	46340733	+	.	74	0	7195058_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7195058_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46327062(+)-21:46340733(-)__21_46305001_46330001D;SPAN=13671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:31 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:0 DR:74 LR:-217.9 LO:217.9);ALT=G[chr21:46340733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46330701	+	chr21	46340735	+	.	116	12	7194697_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=7194697_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CC;SCTG=c_21_46329501_46354501_270C;SPAN=10034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:93 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:12 DR:116 LR:-346.6 LO:346.6);ALT=C[chr21:46340735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46360102	+	chr21	46363597	+	.	0	19	7194761_1	41.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7194761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_46354001_46379001_160C;SPAN=3495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:79 GQ:41.3 PL:[41.3, 0.0, 150.2] SR:19 DR:0 LR:-41.32 LO:44.8);ALT=G[chr21:46363597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	46957868	+	chr21	46962282	+	.	8	0	7196332_1	13.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7196332_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:46957868(+)-21:46962282(-)__21_46942001_46967001D;SPAN=4414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=C[chr21:46962282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	47012808	+	chr21	47011273	+	.	8	0	7196482_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7196482_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:47011273(-)-21:47012808(+)__21_46991001_47016001D;SPAN=1535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:122 GQ:6.3 PL:[0.0, 6.3, 306.9] SR:0 DR:8 LR:6.645 LO:13.98);ALT=]chr21:47012808]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	47235664	+	chr21	47234175	+	.	41	0	7197435_1	99.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=7197435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:47234175(-)-21:47235664(+)__21_47211501_47236501D;SPAN=1489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:126 GQ:99 PL:[101.3, 0.0, 203.6] SR:0 DR:41 LR:-101.2 LO:103.1);ALT=]chr21:47235664]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	47588574	+	chr21	47604270	+	.	70	7	7198409_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7198409_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_47603501_47628501_296C;SPAN=15696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:50 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:7 DR:70 LR:-208.0 LO:208.0);ALT=T[chr21:47604270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	47657352	+	chr21	47658674	+	.	63	78	7198496_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=7198496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_47652501_47677501_351C;SPAN=1322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:34 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:78 DR:63 LR:-359.8 LO:359.8);ALT=T[chr21:47658674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	47711378	+	chr21	47717450	+	GACGGCCACCCACGGACTCTGTCACTTGCTGGGATTCACACACGGCACGGAGGCAGAGTGGCAG	0	16	7199026_1	33.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=GACGGCCACCCACGGACTCTGTCACTTGCTGGGATTCACACACGGCACGGAGGCAGAGTGGCAG;MAPQ=60;MATEID=7199026_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_47701501_47726501_338C;SPAN=6072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:72 GQ:33.5 PL:[33.5, 0.0, 139.1] SR:16 DR:0 LR:-33.31 LO:37.09);ALT=T[chr21:47717450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48019418	+	chr21	48022190	+	.	3	62	7199686_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7199686_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_21_47995501_48020501_54C;SPAN=2772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:55 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:62 DR:3 LR:-191.4 LO:191.4);ALT=T[chr21:48022190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48019466	+	chr21	48024931	+	.	69	0	7199687_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7199687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:48019466(+)-21:48024931(-)__21_47995501_48020501D;SPAN=5465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:44 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:0 DR:69 LR:-204.7 LO:204.7);ALT=G[chr21:48024931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48022331	+	chr21	48024925	+	.	64	14	7199712_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7199712_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_48020001_48045001_29C;SPAN=2594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:90 GQ:8.6 PL:[209.9, 0.0, 8.6] SR:14 DR:64 LR:-221.2 LO:221.2);ALT=T[chr21:48024925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48055675	+	chr21	48056806	+	.	22	5	7199793_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7199793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_48044501_48069501_33C;SPAN=1131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:103 GQ:51.5 PL:[51.5, 0.0, 196.7] SR:5 DR:22 LR:-51.32 LO:56.21);ALT=G[chr21:48056806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48055718	+	chr21	48063442	+	.	36	0	7199795_1	87.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7199795_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:48055718(+)-21:48063442(-)__21_48044501_48069501D;SPAN=7724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:117 GQ:87.2 PL:[87.2, 0.0, 196.1] SR:0 DR:36 LR:-87.14 LO:89.47);ALT=A[chr21:48063442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48056903	+	chr21	48063443	+	.	5	38	7199799_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCAGG;MAPQ=60;MATEID=7199799_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_21_48044501_48069501_31C;SPAN=6540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:91 GQ:99 PL:[110.9, 0.0, 107.6] SR:38 DR:5 LR:-110.7 LO:110.7);ALT=G[chr21:48063443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	48056947	+	chr21	48064213	+	.	8	0	7199801_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7199801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:48056947(+)-21:48064213(-)__21_48044501_48069501D;SPAN=7266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=G[chr21:48064213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
