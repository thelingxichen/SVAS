chr21	33623598	-	chr21	33624610	+	.	8	0	10756488_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=10756488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:33623598(-)-21:33624610(-)__21_33614001_33639001D;SPAN=1012;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:0 DR:8 LR:5.29 LO:14.13);ALT=[chr21:33624610[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
