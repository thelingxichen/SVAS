chr9	101309048	+	chr9	101311665	+	.	48	56	5941142_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCTCA;MAPQ=60;MATEID=5941142_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_101307501_101332501_215C;SPAN=2617;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:20 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:56 DR:48 LR:-254.2 LO:254.2);ALT=A[chr9:101311665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
