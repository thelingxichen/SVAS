chr4	88847164	-	chr4	88858700	+	A	71	62	2781227_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=2781227_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_88837001_88862001_219C;SPAN=11536;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:110 DP:33 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:62 DR:71 LR:-326.8 LO:326.8);ALT=[chr4:88858700[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	89497059	+	chr4	89542720	+	.	74	42	2782337_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGG;MAPQ=60;MATEID=2782337_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_89474001_89499001_61C;SPAN=45661;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:8 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:42 DR:74 LR:-290.5 LO:290.5);ALT=G[chr4:89542720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
