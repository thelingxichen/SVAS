chr1	194451086	+	chr1	194454312	+	.	11	0	471845_1	29.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=471845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:194451086(+)-1:194454312(-)__1_194432001_194457001D;SPAN=3226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:11 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:11 LR:-29.71 LO:29.71);ALT=T[chr1:194454312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
