chr2	146862621	+	chr2	146876863	+	.	24	17	1031847_1	96.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=1031847_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_146853001_146878001_230C;SPAN=14242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:57 GQ:40.7 PL:[96.8, 0.0, 40.7] SR:17 DR:24 LR:-97.99 LO:97.99);ALT=T[chr2:146876863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
