chr15	39372396	+	chr15	39373461	+	.	114	11	8860650_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TTCTCCTGCCTCAGCCTCCCGAGTAGCTGGGATTACAGGCAT;MAPQ=60;MATEID=8860650_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_15_39347001_39372001_252C;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:123 DP:0 GQ:33 PL:[363.0, 33.0, 0.0] SR:11 DR:114 LR:-363.1 LO:363.1);ALT=T[chr15:39373461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
