chrX	23685928	+	chrX	23689646	+	.	0	18	7382373_1	43.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7382373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_23667001_23692001_31C;SPAN=3718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:18 DR:0 LR:-43.7 LO:44.82);ALT=A[chrX:23689646[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23697404	+	chrX	23700511	+	.	2	9	7382476_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7382476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_23691501_23716501_9C;SPAN=3107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:9 DR:2 LR:-23.31 LO:25.67);ALT=G[chrX:23700511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23700643	+	chrX	23704402	+	TCTGCCCTGCTGGCTGGAAACCTGGTAGTGAAACA	0	40	7382486_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TCTGCCCTGCTGGCTGGAAACCTGGTAGTGAAACA;MAPQ=60;MATEID=7382486_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_23691501_23716501_122C;SPAN=3759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:63 GQ:35.9 PL:[115.1, 0.0, 35.9] SR:40 DR:0 LR:-117.1 LO:117.1);ALT=G[chrX:23704402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23749105	+	chrX	23761241	+	CCAGTTTGTGGATGCTCCTACTATCTCCCGCAACTTATCTCGAACATGATTCACATGTATAGATGAACATGCTTCATGAATGTGGAAGATTCCCTGTTTCTTGGGGTTCTGGGGTCCTTGAGTCAGTCCTCTTCCAGGAGTAAGCTGCCCTTTGCCCAAGGCACAAAG	3	23	7382597_1	61.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CCAGTTTGTGGATGCTCCTACTATCTCCCGCAACTTATCTCGAACATGATTCACATGTATAGATGAACATGCTTCATGAATGTGGAAGATTCCCTGTTTCTTGGGGTTCTGGGGTCCTTGAGTCAGTCCTCTTCCAGGAGTAAGCTGCCCTTTGCCCAAGGCACAAAG;MAPQ=60;MATEID=7382597_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_23740501_23765501_4C;SPAN=12136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:66 GQ:61.4 PL:[61.4, 0.0, 97.7] SR:23 DR:3 LR:-61.34 LO:61.82);ALT=T[chrX:23761241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23754183	+	chrX	23761319	+	.	21	0	7382608_1	50.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7382608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:23754183(+)-23:23761319(-)__23_23740501_23765501D;SPAN=7136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:69 GQ:50.6 PL:[50.6, 0.0, 116.6] SR:0 DR:21 LR:-50.63 LO:52.07);ALT=C[chrX:23761319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23802001	+	chrX	23803443	+	.	11	10	7382922_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7382922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_23789501_23814501_37C;SPAN=1442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:20 DP:294 GQ:13.3 PL:[0.0, 13.3, 739.3] SR:10 DR:11 LR:13.63 LO:35.29);ALT=G[chrX:23803443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	23899071	+	chrX	23925809	+	.	0	8	7382976_1	19.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=7382976_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_23887501_23912501_211C;SPAN=26738;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:25 GQ:19.7 PL:[19.7, 0.0, 39.5] SR:8 DR:0 LR:-19.64 LO:20.05);ALT=T[chrX:23925809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	24073159	+	chrX	24075747	+	.	15	0	7383406_1	34.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7383406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:24073159(+)-23:24075747(-)__23_24059001_24084001D;SPAN=2588;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:56 GQ:34.4 PL:[34.4, 0.0, 100.4] SR:0 DR:15 LR:-34.34 LO:36.19);ALT=G[chrX:24075747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	24073164	+	chrX	24075532	+	.	44	0	7383407_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=7383407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:24073164(+)-23:24075532(-)__23_24059001_24084001D;SPAN=2368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:57 GQ:7.7 PL:[129.8, 0.0, 7.7] SR:0 DR:44 LR:-136.1 LO:136.1);ALT=T[chrX:24075532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
