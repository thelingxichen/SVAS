chr4	115175128	+	chr4	115183836	+	.	32	18	2855878_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=2855878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_115150001_115175001_312C;SPAN=8708;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:0 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:18 DR:32 LR:-141.9 LO:141.9);ALT=A[chr4:115183836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115507821	+	chr4	115511041	+	.	19	47	2856376_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2856376_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_115493001_115518001_103C;SPAN=3220;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:81 GQ:34.4 PL:[159.8, 0.0, 34.4] SR:47 DR:19 LR:-163.9 LO:163.9);ALT=G[chr4:115511041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115507821	+	chr4	115513865	+	TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT	43	76	2856377_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=GGTTATGTAGGGGTTTTCACACAAAAGCCCTTGATATCTTAACATCCTAGGGTTAGAAAGCCAGCGATGCCCACTCTGCTCCATCAGGGTGA;INSERTION=TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT;MAPQ=60;MATEID=2856377_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_115493001_115518001_103C;SECONDARY;SPAN=6044;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:108 DP:83 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:76 DR:43 LR:-320.2 LO:320.2);ALT=G[chr4:115513865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115511096	+	chr4	115513865	+	GTTGAGT	11	31	2856382_1	98.0	.	DISC_MAPQ=38;EVDNC=TSI_L;HOMSEQ=AG;INSERTION=GTTGAGT;MAPQ=44;MATEID=2856382_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_4_115493001_115518001_103C;SPAN=2769;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:89 GQ:98 PL:[98.0, 0.0, 117.8] SR:31 DR:11 LR:-98.03 LO:98.13);ALT=G[chr4:115513865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115890302	+	chr4	115891635	+	.	5	6	2858033_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=2858033_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_115885001_115910001_127C;SPAN=1333;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:128 GQ:8.1 PL:[0.0, 8.1, 326.7] SR:6 DR:5 LR:8.27 LO:13.81);ALT=T[chr4:115891635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115928723	+	chr4	115931874	+	.	139	119	2858160_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTGA;MAPQ=60;MATEID=2858160_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_115909501_115934501_342C;SPAN=3151;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:211 DP:43 GQ:56.8 PL:[623.8, 56.8, 0.0] SR:119 DR:139 LR:-623.9 LO:623.9);ALT=A[chr4:115931874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	116166907	+	chr4	116177181	+	GAATCAGAAAGCTAAGAAAAGACTGCCTGAATGTAAATTAGCCTGACAAATTATAATAGCACTTCTCATTTCTAAG	30	78	2858725_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GAATA;INSERTION=GAATCAGAAAGCTAAGAAAAGACTGCCTGAATGTAAATTAGCCTGACAAATTATAATAGCACTTCTCATTTCTAAG;MAPQ=60;MATEID=2858725_2;MATENM=4;NM=1;NUMPARTS=3;SCTG=c_4_116154501_116179501_265C;SPAN=10274;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:78 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:78 DR:30 LR:-287.2 LO:287.2);ALT=A[chr4:116177181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	116166907	+	chr4	116172035	-	.	14	44	2858724_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TTA;MAPQ=60;MATEID=2858724_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_116154501_116179501_265C;SPAN=5128;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:70 GQ:17.3 PL:[152.6, 0.0, 17.3] SR:44 DR:14 LR:-159.0 LO:159.0);ALT=A]chr4:116172035];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	116171952	-	chr4	116177181	+	.	20	38	2858728_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GAATA;MAPQ=60;MATEID=2858728_2;MATENM=4;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_116154501_116179501_265C;SPAN=5229;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:51 DP:56 GQ:15 PL:[165.0, 15.0, 0.0] SR:38 DR:20 LR:-165.0 LO:165.0);ALT=[chr4:116177181[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
