chr4	148357049	-	chr4	148391407	+	.	8	0	2260749_1	12.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=2260749_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:148357049(-)-4:148391407(-)__4_148347501_148372501D;SPAN=34358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.59 LO:17.19);ALT=[chr4:148391407[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
