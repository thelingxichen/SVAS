chr3	87276706	+	chr3	87294863	+	ATGTAATAAAGGAACAGAATCGAGAGTTACGAGGTACACAGAGGGCTATAATCAGAGATCGAGCAGCTTTAGAGAAACAAGAAAAACAGCT	2	10	1524919_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATGTAATAAAGGAACAGAATCGAGAGTTACGAGGTACACAGAGGGCTATAATCAGAGATCGAGCAGCTTTAGAGAAACAAGAAAAACAGCT;MAPQ=60;MATEID=1524919_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_87269001_87294001_372C;SPAN=18157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:10 DR:2 LR:-18.65 LO:22.38);ALT=G[chr3:87294863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	87276706	+	chr3	87289848	+	.	4	6	1524918_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1524918_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_87269001_87294001_372C;SPAN=13142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:112 GQ:3.6 PL:[0.0, 3.6, 277.2] SR:6 DR:4 LR:3.936 LO:14.29);ALT=G[chr3:87289848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	87842420	+	chr3	87871155	+	.	14	0	1526550_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1526550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:87842420(+)-3:87871155(-)__3_87857001_87882001D;SPAN=28735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:45 GQ:34.1 PL:[34.1, 0.0, 73.7] SR:0 DR:14 LR:-34.02 LO:34.88);ALT=A[chr3:87871155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	88199335	+	chr3	88202378	+	.	8	8	1527714_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1527714_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_3_88175501_88200501_87C;SPAN=3043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:8 DR:8 LR:-21.68 LO:25.03);ALT=G[chr3:88202378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
