chr1	63195091	+	chr1	63196336	-	.	8	0	305156_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=305156_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:63195091(+)-1:63196336(+)__1_63185501_63210501D;SPAN=1245;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:123 GQ:6.6 PL:[0.0, 6.6, 310.2] SR:0 DR:8 LR:6.916 LO:13.95);ALT=A]chr1:63196336];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	64291837	+	chr1	64188218	+	.	70	57	309740_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GTT;MAPQ=60;MATEID=309740_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_64165501_64190501_3C;SPAN=103619;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:78 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:57 DR:70 LR:-300.4 LO:300.4);ALT=]chr1:64291837]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	64839517	-	chr1	64854683	+	.	48	0	312920_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=312920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:64839517(-)-1:64854683(-)__1_64851501_64876501D;SPAN=15166;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:48 DP:90 GQ:84.5 PL:[134.0, 0.0, 84.5] SR:0 DR:48 LR:-134.7 LO:134.7);ALT=[chr1:64854683[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	65461603	-	chr10	3293111	+	.	8	0	6065527_1	5.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6065527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3283001_3308001_155C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:77 GQ:5.6 PL:[5.6, 0.0, 180.5] SR:0 DR:8 LR:-5.547 LO:15.65);ALT=[chr10:3293111[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	66024188	+	chr1	66030268	+	.	66	44	318493_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTTTCTTAATGTTTT;MAPQ=60;MATEID=318493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_66003001_66028001_275C;SPAN=6080;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:27 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:44 DR:66 LR:-260.8 LO:260.8);ALT=T[chr1:66030268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	66263923	+	chr2	196672057	+	.	10	44	1599941_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTTTTAGTAGAGATGGGGTTTCACCATGTTGGCCAGGCTAGTCTT;MAPQ=60;MATEID=1599941_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_196661501_196686501_63C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:88 GQ:62 PL:[151.1, 0.0, 62.0] SR:44 DR:10 LR:-153.1 LO:153.1);ALT=T[chr2:196672057[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	196672162	+	chr1	66264255	+	.	27	0	319234_1	79.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=319234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:66264255(-)-2:196672162(+)__1_66248001_66273001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:27 DP:25 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:0 DR:27 LR:-79.22 LO:79.22);ALT=]chr2:196672162]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	67297604	+	chr1	67001359	+	.	57	22	323751_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=323751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_67277001_67302001_404C;SPAN=296245;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:65 DP:81 GQ:1.4 PL:[192.8, 0.0, 1.4] SR:22 DR:57 LR:-203.7 LO:203.7);ALT=]chr1:67297604]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	197613646	-	chr2	197614859	+	.	17	0	1604328_1	26.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=1604328_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:197613646(-)-2:197614859(-)__2_197592501_197617501D;SPAN=1213;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:111 GQ:26.3 PL:[26.3, 0.0, 240.8] SR:0 DR:17 LR:-26.04 LO:36.34);ALT=[chr2:197614859[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	198328510	+	chr2	198330045	-	.	9	0	1607558_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1607558_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198328510(+)-2:198330045(+)__2_198303001_198328001D;SPAN=1535;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:9 DP:0 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=T]chr2:198330045];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	198629113	-	chr2	198630526	+	.	9	0	1608490_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1608490_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198629113(-)-2:198630526(-)__2_198621501_198646501D;SPAN=1413;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:134 GQ:6.3 PL:[0.0, 6.3, 336.6] SR:0 DR:9 LR:6.595 LO:15.83);ALT=[chr2:198630526[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	4290063	+	chr10	4291683	+	.	92	70	6067387_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6067387_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_4287501_4312501_146C;SPAN=1620;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:131 DP:23 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:70 DR:92 LR:-386.2 LO:386.2);ALT=C[chr10:4291683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	4708518	+	chr10	4710523	+	ATAG	59	38	6068109_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=ATAG;MAPQ=60;MATEID=6068109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_4704001_4729001_54C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:15 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:38 DR:59 LR:-241.0 LO:241.0);ALT=T[chr10:4710523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
