chr3	135969294	+	chr3	135974697	+	.	10	0	1672762_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1672762_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:135969294(+)-3:135974697(-)__3_135950501_135975501D;SPAN=5403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:121 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.2281 LO:18.52);ALT=G[chr3:135974697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	136021013	+	chr3	136026200	+	A	0	58	1673010_1	99.0	.	EVDNC=ASSMB;INSERTION=A;MAPQ=60;MATEID=1673010_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_136024001_136049001_275C;SPAN=5187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:34 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:58 DR:0 LR:-171.6 LO:171.6);ALT=C[chr3:136026200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	136349825	+	chr3	136471036	+	.	12	11	1674704_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1674704_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_136465001_136490001_120C;SPAN=121211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:11 DR:12 LR:-44.2 LO:44.37);ALT=T[chr3:136471036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	136462111	-	chr3	136463729	+	.	9	0	1674690_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=1674690_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:136462111(-)-3:136463729(-)__3_136440501_136465501D;SPAN=1618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:117 GQ:1.8 PL:[0.0, 1.8, 287.1] SR:0 DR:9 LR:1.989 LO:16.38);ALT=[chr3:136463729[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	136581195	+	chr3	136646824	+	.	21	4	1675382_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1675382_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_136636501_136661501_362C;SPAN=65629;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:52 GQ:58.7 PL:[65.3, 0.0, 58.7] SR:4 DR:21 LR:-65.14 LO:65.14);ALT=G[chr3:136646824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	137314508	+	chr3	137316442	+	.	65	0	1677698_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1677698_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:137314508(+)-3:137316442(-)__3_137298001_137323001D;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:80 GQ:1.4 PL:[192.8, 0.0, 1.4] SR:0 DR:65 LR:-204.6 LO:204.6);ALT=G[chr3:137316442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	137906485	+	chr3	137940766	+	.	9	0	1679653_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1679653_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:137906485(+)-3:137940766(-)__3_137886001_137911001D;SPAN=34281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:0 DR:9 LR:-14.27 LO:19.37);ALT=T[chr3:137940766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	138478203	+	chr3	138553536	+	.	5	2	1682443_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1682443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_138547501_138572501_25C;SPAN=75333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:62 GQ:0 PL:[0.0, 0.0, 148.5] SR:2 DR:5 LR:0.2923 LO:9.206);ALT=T[chr3:138553536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	139063040	+	chr3	139065719	+	.	17	12	1684038_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1684038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_139062001_139087001_235C;SPAN=2679;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:121 GQ:36.8 PL:[36.8, 0.0, 254.6] SR:12 DR:17 LR:-36.54 LO:46.15);ALT=G[chr3:139065719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	139071634	+	chr3	139075759	+	AATCGATGATGCAACCAACTTGGTCCAGCTGTATCACGTGCTCCATCCAGATGGCCAGTCGGCTCAAGGGGCCAAGGATCAGGCTGCTGAGGGAATAAATTTAATCA	0	13	1684068_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=AATCGATGATGCAACCAACTTGGTCCAGCTGTATCACGTGCTCCATCCAGATGGCCAGTCGGCTCAAGGGGCCAAGGATCAGGCTGCTGAGGGAATAAATTTAATCA;MAPQ=60;MATEID=1684068_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_139062001_139087001_380C;SPAN=4125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:99 GQ:16.1 PL:[16.1, 0.0, 224.0] SR:13 DR:0 LR:-16.09 LO:26.85);ALT=T[chr3:139075759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	139102278	+	chr3	139108390	+	.	6	2	1684261_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1684261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_139086501_139111501_30C;SPAN=6112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:98 GQ:3.3 PL:[0.0, 3.3, 244.2] SR:2 DR:6 LR:3.444 LO:12.5);ALT=C[chr3:139108390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
