chr13	34253777	+	chr13	34261029	+	.	11	0	5450022_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5450022_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:34253777(+)-13:34261029(-)__13_34251001_34276001D;SPAN=7252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:0 DR:11 LR:-9.219 LO:21.81);ALT=T[chr13:34261029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	34392405	+	chr13	34395268	+	.	4	4	5450296_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=5450296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_34373501_34398501_47C;SPAN=2863;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:97 GQ:9.6 PL:[0.0, 9.6, 254.1] SR:4 DR:4 LR:9.775 LO:8.204);ALT=G[chr13:34395268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
