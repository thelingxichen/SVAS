chr19	12550964	+	chr19	12404721	+	.	11	0	10165960_1	21.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=10165960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12404721(-)-19:12550964(+)__19_12544001_12569001D;SPAN=146243;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=]chr19:12550964]C;VARTYPE=BND:DUP-th;JOINTYPE=th
