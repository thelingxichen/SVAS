chr18	23794221	+	chr3	129912866	+	.	20	23	2320436_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=11;MATEID=2320436_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_129899001_129924001_265C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:38 DP:21 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:23 DR:20 LR:-112.2 LO:112.2);ALT=]chr18:23794221]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	129916635	-	chr3	129917734	+	.	8	0	2320486_1	0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2320486_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:129916635(-)-3:129917734(-)__3_129899001_129924001D;SPAN=1099;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:151 GQ:14.2 PL:[0.0, 14.2, 392.7] SR:0 DR:8 LR:14.5 LO:13.22);ALT=[chr3:129917734[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	23747813	+	chr18	23751323	+	.	71	60	9943277_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGTATTTT;MAPQ=60;MATEID=9943277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_23740501_23765501_96C;SPAN=3510;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:90 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:60 DR:71 LR:-326.8 LO:326.8);ALT=T[chr18:23751323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	23763005	+	chr18	23766102	+	.	58	0	9943895_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=9943895_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:23763005(+)-18:23766102(-)__18_23765001_23790001D;SPAN=3097;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:40 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=A[chr18:23766102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
