chr22	26878256	+	chr22	26879660	+	.	13	0	7248154_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7248154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:26878256(+)-22:26879660(-)__22_26876501_26901501D;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:88 GQ:19.1 PL:[19.1, 0.0, 194.0] SR:0 DR:13 LR:-19.07 LO:27.57);ALT=G[chr22:26879660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	26937701	+	chr22	26986015	+	.	32	0	7248459_1	93.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7248459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:26937701(+)-22:26986015(-)__22_26974501_26999501D;SPAN=48314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:45 GQ:14.3 PL:[93.5, 0.0, 14.3] SR:0 DR:32 LR:-96.59 LO:96.59);ALT=A[chr22:26986015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	27168076	+	chr22	27169793	+	.	56	41	7249571_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTTAACCTCT;MAPQ=60;MATEID=7249571_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_22_27146001_27171001_125C;SPAN=1717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:61 GQ:21 PL:[231.0, 21.0, 0.0] SR:41 DR:56 LR:-231.1 LO:231.1);ALT=T[chr22:27169793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
