chr3	106178797	-	chr11	31230228	+	.	37	23	10011507_1	99.0	.	BX=CCGGCAAGTAGGCTCC-1_1,AGCCGTGCACCAACCG-1_1,GATGAGGGTAAACCTC-1_2,GGGTCTGAGTGTCCAT-1_1,ACGCCAGCAATTAAGG-1_1,AGGCGAATCCTATTCA-1_1,CACCAAAAGGAAAGGT-1_1,CATGGCGGTCGTTGGC-1_2,TCGAATGTCCGTCTAC-1_1,GTCCAAAGTTAGAATG-1_2,ATCTCCGTCGACGAAG-1_3,CGATGGCAGGATGTCG-1_1,ATGGGAGCAGTGTAGG-1_5,GGACAGAAGTCTCGGC-1_1,TTCCATAAGCCCGTGT-1_1,TCAACGATCTGAGTAC-1_1,TTCTCCTCAGGGTCAA-1_1,CATATGGTCGTTATCT-1_1,CTGCTGTCAATCGCAT-1_1,CTTATACAGTACCTGT-1_1,AACGTTGGTAGCAAAT-1_1,ACGTATGGTCAAGCGA-1_1,AGGGAACCACACTAAC-1_1,AGCGTATTCTTTCCTC-1_2,TTCGCTGGTGGAAAGA-1_1,GCCGGATAGCTGCATT-1_1,TACTCGCGTGCACCAC-1_1,ACACCAACACAACGGA-1_3,GTGCAGCTCTATGGTG-1_1,GTACGTATCTGAAGCT-1_1,CATCGTCGTCCTGGAC-1_1,GTTCGAAGTACTAGGG-1_1,TGACTTTTCTATGGCA-1_1,GAGCTCGAGGAGCGAG-1_2;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=10011507_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_31213001_31238001_77C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:25 GQ:6.9 PL:[0.0, 6.9, 75.9] SR:0 DR:0 LR:7.024 LO:0.0),OC001T.bam(GT:1/1 AD:50 DP:28 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:23 DR:37 LR:-151.8 LO:151.8);ALT=[chr11:31230228[g;VARTYPE=BND:TRX-hh;JOINTYPE=hh	.
chr3	106178797	-	chr11	31230228	+	.	37	23	10011507_1	99.0	.	BX=CCGGCAAGTAGGCTCC-1_1,AGCCGTGCACCAACCG-1_1,GATGAGGGTAAACCTC-1_2,GGGTCTGAGTGTCCAT-1_1,ACGCCAGCAATTAAGG-1_1,AGGCGAATCCTATTCA-1_1,CACCAAAAGGAAAGGT-1_1,CATGGCGGTCGTTGGC-1_2,TCGAATGTCCGTCTAC-1_1,GTCCAAAGTTAGAATG-1_2,ATCTCCGTCGACGAAG-1_3,CGATGGCAGGATGTCG-1_1,ATGGGAGCAGTGTAGG-1_5,GGACAGAAGTCTCGGC-1_1,TTCCATAAGCCCGTGT-1_1,TCAACGATCTGAGTAC-1_1,TTCTCCTCAGGGTCAA-1_1,CATATGGTCGTTATCT-1_1,CTGCTGTCAATCGCAT-1_1,CTTATACAGTACCTGT-1_1,AACGTTGGTAGCAAAT-1_1,ACGTATGGTCAAGCGA-1_1,AGGGAACCACACTAAC-1_1,AGCGTATTCTTTCCTC-1_2,TTCGCTGGTGGAAAGA-1_1,GCCGGATAGCTGCATT-1_1,TACTCGCGTGCACCAC-1_1,ACACCAACACAACGGA-1_3,GTGCAGCTCTATGGTG-1_1,GTACGTATCTGAAGCT-1_1,CATCGTCGTCCTGGAC-1_1,GTTCGAAGTACTAGGG-1_1,TGACTTTTCTATGGCA-1_1,GAGCTCGAGGAGCGAG-1_2;DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=10011507_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_31213001_31238001_77C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:25 GQ:6.9 PL:[0.0, 6.9, 75.9] SR:0 DR:0 LR:7.024 LO:0.0),OC001T.bam(GT:1/1 AD:50 DP:28 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:23 DR:37 LR:-151.8 LO:151.8);ALT=[chr11:31230228[g;VARTYPE=BND:TRX-hh;JOINTYPE=hh	.
