chr7	54820113	+	chr7	54823472	+	.	3	138	3316122_1	99.0	.	DISC_MAPQ=44;EVDNC=TSI_L;MAPQ=60;MATEID=3316122_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ACCACC;SCTG=c_7_54806501_54831501_329C;SPAN=3359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:141 DP:204 GQ:54.3 PL:[311.8, 0.0, 54.3] SR:138 DR:3 LR:-323.6 LO:323.6);ALT=A[chr7:54823472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	54820113	+	chr7	54825188	+	ACAATGATGTTATTAATAGGAATATGGATCAATTTCACAAAGAAGCCAATGAATCCCATTATAGCAAATCCTATTGCTGTTGCCATGGCAATCTTCTGGAATT	6	254	3316123_1	99.0	.	DISC_MAPQ=46;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ACAATGATGTTATTAATAGGAATATGGATCAATTTCACAAAGAAGCCAATGAATCCCATTATAGCAAATCCTATTGCTGTTGCCATGGCAATCTTCTGGAATT;MAPQ=60;MATEID=3316123_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_54806501_54831501_329C;SPAN=5075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:256 DP:191 GQ:69.1 PL:[759.1, 69.1, 0.0] SR:254 DR:6 LR:-759.2 LO:759.2);ALT=A[chr7:54825188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	54820167	+	chr7	54826797	+	.	36	0	3316124_1	87.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=3316124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:54820167(+)-7:54826797(-)__7_54806501_54831501D;SPAN=6630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:116 GQ:87.5 PL:[87.5, 0.0, 193.1] SR:0 DR:36 LR:-87.41 LO:89.64);ALT=T[chr7:54826797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	54823619	+	chr7	54826848	+	.	59	0	3316134_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=3316134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:54823619(+)-7:54826848(-)__7_54806501_54831501D;SPAN=3229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:152 GQ:99 PL:[153.8, 0.0, 213.2] SR:0 DR:59 LR:-153.6 LO:154.1);ALT=T[chr7:54826848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	54825289	+	chr7	54826850	+	.	48	51	3316141_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=3316141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_54806501_54831501_32C;SPAN=1561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:88 DP:175 GQ:99 PL:[243.2, 0.0, 180.5] SR:51 DR:48 LR:-243.5 LO:243.5);ALT=T[chr7:54826850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
