chr5	29530256	+	chr5	29540078	+	.	104	0	3324096_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3324096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:29530256(+)-5:29540078(-)__5_29522501_29547501D;SPAN=9822;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:66 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:0 DR:104 LR:-307.0 LO:307.0);ALT=G[chr5:29540078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	29791146	+	chr5	29786795	+	.	8	0	3326351_1	0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=3326351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:29786795(-)-5:29791146(+)__5_29767501_29792501D;SPAN=4351;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:200 GQ:27.7 PL:[0.0, 27.7, 541.3] SR:0 DR:8 LR:27.78 LO:12.23);ALT=]chr5:29791146]T;VARTYPE=BND:DUP-th;JOINTYPE=th
