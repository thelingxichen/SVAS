chr1	2906067	+	chr1	2902382	+	.	12	0	18155_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=18155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:2902382(-)-1:2906067(+)__1_2891001_2916001D;SPAN=3685;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:12 DP:166 GQ:5.2 PL:[0.0, 5.2, 412.6] SR:0 DR:12 LR:5.362 LO:21.5);ALT=]chr1:2906067]A;VARTYPE=BND:DUP-th;JOINTYPE=th
