chr2	106879557	+	chr2	106885916	+	GCCCAG	70	59	1230114_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;INSERTION=GCCCAG;MAPQ=60;MATEID=1230114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_106869001_106894001_331C;SPAN=6359;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:116 DP:26 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:59 DR:70 LR:-343.3 LO:343.3);ALT=C[chr2:106885916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
