chr3	66335967	+	chrX	97207823	-	.	16	0	2078974_1	29.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2078974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:66335967(+)-23:97207823(+)__3_66321501_66346501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:85 GQ:29.9 PL:[29.9, 0.0, 175.1] SR:0 DR:16 LR:-29.79 LO:35.79);ALT=T]chrX:97207823];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chrX	96698346	+	chrX	96648234	+	.	8	0	11323494_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=11323494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:96648234(-)-23:96698346(+)__23_96677001_96702001D;SPAN=50112;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=]chrX:96698346]C;VARTYPE=BND:DUP-th;JOINTYPE=th
