chr5	136878453	+	chr5	136885592	+	.	15	0	3784249_1	36.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=3784249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:136878453(+)-5:136885592(-)__5_136857001_136882001D;SPAN=7139;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:49 GQ:36.2 PL:[36.2, 0.0, 82.4] SR:0 DR:15 LR:-36.24 LO:37.24);ALT=A[chr5:136885592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	136885828	+	chr5	136878802	+	.	20	0	3784251_1	54.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=3784251_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:136878802(-)-5:136885828(+)__5_136857001_136882001D;SPAN=7026;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:42 GQ:44.9 PL:[54.8, 0.0, 44.9] SR:0 DR:20 LR:-54.67 LO:54.67);ALT=]chr5:136885828]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	137022578	+	chr5	137023887	+	.	121	89	3784462_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAATATTACCTCCCT;MAPQ=60;MATEID=3784462_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_137004001_137029001_257C;SPAN=1309;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:172 DP:36 GQ:46.3 PL:[508.3, 46.3, 0.0] SR:89 DR:121 LR:-508.3 LO:508.3);ALT=T[chr5:137023887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
