chr3	50759282	+	chr3	50761229	-	.	9	0	2012750_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2012750_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:50759282(+)-3:50761229(+)__3_50739501_50764501D;SPAN=1947;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:136 GQ:6.9 PL:[0.0, 6.9, 343.2] SR:0 DR:9 LR:7.137 LO:15.77);ALT=C]chr3:50761229];VARTYPE=BND:INV-hh;JOINTYPE=hh
