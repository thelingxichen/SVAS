chr21	9660775	+	chr1	143130551	+	.	28	0	10691312_1	52.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=10691312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:143130551(-)-21:9660775(+)__21_9653001_9678001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:28 DP:148 GQ:52.4 PL:[52.4, 0.0, 306.5] SR:0 DR:28 LR:-52.33 LO:62.7);ALT=]chr21:9660775]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	143130729	+	chr21	9661434	+	.	16	0	10691313_1	9.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=10691313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:143130729(+)-21:9661434(-)__21_9653001_9678001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:162 GQ:9.1 PL:[9.1, 0.0, 382.1] SR:0 DR:16 LR:-8.926 LO:30.93);ALT=C[chr21:9661434[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
