chr1	98348932	+	chr1	98386440	+	.	0	8	247869_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=247869_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_98343001_98368001_71C;SPAN=37508;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:8 DR:0 LR:-19.36 LO:19.88);ALT=T[chr1:98386440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
