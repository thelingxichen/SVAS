chr9	113024576	+	chr9	113037094	+	TTATTATTATTAT	18	31	5962308_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TTATTATTATTAT;MAPQ=60;MATEID=5962308_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_113018501_113043501_55C;SPAN=12518;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:42 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:31 DR:18 LR:-125.4 LO:125.4);ALT=T[chr9:113037094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	113037287	+	chr9	113029970	+	.	73	61	5962313_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=5962313_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_113018501_113043501_89C;SPAN=7317;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:115 DP:56 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:61 DR:73 LR:-340.0 LO:340.0);ALT=]chr9:113037287]A;VARTYPE=BND:DUP-th;JOINTYPE=th
