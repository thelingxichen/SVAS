chr4	91084269	+	chr4	91148917	+	CCATGCTTA	0	40	2785020_1	99.0	.	EVDNC=ASSMB;INSERTION=CCATGCTTA;MAPQ=60;MATEID=2785020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_91066501_91091501_175C;SPAN=64648;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:40 DP:8 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:40 DR:0 LR:-118.8 LO:118.8);ALT=A[chr4:91148917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	91596798	+	chr4	91602909	+	.	72	42	2785825_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTGTTTTTATCTT;MAPQ=60;MATEID=2785825_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_4_91581001_91606001_212C;SPAN=6111;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:36 GQ:24 PL:[264.0, 24.0, 0.0] SR:42 DR:72 LR:-264.1 LO:264.1);ALT=T[chr4:91602909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
