chr11	76139879	+	chr2	63328429	-	.	64	0	10273828_1	99.0	.	BX=AAGTCACAGAATTCCC-1_1,GAGGTGACACCGCTAG-1_1,AGTCGATTCTGCTAGA-1_1,ACTACAGCATCCCTTG-1_1,GTCATTTGTGTGTTCA-1_1,CATCAAGTCGCAAGCC-1_1,GACACATGTGAGGGTT-1_1,TTAGTTCTCTGAAGCT-1_1,GCCAAATAGCCCGAAA-1_1,CTGGCGATCAATCGAC-1_1,CCTAACCTCCTATGAG-1_1,ATATTCCCAGTGAATA-1_1,GACCAATAGGTGCTTT-1_2,TGGCATAAGATTCACC-1_2,CTCTTAACAGGTCCCA-1_3,TTGAGCACATTCGTTT-1_1,CGTTAGAAGCAATTGA-1_1,TTGACTTTCCGTAGGC-1_1,CGGAACCTCATAAGCC-1_1,TCCGGAGCATCCTTGC-1_1,GCTATAGTCCGTTAAG-1_1,TACCCACCAATAAGCA-1_1,ACTCAGAAGTGGACGT-1_1,AGCTGGCAGCAGTAGC-1_1,CGTGAGCTCACTACAG-1_1,CAAAGCTCACTTACGA-1_1,GTCACCTCATTCCTCG-1_1,TATTACCTCCAGAAGG-1_1,AGCGGTCCATGTAGAA-1_1,TTTGTGTAGGAATCAT-1_1,TACAAGCAGGTAACGC-1_3,CCAGTGGAGAGTAAGG-1_1,ATTTCTGTCCAACCGG-1_1,GCCGGATAGATTGAGT-1_2,ACTAAGCGTTTGACAC-1_1,GTCGTGGTCGCTTGAA-1_1,CTCTTAAAGCCCGTTG-1_1,GTTAAGCCAGACAGGT-1_2,ACATGTGGTTGAGGTG-1_1,CTATGAGAGGTATCAA-1_1,GTTGCCTTCCACTCGT-1_1,TCGGGCAAGAAGTGCC-1_2,AGGGCAATCCTCTACG-1_1,CCGGGATCACGCTTTC-1_1,CTCGAAACAGACACGA-1_1,AGCAATCAGAGGGTTC-1_1,GGGTCTGCAGATCACT-1_1,ACGCTCTAGTTCTGTG-1_3,CAGGTATTCCGACGTG-1_1,CACATTTGTGAGCACA-1_1,ATCACCCTCTCCACTG-1_1,CGGTGTGTCTGTGCAA-1_1;DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=10273828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63328429(+)-11:76139879(+)__11_76121501_76146501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:31 GQ:8.4 PL:[0.0, 8.4, 92.4] SR:0 DR:0 LR:8.71 LO:0.0),OC001T.bam(GT:0/1 AD:64 DP:81 GQ:13.7 PL:[188.6, 0.0, 13.7] SR:0 DR:64 LR:-197.2 LO:197.2);ALT=t]chr11:76139879];VARTYPE=BND:TRX-tt;JOINTYPE=tt	.
chr11	76139879	+	chr2	63328429	-	.	64	0	10273828_1	99.0	.	BX=AAGTCACAGAATTCCC-1_1,GAGGTGACACCGCTAG-1_1,AGTCGATTCTGCTAGA-1_1,ACTACAGCATCCCTTG-1_1,GTCATTTGTGTGTTCA-1_1,CATCAAGTCGCAAGCC-1_1,GACACATGTGAGGGTT-1_1,TTAGTTCTCTGAAGCT-1_1,GCCAAATAGCCCGAAA-1_1,CTGGCGATCAATCGAC-1_1,CCTAACCTCCTATGAG-1_1,ATATTCCCAGTGAATA-1_1,GACCAATAGGTGCTTT-1_2,TGGCATAAGATTCACC-1_2,CTCTTAACAGGTCCCA-1_3,TTGAGCACATTCGTTT-1_1,CGTTAGAAGCAATTGA-1_1,TTGACTTTCCGTAGGC-1_1,CGGAACCTCATAAGCC-1_1,TCCGGAGCATCCTTGC-1_1,GCTATAGTCCGTTAAG-1_1,TACCCACCAATAAGCA-1_1,ACTCAGAAGTGGACGT-1_1,AGCTGGCAGCAGTAGC-1_1,CGTGAGCTCACTACAG-1_1,CAAAGCTCACTTACGA-1_1,GTCACCTCATTCCTCG-1_1,TATTACCTCCAGAAGG-1_1,AGCGGTCCATGTAGAA-1_1,TTTGTGTAGGAATCAT-1_1,TACAAGCAGGTAACGC-1_3,CCAGTGGAGAGTAAGG-1_1,ATTTCTGTCCAACCGG-1_1,GCCGGATAGATTGAGT-1_2,ACTAAGCGTTTGACAC-1_1,GTCGTGGTCGCTTGAA-1_1,CTCTTAAAGCCCGTTG-1_1,GTTAAGCCAGACAGGT-1_2,ACATGTGGTTGAGGTG-1_1,CTATGAGAGGTATCAA-1_1,GTTGCCTTCCACTCGT-1_1,TCGGGCAAGAAGTGCC-1_2,AGGGCAATCCTCTACG-1_1,CCGGGATCACGCTTTC-1_1,CTCGAAACAGACACGA-1_1,AGCAATCAGAGGGTTC-1_1,GGGTCTGCAGATCACT-1_1,ACGCTCTAGTTCTGTG-1_3,CAGGTATTCCGACGTG-1_1,CACATTTGTGAGCACA-1_1,ATCACCCTCTCCACTG-1_1,CGGTGTGTCTGTGCAA-1_1;DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=10273828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63328429(+)-11:76139879(+)__11_76121501_76146501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:31 GQ:8.4 PL:[0.0, 8.4, 92.4] SR:0 DR:0 LR:8.71 LO:0.0),OC001T.bam(GT:0/1 AD:64 DP:81 GQ:13.7 PL:[188.6, 0.0, 13.7] SR:0 DR:64 LR:-197.2 LO:197.2);ALT=t]chr11:76139879];VARTYPE=BND:TRX-tt;JOINTYPE=tt	.
