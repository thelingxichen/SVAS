chr10	51565329	+	chr10	51579126	+	.	13	0	4595101_1	34.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4595101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:51565329(+)-10:51579126(-)__10_51572501_51597501D;SPAN=13797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:32 GQ:34.4 PL:[34.4, 0.0, 41.0] SR:0 DR:13 LR:-34.24 LO:34.3);ALT=T[chr10:51579126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	51565341	+	chr10	51580553	+	.	16	0	4595102_1	44.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4595102_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:51565341(+)-10:51580553(-)__10_51572501_51597501D;SPAN=15212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:30 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:0 DR:16 LR:-44.89 LO:44.89);ALT=C[chr10:51580553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
