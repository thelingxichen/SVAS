chr5	15133086	+	chr10	93500789	+	GTGGGGGTCGTGGGGTCTCTTGCTGCCAGGATTCCAG	40	146	6438818_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=GTGGGGGTCGTGGGGTCTCTTGCTGCCAGGATTCCAG;MAPQ=60;MATEID=6438818_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_10_93492001_93517001_114C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:157 DP:77 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:146 DR:40 LR:-465.4 LO:465.4);ALT=C[chr10:93500789[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	93633338	+	chr10	93634563	+	.	0	112	6438681_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CAC;MAPQ=60;MATEID=6438681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_93614501_93639501_258C;SPAN=1225;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:112 DP:49 GQ:30 PL:[330.0, 30.0, 0.0] SR:112 DR:0 LR:-330.1 LO:330.1);ALT=C[chr10:93634563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	94134599	+	chr10	94137654	+	GTTGACTTATCTTTT	142	77	6441966_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;INSERTION=GTTGACTTATCTTTT;MAPQ=60;MATEID=6441966_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_94129001_94154001_419C;SPAN=3055;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:183 DP:88 GQ:49.3 PL:[541.3, 49.3, 0.0] SR:77 DR:142 LR:-541.3 LO:541.3);ALT=A[chr10:94137654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
