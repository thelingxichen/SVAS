chr1	40966776	+	chr1	40970572	+	.	75	59	206123_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGAT;MAPQ=60;MATEID=206123_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_40964001_40989001_376C;SPAN=3796;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:107 DP:116 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:59 DR:75 LR:-343.3 LO:343.3);ALT=T[chr1:40970572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
