chr1	146779562	-	chr9	1422881	+	.	15	0	515103_1	32.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=515103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146779562(-)-9:1422881(-)__1_146779501_146804501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:0 DR:15 LR:-32.72 LO:35.42);ALT=[chr9:1422881[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	147737793	+	chr4	64751670	-	.	35	16	520154_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=AGGAAGGAAGGAAGGAAGGAAGGAAGGAA;MAPQ=31;MATEID=520154_2;MATENM=1;NM=3;NUMPARTS=2;SCTG=c_1_147735001_147760001_249C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:50 DP:31 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:16 DR:35 LR:-148.5 LO:148.5);ALT=T]chr4:64751670];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	147752841	-	chr1	147775507	+	.	36	40	519603_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GCCTCTCAGGTTTTCCGAGGCTTTGGAGCCTGCACA;MAPQ=60;MATEID=519603_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_1_147759501_147784501_447C;SPAN=22666;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:76 DP:25 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:40 DR:36 LR:-224.5 LO:224.5);ALT=[chr1:147775507[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	109310554	+	chr2	109312123	+	TTCTGCTTGCC	58	37	1241599_1	99.0	.	DISC_MAPQ=34;EVDNC=ASDIS;INSERTION=TTCTGCTTGCC;MAPQ=0;MATEID=1241599_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=CGCG;SCTG=c_2_109294501_109319501_365C;SECONDARY;SPAN=1569;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:83 DP:113 GQ:29 PL:[243.5, 0.0, 29.0] SR:37 DR:58 LR:-252.9 LO:252.9);ALT=C[chr2:109312123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	109639512	+	chr9	817682	+	.	7	12	5763590_1	51.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=ACTCCAGCCTGGGCGACAGAGCGAGACTCCATCTCAAAAAA;MAPQ=43;MATEID=5763590_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_9_808501_833501_18C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:31 GQ:21.5 PL:[51.2, 0.0, 21.5] SR:12 DR:7 LR:-51.54 LO:51.54);ALT=A[chr9:817682[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	137072366	+	chr3	137073447	+	.	54	44	2349206_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAC;MAPQ=60;MATEID=2349206_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_137053001_137078001_331C;SPAN=1081;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:82 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:44 DR:54 LR:-241.0 LO:241.0);ALT=C[chr3:137073447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	2397101	+	chr3	137221712	+	CAGTACATCCCAAGTGGCTGAGCAGTAATCTTTTTTTTTTT	8	59	2349528_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;INSERTION=CAGTACATCCCAAGTGGCTGAGCAGTAATCTTTTTTTTTTT;MAPQ=21;MATEID=2349528_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_3_137200001_137225001_226C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:66 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:59 DR:8 LR:-194.7 LO:194.7);ALT=]chr9:2397101]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	138129860	+	chr11	43756679	+	.	8	0	6773584_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6773584_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_43732501_43757501_154C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:102 GQ:0.9 PL:[0.0, 0.9, 247.5] SR:0 DR:8 LR:1.226 LO:14.63);ALT=G[chr11:43756679[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	139318061	+	chr3	138920642	+	CAAGCTTTAAGTTTCTGT	28	32	2360102_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CAAGCTTTAAGTTTCTGT;MAPQ=60;MATEID=2360102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_139307001_139332001_366C;SPAN=397419;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:63 GQ:2.9 PL:[148.1, 0.0, 2.9] SR:32 DR:28 LR:-156.1 LO:156.1);ALT=]chr3:139318061]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	65719085	+	chr4	65721141	-	.	5	50	2738108_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=TGT;MAPQ=60;MATEID=2738108_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_65709001_65734001_167C;SPAN=2056;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:52 DP:50 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:50 DR:5 LR:-151.8 LO:151.8);ALT=A]chr4:65721141];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	65719561	-	chr4	65721074	+	CTGGTGTGAACCCGGGAGGCGGAGCTATCTG	17	72	2738111_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGGTGTGAACCCGGGAGGCGGAGCTATCTG;MAPQ=60;MATEID=2738111_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_65709001_65734001_69C;SPAN=1513;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:66 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:72 DR:17 LR:-234.4 LO:234.4);ALT=[chr4:65721074[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	4190435	+	chr9	3107626	+	.	33	25	5769611_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=CGATCAACTGGAAGAAAGGGTATCAGTGA;MAPQ=60;MATEID=5769611_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_4189501_4214501_17C;SPAN=1082809;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:49 DP:20 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:25 DR:33 LR:-145.2 LO:145.2);ALT=]chr9:4190435]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	3107812	+	chr9	4190646	+	.	11	0	5769612_1	26.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5769612_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:3107812(+)-9:4190646(-)__9_4189501_4214501D;SPAN=1082834;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:0 DR:11 LR:-26.29 LO:27.14);ALT=G[chr9:4190646[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
