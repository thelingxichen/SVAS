chr8	141467775	+	chr8	141446090	+	.	5	4	5739447_1	18.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=5739447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_141463001_141488001_252C;SPAN=21685;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:4 DR:5 LR:-18.82 LO:19.57);ALT=]chr8:141467775]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	142089039	+	chr8	141958591	+	AAC	61	20	5741812_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AAC;MAPQ=60;MATEID=5741812_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_141953001_141978001_38C;SPAN=130448;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:79 GQ:8.1 PL:[207.9, 8.1, 0.0] SR:20 DR:61 LR:-214.3 LO:214.3);ALT=]chr8:142089039]A;VARTYPE=BND:DUP-th;JOINTYPE=th
