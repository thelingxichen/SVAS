chr6	24325366	+	chr6	24327808	+	.	145	75	4081924_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TCTCC;MAPQ=60;MATEID=4081924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24304001_24329001_20C;SPAN=2442;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:187 DP:25 GQ:50.5 PL:[554.5, 50.5, 0.0] SR:75 DR:145 LR:-554.5 LO:554.5);ALT=C[chr6:24327808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24811887	+	chr6	24817951	+	.	103	99	4084294_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CGTTTAGTACTT;MAPQ=60;MATEID=4084294_2;MATENM=13;NM=3;NUMPARTS=2;SCTG=c_6_24794001_24819001_389C;SPAN=6064;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:170 DP:45 GQ:46 PL:[505.0, 46.0, 0.0] SR:99 DR:103 LR:-505.0 LO:505.0);ALT=T[chr6:24817951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
