chr13	78997624	+	chr13	78998720	+	.	58	32	8171526_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AACATGGTGAAACCC;MAPQ=60;MATEID=8171526_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_78988001_79013001_361C;SPAN=1096;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:87 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:32 DR:58 LR:-256.6 LO:256.6);ALT=C[chr13:78998720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
