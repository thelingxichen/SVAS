chr10	114112183	+	chr10	114116659	+	.	122	112	6529653_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6529653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_114096501_114121501_10C;SPAN=4476;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:198 DP:42 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:112 DR:122 LR:-587.5 LO:587.5);ALT=G[chr10:114116659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
