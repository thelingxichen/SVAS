chr12	75107858	+	chr12	75110750	-	.	42	68	7754631_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=7754631_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75092501_75117501_326C;SPAN=2892;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:95 DP:218 GQ:99 PL:[254.6, 0.0, 274.4] SR:68 DR:42 LR:-254.5 LO:254.6);ALT=A]chr12:75110750];VARTYPE=BND:INV-hh;JOINTYPE=hh
