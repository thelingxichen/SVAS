chr14	80106290	+	chr14	80115050	+	.	60	44	8630786_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=8630786_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_80115001_80140001_123C;SPAN=8760;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:39 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:44 DR:60 LR:-260.8 LO:260.8);ALT=G[chr14:80115050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
