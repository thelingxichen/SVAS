chr7	155471378	+	chr7	155473282	+	.	5	3	3701290_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3701290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_155452501_155477501_137C;SPAN=1904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:60 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:3 DR:5 LR:-6.852 LO:14.07);ALT=G[chr7:155473282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
