chrX	16876973	+	chrX	16881078	+	.	3	3	7372564_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7372564_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_16880501_16905501_43C;SPAN=4105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:30 GQ:8.3 PL:[8.3, 0.0, 64.4] SR:3 DR:3 LR:-8.377 LO:10.89);ALT=C[chrX:16881078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
