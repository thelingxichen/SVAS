chr1	198773749	+	chr1	198775415	+	.	0	55	741122_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=741122_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_198768501_198793501_381C;SPAN=1666;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:85 GQ:46.4 PL:[158.6, 0.0, 46.4] SR:55 DR:0 LR:-161.8 LO:161.8);ALT=T[chr1:198775415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	199438743	+	chr1	199440234	+	.	128	54	743821_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAATATTGGGTCTCA;MAPQ=60;MATEID=743821_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_199430001_199455001_309C;SPAN=1491;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:166 DP:201 GQ:7.9 PL:[501.7, 7.9, 0.0] SR:54 DR:128 LR:-525.6 LO:525.6);ALT=A[chr1:199440234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	199530641	-	chr1	199531851	+	.	12	0	743696_1	14.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=743696_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:199530641(-)-1:199531851(-)__1_199528001_199553001D;SPAN=1210;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:92 GQ:14.9 PL:[14.9, 0.0, 206.3] SR:0 DR:12 LR:-14.69 LO:24.74);ALT=[chr1:199531851[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
