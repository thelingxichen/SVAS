chrX	110924572	+	chrX	110928189	+	.	9	0	7497856_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7497856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:110924572(+)-23:110928189(-)__23_110911501_110936501D;SPAN=3617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:0 DR:9 LR:-11.83 LO:18.75);ALT=C[chrX:110928189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	110925524	+	chrX	110928191	+	.	0	7	7497858_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=7497858_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_110911501_110936501_39C;SPAN=2667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:52 GQ:9.2 PL:[9.2, 0.0, 114.8] SR:7 DR:0 LR:-9.019 LO:14.54);ALT=T[chrX:110928191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
