chrX	15056111	+	chrX	15024945	+	TGTAA	0	64	10986410_1	99.0	.	EVDNC=ASSMB;INSERTION=TGTAA;MAPQ=60;MATEID=10986410_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_15043001_15068001_362C;SPAN=31166;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:96 GQ:46.7 PL:[185.3, 0.0, 46.7] SR:64 DR:0 LR:-189.8 LO:189.8);ALT=]chrX:15056111]A;VARTYPE=BND:DUP-th;JOINTYPE=th
