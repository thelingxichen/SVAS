chr2	109310554	+	chr2	109312110	+	.	52	48	935930_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=C;MAPQ=0;MATEID=935930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_109294501_109319501_75C;SPAN=1556;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:53 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:48 DR:52 LR:-244.3 LO:244.3);ALT=C[chr2:109312110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
