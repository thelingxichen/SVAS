chr8	15289364	+	chr13	74314062	-	.	34	60	8153371_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TATGTT;MAPQ=60;MATEID=8153371_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_74308501_74333501_186C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:85 DP:72 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:60 DR:34 LR:-250.9 LO:250.9);ALT=T]chr13:74314062];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	15289367	-	chr13	74313858	+	.	47	67	8153373_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCCA;MAPQ=60;MATEID=8153373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_74308501_74333501_65C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:102 DP:68 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:67 DR:47 LR:-300.4 LO:300.4);ALT=[chr13:74313858[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
