chr12	19508861	-	chr12	19510192	+	.	10	0	5114674_1	10.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5114674_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:19508861(-)-12:19510192(-)__12_19502001_19527001D;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:0 DR:10 LR:-10.52 LO:20.25);ALT=[chr12:19510192[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
