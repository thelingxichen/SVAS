chr3	148281440	+	chr3	148285420	+	.	49	47	2394860_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=GTCCTG;MAPQ=60;MATEID=2394860_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148274001_148299001_378C;SPAN=3980;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:86 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:47 DR:49 LR:-254.2 LO:254.2);ALT=G[chr3:148285420[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
