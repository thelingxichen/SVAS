chr9	75766840	+	chr9	75773436	+	.	131	27	4273448_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4273448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_75754001_75779001_178C;SPAN=6596;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:150 DP:287 GQ:99 PL:[417.5, 0.0, 278.8] SR:27 DR:131 LR:-418.9 LO:418.9);ALT=G[chr9:75773436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75766868	+	chr9	75773668	+	.	31	0	4273450_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75766868(+)-9:75773668(-)__9_75754001_75779001D;SPAN=6800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:272 GQ:28.9 PL:[28.9, 0.0, 629.6] SR:0 DR:31 LR:-28.64 LO:61.98);ALT=T[chr9:75773668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75775317	+	chr9	75777696	+	.	9	0	4273487_1	1.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4273487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75775317(+)-9:75777696(-)__9_75754001_75779001D;SPAN=2379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:106 GQ:1.1 PL:[1.1, 0.0, 255.2] SR:0 DR:9 LR:-0.991 LO:16.78);ALT=T[chr9:75777696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75775325	+	chr9	75778389	+	.	9	0	4273488_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75775325(+)-9:75778389(-)__9_75754001_75779001D;SPAN=3064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:0 DR:9 LR:-0.7201 LO:16.74);ALT=T[chr9:75778389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75775809	+	chr9	75780031	+	AACTGAAGAGAGATCTGGCCAAAGACATAACCTCAGACACATCTGGAGATTTTCGGAACGCTTTGCTTTCTCTTGCTAAGGGTGACCGATCTGAGGACTTTGGTGTGAATGAAGACTTGGCTGATTCAGATGCCAG	9	56	4273714_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AACTGAAGAGAGATCTGGCCAAAGACATAACCTCAGACACATCTGGAGATTTTCGGAACGCTTTGCTTTCTCTTGCTAAGGGTGACCGATCTGAGGACTTTGGTGTGAATGAAGACTTGGCTGATTCAGATGCCAG;MAPQ=60;MATEID=4273714_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_9_75778501_75803501_170C;SPAN=4222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:72 GQ:0.5 PL:[172.1, 0.0, 0.5] SR:56 DR:9 LR:-182.0 LO:182.0);ALT=G[chr9:75780031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75775809	+	chr9	75777697	+	.	5	26	4273490_1	65.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4273490_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_9_75754001_75779001_65C;SPAN=1888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:113 GQ:65.3 PL:[65.3, 0.0, 207.2] SR:26 DR:5 LR:-65.12 LO:69.34);ALT=G[chr9:75777697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75775853	+	chr9	75778389	+	.	13	0	4273492_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75775853(+)-9:75778389(-)__9_75754001_75779001D;SPAN=2536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:97 GQ:16.7 PL:[16.7, 0.0, 218.0] SR:0 DR:13 LR:-16.63 LO:26.97);ALT=G[chr9:75778389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75777807	+	chr9	75780030	+	.	22	0	4273716_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75777807(+)-9:75780030(-)__9_75778501_75803501D;SPAN=2223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:71 GQ:53.6 PL:[53.6, 0.0, 116.3] SR:0 DR:22 LR:-53.39 LO:54.76);ALT=C[chr9:75780030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75777821	+	chr9	75781010	+	.	8	0	4273717_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75777821(+)-9:75781010(-)__9_75778501_75803501D;SPAN=3189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:0 DR:8 LR:0.9554 LO:14.66);ALT=A[chr9:75781010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75778449	+	chr9	75780031	+	.	9	41	4273719_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4273719_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GGG;SCTG=c_9_75778501_75803501_170C;SPAN=1582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:92 GQ:84.2 PL:[137.0, 0.0, 84.2] SR:41 DR:9 LR:-137.4 LO:137.4);ALT=G[chr9:75780031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75780172	+	chr9	75783947	+	.	9	0	4273725_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273725_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75780172(+)-9:75783947(-)__9_75778501_75803501D;SPAN=3775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:157 GQ:12.7 PL:[0.0, 12.7, 405.9] SR:0 DR:9 LR:12.83 LO:15.19);ALT=T[chr9:75783947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75781108	+	chr9	75783948	+	TGAAGTGCGCCACAAGCAAACCAGCTTTCTTTGCAGAGAAGCTTCATCAAGCCATGAAA	23	45	4273734_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TGAAGTGCGCCACAAGCAAACCAGCTTTCTTTGCAGAGAAGCTTCATCAAGCCATGAAA;MAPQ=60;MATEID=4273734_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_75778501_75803501_194C;SPAN=2840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:148 GQ:99 PL:[151.4, 0.0, 207.5] SR:45 DR:23 LR:-151.4 LO:151.8);ALT=G[chr9:75783948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75781108	+	chr9	75782412	+	.	4	16	4273733_1	23.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4273733_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_75778501_75803501_194C;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:134 GQ:23.3 PL:[23.3, 0.0, 300.5] SR:16 DR:4 LR:-23.11 LO:37.37);ALT=G[chr9:75782412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75782472	+	chr9	75783948	+	.	7	33	4273741_1	95.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4273741_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_75778501_75803501_194C;SPAN=1476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:134 GQ:95.9 PL:[95.9, 0.0, 227.9] SR:33 DR:7 LR:-95.74 LO:98.77);ALT=G[chr9:75783948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	75782518	+	chr9	75784965	+	.	18	0	4273742_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4273742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:75782518(+)-9:75784965(-)__9_75778501_75803501D;SPAN=2447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:109 GQ:29.9 PL:[29.9, 0.0, 234.5] SR:0 DR:18 LR:-29.89 LO:39.13);ALT=T[chr9:75784965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
