chr14	21952624	+	chr14	21954663	+	T	56	33	8379267_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=8379267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_21952001_21977001_80C;SPAN=2039;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:73 DP:88 GQ:3.9 PL:[221.1, 3.9, 0.0] SR:33 DR:56 LR:-231.5 LO:231.5);ALT=C[chr14:21954663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
