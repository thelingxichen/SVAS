chr10	45455314	+	chr10	45465612	+	.	4	2	4584960_1	0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4584960_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_10_45447501_45472501_15C;SPAN=10298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:58 GQ:2.4 PL:[0.0, 2.4, 145.2] SR:2 DR:4 LR:2.51 LO:7.082);ALT=G[chr10:45465612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	45455335	+	chr10	45477966	+	.	8	0	4585031_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4585031_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:45455335(+)-10:45477966(-)__10_45472001_45497001D;SPAN=22631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=A[chr10:45477966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	45467297	+	chr10	45477967	+	.	0	9	4584980_1	22.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4584980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_45447501_45472501_240C;SPAN=10670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:9 DR:0 LR:-22.39 LO:22.75);ALT=G[chr10:45477967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	45496468	+	chr10	45498726	+	.	77	0	4585275_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4585275_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:45496468(+)-10:45498726(-)__10_45496501_45521501D;SPAN=2258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:35 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:0 DR:77 LR:-227.8 LO:227.8);ALT=C[chr10:45498726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	45869880	+	chr10	45877930	+	.	21	22	4585631_1	95.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=GGTG;MAPQ=60;MATEID=4585631_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_45864001_45889001_209C;SPAN=8050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:52 GQ:29 PL:[95.0, 0.0, 29.0] SR:22 DR:21 LR:-96.6 LO:96.6);ALT=G[chr10:45877930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
