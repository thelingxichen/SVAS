chr4	42762678	+	chr4	42769543	+	.	20	20	1951197_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1951197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_42752501_42777501_91C;SPAN=6865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:32 GQ:9 PL:[99.0, 9.0, 0.0] SR:20 DR:20 LR:-99.02 LO:99.02);ALT=G[chr4:42769543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
