chr16	46958953	+	chr16	46960105	-	.	8	0	9294463_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=9294463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:46958953(+)-16:46960105(+)__16_46942001_46967001D;SPAN=1152;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:142 GQ:11.7 PL:[0.0, 11.7, 366.3] SR:0 DR:8 LR:12.06 LO:13.44);ALT=C]chr16:46960105];VARTYPE=BND:INV-hh;JOINTYPE=hh
