chr16	14014230	+	chr16	14015886	+	.	0	7	6118871_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6118871_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_13989501_14014501_38C;SPAN=1656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:40 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:7 DR:0 LR:-12.27 LO:15.41);ALT=G[chr16:14015886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	14721195	+	chr16	14723453	+	TTTTAAGCTTCTGATACCTCTCTTCTGGAGTGTCAAAACCATTTGTTAATGCAGAGACTGAAGGTCCATCACTGATT	0	12	6121205_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TTTTAAGCTTCTGATACCTCTCTTCTGGAGTGTCAAAACCATTTGTTAATGCAGAGACTGAAGGTCCATCACTGATT;MAPQ=60;MATEID=6121205_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_14700001_14725001_219C;SPAN=2258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:12 DR:0 LR:-16.31 LO:25.12);ALT=T[chr16:14723453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	14726901	+	chr16	14738129	+	.	36	0	6121293_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6121293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:14726901(+)-16:14738129(-)__16_14724501_14749501D;SPAN=11228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:96 GQ:92.9 PL:[92.9, 0.0, 139.1] SR:0 DR:36 LR:-92.83 LO:93.35);ALT=G[chr16:14738129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15141958	+	chr16	15149747	+	.	8	3	6122986_1	12.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6122986_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_15141001_15166001_410C;SPAN=7789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:3 DR:8 LR:-12.69 LO:20.72);ALT=T[chr16:15149747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15744200	+	chr16	15761140	+	.	21	0	6126363_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6126363_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:15744200(+)-16:15761140(-)__16_15753501_15778501D;SPAN=16940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:41 GQ:38.6 PL:[58.4, 0.0, 38.6] SR:0 DR:21 LR:-58.37 LO:58.37);ALT=C[chr16:15761140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15744203	+	chr16	15758590	+	.	12	0	6126364_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6126364_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:15744203(+)-16:15758590(-)__16_15753501_15778501D;SPAN=14387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=C[chr16:15758590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15758719	+	chr16	15761141	+	.	0	17	6126389_1	33.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6126389_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_15753501_15778501_55C;SPAN=2422;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:17 DR:0 LR:-33.63 LO:38.73);ALT=G[chr16:15761141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15961374	+	chr16	15967348	+	.	0	7	6127074_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6127074_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_15949501_15974501_32C;SPAN=5974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=C[chr16:15967348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15973748	+	chr16	15977865	+	.	0	14	6127228_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6127228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_15974001_15999001_204C;SPAN=4117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:41 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:14 DR:0 LR:-35.11 LO:35.58);ALT=G[chr16:15977865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	15978073	+	chr16	15982413	+	.	23	0	6127242_1	48.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6127242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:15978073(+)-16:15982413(-)__16_15974001_15999001D;SPAN=4340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:103 GQ:48.2 PL:[48.2, 0.0, 200.0] SR:0 DR:23 LR:-48.02 LO:53.38);ALT=T[chr16:15982413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
