chr14	37769602	+	chr16	61079339	-	.	18	0	6226767_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6226767_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:37769602(+)-16:61079339(+)__16_61078501_61103501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:29 GQ:18.5 PL:[51.5, 0.0, 18.5] SR:0 DR:18 LR:-52.4 LO:52.4);ALT=A]chr16:61079339];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr16	60910045	+	chr16	60913925	+	.	0	24	6226414_1	75.0	.	EVDNC=ASSMB;HOMSEQ=AAAAAAAAA;MAPQ=60;MATEID=6226414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_60907001_60932001_240C;SPAN=3880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:28 GQ:4.2 PL:[75.9, 4.2, 0.0] SR:24 DR:0 LR:-77.12 LO:77.12);ALT=A[chr16:60913925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
