chr14	105925443	+	chr14	105926486	+	.	9	0	8738726_1	10.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=8738726_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105925443(+)-14:105926486(-)__14_105913501_105938501D;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=C[chr14:105926486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106449027	+	chr14	106450849	+	.	101	39	8742437_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;MAPQ=60;MATEID=8742437_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106428001_106453001_69C;SPAN=1822;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:124 DP:87 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:39 DR:101 LR:-366.4 LO:366.4);ALT=T[chr14:106450849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106572849	+	chr14	106518045	+	.	20	0	8742652_1	50.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=8742652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106518045(-)-14:106572849(+)__14_106550501_106575501D;SPAN=54804;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:56 GQ:50.9 PL:[50.9, 0.0, 83.9] SR:0 DR:20 LR:-50.85 LO:51.32);ALT=]chr14:106572849]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106518239	+	chr14	106573325	+	.	10	0	8742653_1	19.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=8742653_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106518239(+)-14:106573325(-)__14_106550501_106575501D;SPAN=55086;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:52 GQ:19.1 PL:[19.1, 0.0, 104.9] SR:0 DR:10 LR:-18.92 LO:22.47);ALT=G[chr14:106573325[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106550908	+	chr14	106924658	+	.	8	0	8744692_1	4.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=8744692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106550908(+)-14:106924658(-)__14_106918001_106943001D;SPAN=373750;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=T[chr14:106924658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106650013	+	chr14	106841681	+	.	24	0	8742863_1	64.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=8742863_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106650013(+)-14:106841681(-)__14_106648501_106673501D;SPAN=191668;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:55 GQ:64.4 PL:[64.4, 0.0, 67.7] SR:0 DR:24 LR:-64.32 LO:64.33);ALT=A[chr14:106841681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106842070	+	chr14	106650352	+	.	43	0	8742867_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=8742867_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106650352(-)-14:106842070(+)__14_106648501_106673501D;SPAN=191718;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:43 DP:22 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=]chr14:106842070]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106712928	+	chr14	107011400	+	.	15	0	8743152_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=8743152_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106712928(+)-14:107011400(-)__14_106697501_106722501D;SPAN=298472;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:50 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.97 LO:37.08);ALT=T[chr14:107011400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	107011599	+	chr14	106713056	+	.	10	0	8743153_1	19.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ATCCCGAGGAGATGGCCTAATCCAAGGAGAGGGAGGCTCCAGGTCGTGTGGACTCACACGGGGCTCCTCCTTCTGCCC;MAPQ=0;MATEID=8743153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106697501_106722501_293C;SECONDARY;SPAN=298543;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:52 GQ:19.1 PL:[19.1, 0.0, 104.9] SR:0 DR:10 LR:-18.92 LO:22.47);ALT=]chr14:107011599]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	107273723	+	chr14	107093606	+	CGTGTGC	20	53	8746711_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CGTGTGC;MAPQ=60;MATEID=8746711_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_14_107089501_107114501_123C;SPAN=180117;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:64 DP:60 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:53 DR:20 LR:-188.1 LO:188.1);ALT=]chr14:107273723]C;VARTYPE=BND:DUP-th;JOINTYPE=th
