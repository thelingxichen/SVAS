chr8	5728020	+	chr8	5729354	+	AAAA	0	63	5375952_1	99.0	.	EVDNC=ASSMB;INSERTION=AAAA;MAPQ=60;MATEID=5375952_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_5708501_5733501_227C;SPAN=1334;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:25 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:63 DR:0 LR:-184.8 LO:184.8);ALT=A[chr8:5729354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
