chr5	160680743	+	chr5	160671899	+	.	24	0	3886950_1	48.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3886950_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:160671899(-)-5:160680743(+)__5_160671001_160696001D;SPAN=8844;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:113 GQ:48.8 PL:[48.8, 0.0, 223.7] SR:0 DR:24 LR:-48.61 LO:55.1);ALT=]chr5:160680743]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	160672106	+	chr5	160681111	+	.	8	0	3886951_1	0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=3886951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:160672106(+)-5:160681111(-)__5_160671001_160696001D;SPAN=9005;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:144 GQ:12.3 PL:[0.0, 12.3, 372.9] SR:0 DR:8 LR:12.61 LO:13.39);ALT=C[chr5:160681111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
