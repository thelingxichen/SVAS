chr11	69663331	+	chr19	29642735	-	.	11	0	6892554_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6892554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:69663331(+)-19:29642735(+)__11_69653501_69678501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=T]chr19:29642735];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr19	29950197	+	chr19	29956168	+	.	46	42	10241401_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAGAAATTA;MAPQ=60;MATEID=10241401_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_29939001_29964001_395C;SPAN=5971;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:86 GQ:6.5 PL:[201.2, 0.0, 6.5] SR:42 DR:46 LR:-212.0 LO:212.0);ALT=A[chr19:29956168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	30388804	+	chr19	30393101	+	.	55	36	10243316_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAATTTTTATTTTT;MAPQ=60;MATEID=10243316_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_30380001_30405001_144C;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:118 GQ:70.4 PL:[215.6, 0.0, 70.4] SR:36 DR:55 LR:-219.6 LO:219.6);ALT=T[chr19:30393101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	31298214	+	chr19	31308630	+	.	0	55	10246967_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=10246967_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_31286501_31311501_266C;SPAN=10416;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:55 DP:75 GQ:19.4 PL:[161.3, 0.0, 19.4] SR:55 DR:0 LR:-167.5 LO:167.5);ALT=C[chr19:31308630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
