chr5	42028778	+	chr5	42027701	+	.	4	2	3394223_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCTTGCTTTT;MAPQ=60;MATEID=3394223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_42017501_42042501_62C;SPAN=1077;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:135 GQ:23.1 PL:[0.0, 23.1, 372.9] SR:2 DR:4 LR:23.37 LO:5.59);ALT=]chr5:42028778]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	42165941	+	chr5	42167770	+	.	110	84	3394834_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTAAAACTTTGTT;MAPQ=60;MATEID=3394834_2;MATENM=4;NM=4;NUMPARTS=2;SCTG=c_5_42164501_42189501_55C;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:157 DP:28 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:84 DR:110 LR:-465.4 LO:465.4);ALT=T[chr5:42167770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
