chr2	204566581	+	chr2	204567748	-	.	4	2	1634719_1	0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AGCTTCTGCACAGCAAAAGAAAC;MAPQ=60;MATEID=1634719_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_204550501_204575501_205C;SPAN=1167;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:124 GQ:16.8 PL:[0.0, 16.8, 333.3] SR:2 DR:4 LR:17.09 LO:7.662);ALT=C]chr2:204567748];VARTYPE=BND:INV-hh;JOINTYPE=hh
