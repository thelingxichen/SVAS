chr11	51341203	+	chr11	51362970	+	.	65	28	4862357_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GTTTAACTCTGTGAGATGAATGCACACATCACAAAGC;MAPQ=60;MATEID=4862357_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_11_51327501_51352501_201C;SPAN=21767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:6 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:28 DR:65 LR:-260.8 LO:260.8);ALT=C[chr11:51362970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
