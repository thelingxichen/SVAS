chr1	194451080	+	chr1	194454312	+	.	8	0	724968_1	22.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=724968_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:194451080(+)-1:194454312(-)__1_194432001_194457001D;SPAN=3232;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:14 GQ:9.5 PL:[22.7, 0.0, 9.5] SR:0 DR:8 LR:-22.82 LO:22.82);ALT=A[chr1:194454312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
