chr4	175625169	+	chr4	175626971	+	.	67	42	3082656_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGG;MAPQ=60;MATEID=3082656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_175616001_175641001_128C;SPAN=1802;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:68 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:42 DR:67 LR:-277.3 LO:277.3);ALT=G[chr4:175626971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
