chr1	62175110	+	chr1	62189385	+	.	0	12	175456_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=175456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_62181001_62206001_10C;SPAN=14275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:38 GQ:29.3 PL:[29.3, 0.0, 62.3] SR:12 DR:0 LR:-29.32 LO:29.99);ALT=C[chr1:62189385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	62189458	+	chr1	62190625	+	.	0	9	175496_1	8.0	.	EVDNC=ASSMB;HOMSEQ=ATAT;MAPQ=60;MATEID=175496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_62181001_62206001_137C;SPAN=1167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-7.764 LO:17.89);ALT=T[chr1:62190625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	62903071	+	chr1	62905467	+	.	5	6	177451_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=177451_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_62891501_62916501_302C;SPAN=2396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:6 DR:5 LR:-10.97 LO:16.77);ALT=G[chr1:62905467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
