chr12	82139719	+	chr12	82144320	+	.	74	62	7775359_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AACA;MAPQ=60;MATEID=7775359_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_12_82124001_82149001_128C;SPAN=4601;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:21 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:62 DR:74 LR:-326.8 LO:326.8);ALT=A[chr12:82144320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
