chr14	80106290	+	chr14	80115050	+	.	89	60	5815047_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=5815047_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_80115001_80140001_129C;SPAN=8760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:17 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:60 DR:89 LR:-399.4 LO:399.4);ALT=G[chr14:80115050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
