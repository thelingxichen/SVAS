chr10	127190418	-	chr10	127201102	+	.	23	64	6585311_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6585311_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_165C;SPAN=10684;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:76 DP:156 GQ:99 PL:[208.7, 0.0, 169.1] SR:64 DR:23 LR:-208.8 LO:208.8);ALT=[chr10:127201102[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	127190681	+	chr10	127197222	-	.	45	65	6585312_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCC;MAPQ=60;MATEID=6585312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_230C;SPAN=6541;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:92 DP:134 GQ:56.3 PL:[267.5, 0.0, 56.3] SR:65 DR:45 LR:-275.0 LO:275.0);ALT=C]chr10:127197222];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	127201222	+	chr10	127190797	+	.	35	48	6585315_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCACCAT;MAPQ=60;MATEID=6585315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_115C;SPAN=10425;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:75 DP:161 GQ:99 PL:[204.2, 0.0, 184.4] SR:48 DR:35 LR:-204.0 LO:204.0);ALT=]chr10:127201222]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	127191657	+	chr10	127197235	+	.	93	61	6585328_1	99.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=2;MATEID=6585328_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_143C;SPAN=5578;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:126 DP:129 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:61 DR:93 LR:-382.9 LO:382.9);ALT=C[chr10:127197235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127197257	+	chr10	127201101	+	.	10	0	6585350_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6585350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:127197257(+)-10:127201101(-)__10_127179501_127204501D;SPAN=3844;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:153 GQ:8.2 PL:[0.0, 8.2, 386.1] SR:0 DR:10 LR:8.442 LO:17.47);ALT=C[chr10:127201101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
