chr4	15642508	+	chr4	15656827	+	TAACATTCTTCAGTCCCTTTTCAAAGAGGCTAAGCATCTCGGAGAGTTTATTGTCAGAATGTACATTATAAATGGTCTGGCTGCGTTGTTGAAGCAAACCAATAATGTATTCATTTTCAATCTGCTCATGCATTTTGAACTCCTTGAAAGTAGCATACAAAGACTGCAGAAGAGCACGGAAATCGTTGTTGTTGGAAAAATTGGTTTTAGAAAG	0	10	1910516_1	28.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TAACATTCTTCAGTCCCTTTTCAAAGAGGCTAAGCATCTCGGAGAGTTTATTGTCAGAATGTACATTATAAATGGTCTGGCTGCGTTGTTGAAGCAAACCAATAATGTATTCATTTTCAATCTGCTCATGCATTTTGAACTCCTTGAAAGTAGCATACAAAGACTGCAGAAGAGCACGGAAATCGTTGTTGTTGGAAAAATTGGTTTTAGAAAG;MAPQ=60;MATEID=1910516_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_15631001_15656001_86C;SPAN=14319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:18 GQ:14.9 PL:[28.1, 0.0, 14.9] SR:10 DR:0 LR:-28.33 LO:28.33);ALT=T[chr4:15656827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15642508	+	chr4	15646116	+	.	2	5	1910515_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1910515_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_15631001_15656001_86C;SPAN=3608;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:46 GQ:10.7 PL:[10.7, 0.0, 99.8] SR:5 DR:2 LR:-10.64 LO:14.94);ALT=T[chr4:15646116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15646345	+	chr4	15656883	+	.	8	0	1910527_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1910527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:15646345(+)-4:15656883(-)__4_15631001_15656001D;SPAN=10538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:25 GQ:19.7 PL:[19.7, 0.0, 39.5] SR:0 DR:8 LR:-19.64 LO:20.05);ALT=T[chr4:15656883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15669709	+	chr4	15683031	+	.	8	0	1910455_1	19.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=1910455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:15669709(+)-4:15683031(-)__4_15680001_15705001D;SPAN=13322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:25 GQ:19.7 PL:[19.7, 0.0, 39.5] SR:0 DR:8 LR:-19.64 LO:20.05);ALT=T[chr4:15683031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15683526	+	chr4	15687857	+	.	30	5	1910469_1	91.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1910469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_15680001_15705001_222C;SPAN=4331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:77 GQ:91.4 PL:[91.4, 0.0, 94.7] SR:5 DR:30 LR:-91.37 LO:91.38);ALT=T[chr4:15687857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15704814	+	chr4	15707136	+	.	10	0	1910588_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1910588_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:15704814(+)-4:15707136(-)__4_15704501_15729501D;SPAN=2322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-14.05 LO:21.05);ALT=T[chr4:15707136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	15704956	+	chr4	15709132	+	AACAAGAACTGCACAGCCATCTGGGAAGCCTTTAAAGTGGCGCTGGACAAGGATCCCTGCTCCGTGCTGCCCTCAGACTATGACCTTTTTATTAACTTGTCCAGGCACTCTATTCCCAGAGATA	0	14	1910590_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AACAAGAACTGCACAGCCATCTGGGAAGCCTTTAAAGTGGCGCTGGACAAGGATCCCTGCTCCGTGCTGCCCTCAGACTATGACCTTTTTATTAACTTGTCCAGGCACTCTATTCCCAGAGATA;MAPQ=60;MATEID=1910590_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_15704501_15729501_76C;SPAN=4176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:60 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:14 DR:0 LR:-29.96 LO:32.8);ALT=G[chr4:15709132[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
