chr18	60697980	+	chr18	60779364	+	.	72	42	10040296_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GATAATT;MAPQ=60;MATEID=10040296_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_18_60686501_60711501_123C;SPAN=81384;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:9 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:42 DR:72 LR:-287.2 LO:287.2);ALT=T[chr18:60779364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	61330219	+	chr18	61312560	+	.	13	0	10041598_1	38.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=10041598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:61312560(-)-18:61330219(+)__18_61299001_61324001D;SPAN=17659;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:18 GQ:5 PL:[38.0, 0.0, 5.0] SR:0 DR:13 LR:-39.41 LO:39.41);ALT=]chr18:61330219]C;VARTYPE=BND:DUP-th;JOINTYPE=th
