chr7	158574893	+	chr7	158573702	+	.	9	0	3706917_1	11.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3706917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:158573702(-)-7:158574893(+)__7_158564001_158589001D;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=]chr7:158574893]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	158649441	+	chr7	158663832	+	AGAAGAACCAAAGATGATACCTGGAAAGCAGATGACCTCAGAAAACATCTCTG	8	14	3707009_1	54.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AGAAGAACCAAAGATGATACCTGGAAAGCAGATGACCTCAGAAAACATCTCTG;MAPQ=60;MATEID=3707009_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_158662001_158687001_279C;SPAN=14391;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:31 GQ:18.2 PL:[54.5, 0.0, 18.2] SR:14 DR:8 LR:-55.13 LO:55.13);ALT=G[chr7:158663832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	158649441	+	chr7	158662544	+	.	4	5	3707008_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3707008_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_7_158662001_158687001_279C;SPAN=13103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:16 PL:[16.0, 0.0, 16.0] SR:5 DR:4 LR:-15.94 LO:15.94);ALT=G[chr7:158662544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	158853486	+	chr7	158852427	+	.	17	0	3707214_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3707214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:158852427(-)-7:158853486(+)__7_158833501_158858501D;SPAN=1059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:79 GQ:34.7 PL:[34.7, 0.0, 156.8] SR:0 DR:17 LR:-34.71 LO:39.14);ALT=]chr7:158853486]A;VARTYPE=BND:DUP-th;JOINTYPE=th
