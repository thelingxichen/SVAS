chrX	140476730	+	chrX	140479227	+	.	0	27	7541155_1	79.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=7541155_2;MATENM=7;NM=0;NUMPARTS=2;SCTG=c_23_140458501_140483501_103C;SPAN=2497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:14 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:27 DR:0 LR:-79.22 LO:79.22);ALT=A[chrX:140479227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
