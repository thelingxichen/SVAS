chr18	66377381	+	chr18	66381081	+	ATCTACAAGCCAAATGTCATCATTTCGATTTTCTTTAA	0	7	6661981_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=ATCTACAAGCCAAATGTCATCATTTCGATTTTCTTTAA;MAPQ=60;MATEID=6661981_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_66370501_66395501_138C;SPAN=3700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:54 GQ:8.6 PL:[8.6, 0.0, 120.8] SR:7 DR:0 LR:-8.477 LO:14.41);ALT=A[chr18:66381081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	66379462	+	chr18	66382826	+	.	32	14	6661984_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6661984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_66370501_66395501_98C;SPAN=3364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:57 GQ:20.9 PL:[116.6, 0.0, 20.9] SR:14 DR:32 LR:-120.3 LO:120.3);ALT=G[chr18:66382826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
