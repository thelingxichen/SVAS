chr8	144139901	-	chr8	144141752	+	.	10	0	5751035_1	3.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5751035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144139901(-)-8:144141752(-)__8_144133501_144158501D;SPAN=1851;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:108 GQ:3.8 PL:[3.8, 0.0, 257.9] SR:0 DR:10 LR:-3.75 LO:19.04);ALT=[chr8:144141752[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	144704918	+	chr8	144561423	+	GCTGA	94	25	5753211_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GCTGA;MAPQ=60;MATEID=5753211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144697001_144722001_54C;SPAN=143495;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:43 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:25 DR:94 LR:-326.8 LO:326.8);ALT=]chr8:144704918]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	144634067	+	chr8	144636240	+	.	0	156	5753635_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TGT;MAPQ=60;MATEID=5753635_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_144623501_144648501_79C;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:156 DP:111 GQ:42.1 PL:[462.1, 42.1, 0.0] SR:156 DR:0 LR:-462.1 LO:462.1);ALT=T[chr8:144636240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144700487	+	chr8	144714693	+	.	56	34	5753225_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=5753225_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144697001_144722001_115C;SPAN=14206;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:73 DP:95 GQ:14 PL:[215.3, 0.0, 14.0] SR:34 DR:56 LR:-225.5 LO:225.5);ALT=A[chr8:144714693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144716355	+	chr15	98558153	+	.	20	0	9097648_1	50.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=9097648_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144716355(+)-15:98558153(-)__15_98539001_98564001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:59 GQ:50 PL:[50.0, 0.0, 92.9] SR:0 DR:20 LR:-50.04 LO:50.75);ALT=T[chr15:98558153[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	145104681	+	chr8	144965983	+	.	74	26	5755412_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=5755412_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_145089001_145114001_60C;SPAN=138698;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:68 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:26 DR:74 LR:-267.4 LO:267.4);ALT=]chr8:145104681]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	145788015	+	chr8	145786646	+	.	6	10	5757963_1	4.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=ACCCCAGTGGTTTCCATC;MAPQ=10;MATEID=5757963_2;MATENM=1;NM=0;NUMPARTS=2;REPSEQ=CCCC;SCTG=c_8_145775001_145800001_153C;SECONDARY;SPAN=1369;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:180 GQ:4 PL:[4.0, 0.0, 433.1] SR:10 DR:6 LR:-4.05 LO:30.16);ALT=]chr8:145788015]A;VARTYPE=BND:DUP-th;JOINTYPE=th
