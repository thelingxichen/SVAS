chrX	97163465	+	chrX	97164469	+	.	13	0	7479812_1	33.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=7479812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:97163465(+)-23:97164469(-)__23_97142501_97167501D;SPAN=1004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:0 DR:13 LR:-33.7 LO:33.85);ALT=G[chrX:97164469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
