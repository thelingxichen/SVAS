chr3	186327788	+	chr3	119049964	+	.	0	37	4082317_1	99.0	.	BX=GCCACTTAGGCATTTC-1_1,CCAATCCAGTATCTCG-1_1,GTGGCACTCCCAACGG-1_1,AGGCGAAGTCGTTGGC-1_2,TACTTGTTCGTGGTCG-1_1,TGCCCTAGTGAAATCA-1_1,GGCAATTTCGTATCAG-1_2,CTGGTCTAGCTCGCTG-1_1,CTGTAAGTCTTCACGC-1_1,ATGCGGCCAAACCGAG-1_2,ATCTATCGTAACGACG-1_2,GTTGCCTGTAAGAGAG-1_1,GACACATTCAACGATC-1_1,CTATCTAGTCTTACCC-1_2,GGGCCATGTCAACCGC-1_2,CTCACACGTACGAAAT-1_1,ACACCGGAGTGGACAC-1_1,GAGATGGAGCAGTCTT-1_1,CCACCTAAGTGAGAAG-1_1,GTTTGAGTCACGACGC-1_2,AGTAGTCAGACAGATT-1_1,ATGCGGCGTCTCAACA-1_1,CGGTGACTCGAGAAGC-1_1,CTACCCACACTTGGAT-1_1,CGCAAGCAGCACAGGT-1_1,GCTCTGTGTTGCGGCT-1_1,TCGAAACCAACGCACC-1_1;EVDNC=ASSMB;HOMSEQ=TGA;MAPQ=60;MATEID=4082317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_186322501_186347501_50C;SPAN=67277824;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:19 GQ:5.1 PL:[0.0, 5.1, 56.1] SR:0 DR:0 LR:5.338 LO:0.0),OC001T.bam(GT:0/1 AD:37 DP:54 GQ:27.8 PL:[107.0, 0.0, 27.8] SR:37 DR:0 LR:-109.5 LO:109.5);ALT=]chr3:186327788]T;VARTYPE=BND:DUP-th;JOINTYPE=th	.
chr3	186327788	+	chr3	119049964	+	.	0	37	4082317_1	99.0	.	BX=GCCACTTAGGCATTTC-1_1,CCAATCCAGTATCTCG-1_1,GTGGCACTCCCAACGG-1_1,AGGCGAAGTCGTTGGC-1_2,TACTTGTTCGTGGTCG-1_1,TGCCCTAGTGAAATCA-1_1,GGCAATTTCGTATCAG-1_2,CTGGTCTAGCTCGCTG-1_1,CTGTAAGTCTTCACGC-1_1,ATGCGGCCAAACCGAG-1_2,ATCTATCGTAACGACG-1_2,GTTGCCTGTAAGAGAG-1_1,GACACATTCAACGATC-1_1,CTATCTAGTCTTACCC-1_2,GGGCCATGTCAACCGC-1_2,CTCACACGTACGAAAT-1_1,ACACCGGAGTGGACAC-1_1,GAGATGGAGCAGTCTT-1_1,CCACCTAAGTGAGAAG-1_1,GTTTGAGTCACGACGC-1_2,AGTAGTCAGACAGATT-1_1,ATGCGGCGTCTCAACA-1_1,CGGTGACTCGAGAAGC-1_1,CTACCCACACTTGGAT-1_1,CGCAAGCAGCACAGGT-1_1,GCTCTGTGTTGCGGCT-1_1,TCGAAACCAACGCACC-1_1;EVDNC=ASSMB;HOMSEQ=TGA;MAPQ=60;MATEID=4082317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_186322501_186347501_50C;SPAN=67277824;SVTYPE=BND;TOOL=svaba;GENOTYPE=OC001B.bam(GT:0/0 AD:0 DP:19 GQ:5.1 PL:[0.0, 5.1, 56.1] SR:0 DR:0 LR:5.338 LO:0.0),OC001T.bam(GT:0/1 AD:37 DP:54 GQ:27.8 PL:[107.0, 0.0, 27.8] SR:37 DR:0 LR:-109.5 LO:109.5);ALT=]chr3:186327788]T;VARTYPE=BND:DUP-th;JOINTYPE=th	.
