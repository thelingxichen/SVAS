chr8	110106059	-	chr8	110107260	+	.	4	2	5614623_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAGCAAAAGTT;MAPQ=60;MATEID=5614623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110103001_110128001_76C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:141 GQ:18 PL:[0.0, 18.0, 376.2] SR:2 DR:4 LR:18.39 LO:9.336);ALT=[chr8:110107260[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
