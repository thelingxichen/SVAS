chr12	39242466	+	chr12	39299239	+	CTCTCCATTCTTTATTTCCAACTCCTTGTACATATAAGACACAAATTGGATCAGATTTAGAAAATGTGTCTCTGTCAAGAAGATTT	0	24	5156827_1	67.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTCTCCATTCTTTATTTCCAACTCCTTGTACATATAAGACACAAATTGGATCAGATTTAGAAAATGTGTCTCTGTCAAGAAGATTT;MAPQ=60;MATEID=5156827_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_39298001_39323001_346C;SPAN=56773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:43 GQ:34.7 PL:[67.7, 0.0, 34.7] SR:24 DR:0 LR:-68.06 LO:68.06);ALT=T[chr12:39299239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
