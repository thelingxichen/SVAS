chr12	69172523	+	chr12	69174356	-	.	8	0	7701627_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=7701627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69172523(+)-12:69174356(+)__12_69163501_69188501D;SPAN=1833;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:322 GQ:60.5 PL:[0.0, 60.5, 901.1] SR:0 DR:8 LR:60.83 LO:10.57);ALT=T]chr12:69174356];VARTYPE=BND:INV-hh;JOINTYPE=hh
