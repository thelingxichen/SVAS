chr20	1389146	+	chr20	1390815	+	.	96	66	10398953_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=10398953_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_20_1372001_1397001_239C;SPAN=1669;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:133 DP:22 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:66 DR:96 LR:-392.8 LO:392.8);ALT=A[chr20:1390815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
