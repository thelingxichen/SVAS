chrX	88462513	+	chrX	88460958	+	GTTTT	65	24	7469846_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;INSERTION=GTTTT;MAPQ=60;MATEID=7469846_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_23_88445001_88470001_229C;SPAN=1555;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:145 GQ:99 PL:[228.2, 0.0, 122.6] SR:24 DR:65 LR:-229.8 LO:229.8);ALT=]chrX:88462513]T;VARTYPE=BND:DUP-th;JOINTYPE=th
