chr8	47405851	+	chr8	47407911	+	.	35	25	3843975_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGAGCT;MAPQ=60;MATEID=3843975_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_47383001_47408001_185C;SPAN=2060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:60 GQ:3 PL:[151.8, 3.0, 0.0] SR:25 DR:35 LR:-158.8 LO:158.8);ALT=T[chr8:47407911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	47768069	+	chr8	47769814	+	.	58	28	3844931_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCCTGGTTTCTGCCCACAT;MAPQ=60;MATEID=3844931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_47750501_47775501_237C;SPAN=1745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:67 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:28 DR:58 LR:-224.5 LO:224.5);ALT=T[chr8:47769814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	48711953	+	chr8	48713352	+	.	3	2	3847524_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=3847524_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_48706001_48731001_315C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:87 GQ:10.2 PL:[0.0, 10.2, 231.0] SR:2 DR:3 LR:10.37 LO:6.36);ALT=T[chr8:48713352[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	48868510	+	chr8	48869731	+	.	0	9	3847948_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3847948_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_48853001_48878001_86C;SPAN=1221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-8.035 LO:17.94);ALT=T[chr8:48869731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	48869992	+	chr8	48872533	+	.	0	10	3847956_1	8.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=3847956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_48853001_48878001_237C;SPAN=2541;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:10 DR:0 LR:-8.085 LO:19.77);ALT=C[chr8:48872533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	48921078	+	chr8	48955607	+	.	8	0	3848348_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3848348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:48921078(+)-8:48955607(-)__8_48951001_48976001D;SPAN=34529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.57 LO:18.13);ALT=T[chr8:48955607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
