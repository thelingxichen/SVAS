chr16	55814267	-	chr16	55850425	+	.	12	0	9332058_1	23.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=9332058_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:55814267(-)-16:55850425(-)__16_55811001_55836001D;SPAN=36158;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:61 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:0 DR:12 LR:-23.09 LO:27.1);ALT=[chr16:55850425[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	57002919	+	chr16	56846831	+	A	80	29	9336889_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=9336889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_56987001_57012001_293C;SPAN=156088;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:77 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:29 DR:80 LR:-283.9 LO:283.9);ALT=]chr16:57002919]C;VARTYPE=BND:DUP-th;JOINTYPE=th
