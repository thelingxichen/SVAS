chr21	16588380	+	chr21	16591453	+	.	80	47	10712126_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=10712126_2;MATENM=2;NM=3;NUMPARTS=2;SCTG=c_21_16586501_16611501_167C;SPAN=3073;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:23 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:47 DR:80 LR:-310.3 LO:310.3);ALT=T[chr21:16591453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
