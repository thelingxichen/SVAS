chr16	76539133	+	chr16	76544026	+	C	152	128	9427720_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=9427720_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_76538001_76563001_141C;SPAN=4893;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:217 DP:47 GQ:58.6 PL:[643.6, 58.6, 0.0] SR:128 DR:152 LR:-643.7 LO:643.7);ALT=G[chr16:76544026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
