chrX	66198859	-	chrX	66200135	+	.	11	0	11211158_1	20.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=11211158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:66198859(-)-23:66200135(-)__23_66174501_66199501D;SPAN=1276;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:60 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-20.06 LO:24.46);ALT=[chrX:66200135[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	66483150	+	chrX	66484329	+	.	0	47	11212109_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GTTT;MAPQ=60;MATEID=11212109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_66468501_66493501_28C;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:47 DP:87 GQ:78.8 PL:[131.6, 0.0, 78.8] SR:47 DR:0 LR:-132.3 LO:132.3);ALT=T[chrX:66484329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
