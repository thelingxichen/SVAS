chr3	120911834	+	chr3	121577522	-	.	24	0	2281508_1	60.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2281508_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:120911834(+)-3:121577522(+)__3_121569001_121594001D;SPAN=665688;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:24 DP:69 GQ:60.5 PL:[60.5, 0.0, 106.7] SR:0 DR:24 LR:-60.53 LO:61.24);ALT=T]chr3:121577522];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	120912265	-	chr3	121577015	+	.	39	0	2281509_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=2281509_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:120912265(-)-3:121577015(-)__3_121569001_121594001D;SPAN=664750;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:87 GQ:99 PL:[105.2, 0.0, 105.2] SR:0 DR:39 LR:-105.2 LO:105.2);ALT=[chr3:121577015[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
