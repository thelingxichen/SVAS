chr4	73552249	+	chr4	73561109	+	CCATGA	38	40	2029082_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAACATG;INSERTION=CCATGA;MAPQ=60;MATEID=2029082_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_73549001_73574001_257C;SPAN=8860;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:78 GQ:7.8 PL:[204.6, 7.8, 0.0] SR:40 DR:38 LR:-210.9 LO:210.9);ALT=A[chr4:73561109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
