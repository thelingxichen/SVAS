chr3	3215994	+	chr3	3221304	+	.	31	0	1271241_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1271241_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:3215994(+)-3:3221304(-)__3_3209501_3234501D;SPAN=5310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:47 GQ:23.6 PL:[89.6, 0.0, 23.6] SR:0 DR:31 LR:-91.67 LO:91.67);ALT=A[chr3:3221304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	3216954	+	chr3	3221305	+	.	11	4	1271242_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1271242_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_3209501_3234501_121C;SPAN=4351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:54 GQ:25.1 PL:[25.1, 0.0, 104.3] SR:4 DR:11 LR:-24.98 LO:27.82);ALT=C[chr3:3221305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	4066937	+	chr3	4069556	+	.	44	35	1272384_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACAAAATATATAT;MAPQ=60;MATEID=1272384_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_4067001_4092001_94C;SPAN=2619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:11 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:35 DR:44 LR:-178.2 LO:178.2);ALT=T[chr3:4069556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	4899428	-	chr3	4900643	+	.	10	0	1273697_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1273697_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:4899428(-)-3:4900643(-)__3_4900001_4925001D;SPAN=1215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:38 GQ:22.7 PL:[22.7, 0.0, 68.9] SR:0 DR:10 LR:-22.72 LO:24.04);ALT=[chr3:4900643[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
