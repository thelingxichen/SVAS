chr20	50759206	+	chr20	50760929	+	.	96	73	10612051_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CAACATGGTGAAACCC;MAPQ=8;MATEID=10612051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_50739501_50764501_333C;SPAN=1723;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:141 DP:124 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:73 DR:96 LR:-415.9 LO:415.9);ALT=C[chr20:50760929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
