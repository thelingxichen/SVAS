chr4	188495200	-	chr4	188496243	+	.	8	0	3128959_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3128959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:188495200(-)-4:188496243(-)__4_188478501_188503501D;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.374 LO:14.01);ALT=[chr4:188496243[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	188812926	+	chr4	189257567	-	.	10	0	3131168_1	24.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3131168_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:188812926(+)-4:189257567(+)__4_189238001_189263001D;SPAN=444641;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:31 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:0 DR:10 LR:-24.61 LO:25.11);ALT=C]chr4:189257567];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	188813069	-	chr4	189257420	+	.	18	0	3131169_1	50.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3131169_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:188813069(-)-4:189257420(-)__4_189238001_189263001D;SPAN=444351;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:35 GQ:33.5 PL:[50.0, 0.0, 33.5] SR:0 DR:18 LR:-50.08 LO:50.08);ALT=[chr4:189257420[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	189071570	+	chr4	189433213	+	GGG	60	30	3131511_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;INSERTION=GGG;MAPQ=60;MATEID=3131511_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_189409501_189434501_143C;SPAN=361643;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:53 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:30 DR:60 LR:-247.6 LO:247.6);ALT=A[chr4:189433213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	189437078	+	chr4	189438907	+	.	54	37	3131602_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=3131602_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_189434001_189459001_105C;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:72 DP:78 GQ:21 PL:[231.0, 21.0, 0.0] SR:37 DR:54 LR:-231.1 LO:231.1);ALT=G[chr4:189438907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	189463410	+	chr4	189467440	+	.	67	54	3131792_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3131792_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_4_189458501_189483501_5C;SPAN=4030;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:65 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:54 DR:67 LR:-280.6 LO:280.6);ALT=T[chr4:189467440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	190058014	+	chr4	190064273	+	.	58	52	3134096_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGACTGGGTAATTTAT;MAPQ=60;MATEID=3134096_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_190046501_190071501_407C;SPAN=6259;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:78 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:52 DR:58 LR:-303.7 LO:303.7);ALT=T[chr4:190064273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
