chr9	71895379	+	chr9	71896579	+	.	29	0	5884040_1	92.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5884040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:71895379(+)-9:71896579(-)__9_71883001_71908001D;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:32 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:29 LR:-92.42 LO:92.42);ALT=C[chr9:71896579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
