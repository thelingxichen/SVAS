chr13	111563120	+	chr13	111567072	+	.	0	7	5647948_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CTT;MAPQ=60;MATEID=5647948_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_111548501_111573501_59C;SPAN=3952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:68 GQ:4.7 PL:[4.7, 0.0, 159.8] SR:7 DR:0 LR:-4.684 LO:13.67);ALT=T[chr13:111567072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
