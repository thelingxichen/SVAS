chr10	122226705	+	chr10	122228783	+	.	134	0	6563219_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=6563219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:122226705(+)-10:122228783(-)__10_122206001_122231001D;SPAN=2078;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:134 DP:23 GQ:36 PL:[396.0, 36.0, 0.0] SR:0 DR:134 LR:-396.1 LO:396.1);ALT=C[chr10:122228783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
