chr6	161275015	+	chr6	161273854	+	.	25	0	3100728_1	68.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=3100728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:161273854(-)-6:161275015(+)__6_161259001_161284001D;SPAN=1161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:50 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:0 DR:25 LR:-69.1 LO:69.1);ALT=]chr6:161275015]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	161851868	+	chr6	161486970	+	.	15	25	3103229_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAAAAAAAA;MAPQ=60;MATEID=3103229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_161847001_161872001_30C;SPAN=364898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:34 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:25 DR:15 LR:-112.2 LO:112.2);ALT=]chr6:161851868]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	161653336	+	chr6	161694970	+	.	4	2	3102650_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3102650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_161651001_161676001_56C;SPAN=41634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:36 GQ:6.8 PL:[6.8, 0.0, 79.4] SR:2 DR:4 LR:-6.752 LO:10.46);ALT=T[chr6:161694970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	161726309	+	chr6	161727860	+	.	49	48	3102736_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGCACTTTGGGAGGC;MAPQ=60;MATEID=3102736_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_161724501_161749501_69C;SPAN=1551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:69 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:48 DR:49 LR:-227.8 LO:227.8);ALT=C[chr6:161727860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	161833926	+	chr6	161832731	+	.	17	0	3102982_1	32.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=3102982_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:161832731(-)-6:161833926(+)__6_161822501_161847501D;SPAN=1195;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:89 GQ:32 PL:[32.0, 0.0, 183.8] SR:0 DR:17 LR:-32.01 LO:38.15);ALT=]chr6:161833926]T;VARTYPE=BND:DUP-th;JOINTYPE=th
