chr21	35139286	+	chr21	35140725	-	.	8	0	10763854_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=10763854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:35139286(+)-21:35140725(+)__21_35133001_35158001D;SPAN=1439;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:151 GQ:14.2 PL:[0.0, 14.2, 392.7] SR:0 DR:8 LR:14.5 LO:13.22);ALT=A]chr21:35140725];VARTYPE=BND:INV-hh;JOINTYPE=hh
