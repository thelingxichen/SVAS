chr1	83125976	+	chr1	83127570	+	.	56	41	383319_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAAATGGTTCATGC;MAPQ=60;MATEID=383319_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_83104001_83129001_323C;SPAN=1594;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:82 DP:76 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:41 DR:56 LR:-241.0 LO:241.0);ALT=C[chr1:83127570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	83479305	+	chr1	208739015	-	.	12	31	785229_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=GAATAGAATAGAATAGAATAGAATAGAATAGAATAGAATAG;MAPQ=60;MATEID=785229_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_208715501_208740501_160C;SPAN=125259710;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:52 GQ:9.2 PL:[114.8, 0.0, 9.2] SR:31 DR:12 LR:-119.6 LO:119.6);ALT=G]chr1:208739015];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	209627215	+	chr1	213087955	+	.	13	0	804816_1	21.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=804816_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:209627215(+)-1:213087955(-)__1_213076501_213101501D;SPAN=3460740;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:78 GQ:21.8 PL:[21.8, 0.0, 167.0] SR:0 DR:13 LR:-21.78 LO:28.31);ALT=T[chr1:213087955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	209936059	+	chr1	209935008	+	GCTGCCCCAGCTCACTTAGTAA	0	42	790169_1	99.0	.	EVDNC=ASSMB;INSERTION=GCTGCCCCAGCTCACTTAGTAA;MAPQ=60;MATEID=790169_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_1_209916001_209941001_162C;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:42 DP:131 GQ:99 PL:[103.4, 0.0, 212.3] SR:42 DR:0 LR:-103.2 LO:105.3);ALT=]chr1:209936059]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	212264750	+	chr1	212266287	-	.	8	0	800134_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=800134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:212264750(+)-1:212266287(+)__1_212243501_212268501D;SPAN=1537;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:134 GQ:9.6 PL:[0.0, 9.6, 343.2] SR:0 DR:8 LR:9.896 LO:13.65);ALT=G]chr1:212266287];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	212471153	+	chr1	212472617	+	.	45	30	801362_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGATGAAGTGAATTGTT;MAPQ=60;MATEID=801362_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212464001_212489001_163C;SPAN=1464;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:64 DP:62 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:30 DR:45 LR:-188.1 LO:188.1);ALT=T[chr1:212472617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	213380313	+	chr1	213381320	-	.	9	0	806076_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=806076_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:213380313(+)-1:213381320(+)__1_213370501_213395501D;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:134 GQ:6.3 PL:[0.0, 6.3, 336.6] SR:0 DR:9 LR:6.595 LO:15.83);ALT=G]chr1:213381320];VARTYPE=BND:INV-hh;JOINTYPE=hh
