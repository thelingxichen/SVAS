chr3	111261157	+	chr3	111263892	+	.	51	19	1589570_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1589570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_111254501_111279501_306C;SPAN=2735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:126 GQ:99 PL:[147.5, 0.0, 157.4] SR:19 DR:51 LR:-147.4 LO:147.4);ALT=G[chr3:111263892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	111286495	+	chr3	111297873	+	.	3	3	1589125_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1589125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_111279001_111304001_173C;SPAN=11378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:100 GQ:10.5 PL:[0.0, 10.5, 264.0] SR:3 DR:3 LR:10.59 LO:8.136);ALT=G[chr3:111297873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	111698050	+	chr3	111700629	+	.	8	9	1590855_1	8.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1590855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_111695501_111720501_348C;SPAN=2579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:105 GQ:8 PL:[8.0, 0.0, 245.6] SR:9 DR:8 LR:-7.864 LO:21.56);ALT=G[chr3:111700629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112052113	+	chr3	112063806	+	.	26	0	1591749_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1591749_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:112052113(+)-3:112063806(-)__3_112063001_112088001D;SPAN=11693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:61 GQ:69.5 PL:[69.5, 0.0, 76.1] SR:0 DR:26 LR:-69.3 LO:69.33);ALT=C[chr3:112063806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112253186	+	chr3	112255321	+	.	3	8	1592408_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1592408_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_112234501_112259501_211C;SPAN=2135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:8 DR:3 LR:-5.918 LO:19.39);ALT=T[chr3:112255321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112256739	+	chr3	112262903	+	CATCTGTTTCCAACAATCCACTCTCTTCATATTCTTCCATATCTGCAGCTTCTCCTTCATCTTCATCTTCTTCCTCTTCACATAGTGCTGAGCAATCTTGAAGCCTTATATTGT	3	18	1592683_1	49.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTT;INSERTION=CATCTGTTTCCAACAATCCACTCTCTTCATATTCTTCCATATCTGCAGCTTCTCCTTCATCTTCATCTTCTTCCTCTTCACATAGTGCTGAGCAATCTTGAAGCCTTATATTGT;MAPQ=60;MATEID=1592683_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_112259001_112284001_416C;SPAN=6164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:49 GQ:49.4 PL:[49.4, 0.0, 69.2] SR:18 DR:3 LR:-49.44 LO:49.63);ALT=T[chr3:112262903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112260761	+	chr3	112267376	+	.	8	0	1592691_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1592691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:112260761(+)-3:112267376(-)__3_112259001_112284001D;SPAN=6615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=T[chr3:112267376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112267488	+	chr3	112269039	+	.	0	14	1592710_1	17.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1592710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_112259001_112284001_148C;SPAN=1551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:108 GQ:17 PL:[17.0, 0.0, 244.7] SR:14 DR:0 LR:-16.95 LO:28.83);ALT=C[chr3:112269039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112269110	+	chr3	112280303	+	ATTGCCATGTTGGACAGTGGTGGACTAGGTGATCTCCAGCTGCCACAAACTCTTCTGGGGTAATTACACCTGTTTCCTTAAACTTTGATT	6	50	1592720_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=ATTGCCATGTTGGACAGTGGTGGACTAGGTGATCTCCAGCTGCCACAAACTCTTCTGGGGTAATTACACCTGTTTCCTTAAACTTTGATT;MAPQ=60;MATEID=1592720_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_112259001_112284001_5C;SPAN=11193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:120 GQ:99 PL:[132.5, 0.0, 158.9] SR:50 DR:6 LR:-132.5 LO:132.7);ALT=C[chr3:112280303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112272230	+	chr3	112280423	+	.	8	0	1592729_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1592729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:112272230(+)-3:112280423(-)__3_112259001_112284001D;SPAN=8193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:0 DR:8 LR:5.29 LO:14.13);ALT=C[chr3:112280423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112281124	+	chr3	112282230	+	.	4	4	1592763_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTAA;MAPQ=60;MATEID=1592763_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_112259001_112284001_402C;SPAN=1106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:115 GQ:7.8 PL:[0.0, 7.8, 293.7] SR:4 DR:4 LR:8.049 LO:12.0);ALT=A[chr3:112282230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	112736476	+	chr3	112738450	+	.	8	0	1593900_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1593900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:112736476(+)-3:112738450(-)__3_112724501_112749501D;SPAN=1974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:119 GQ:5.7 PL:[0.0, 5.7, 300.3] SR:0 DR:8 LR:5.832 LO:14.07);ALT=T[chr3:112738450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	113345064	+	chr3	113346492	+	.	0	4	1595946_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=1595946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_113337001_113362001_300C;SPAN=1428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:108 GQ:15.9 PL:[0.0, 15.9, 293.7] SR:4 DR:0 LR:16.06 LO:5.98);ALT=T[chr3:113346492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	113442943	+	chr3	113464789	+	.	5	4	1596399_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1596399_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_113459501_113484501_169C;SPAN=21846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:61 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:4 DR:5 LR:-13.18 LO:19.08);ALT=C[chr3:113464789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	113466001	+	chr3	113499895	+	.	10	0	1596621_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1596621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:113466001(+)-3:113499895(-)__3_113484001_113509001D;SPAN=33894;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:0 DR:10 LR:-15.67 LO:21.47);ALT=G[chr3:113499895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
