chr2	45292658	+	chr2	45302937	-	.	16	0	982763_1	43.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=982763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:45292658(+)-2:45302937(+)__2_45276001_45301001D;SPAN=10279;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:35 GQ:40.1 PL:[43.4, 0.0, 40.1] SR:0 DR:16 LR:-43.34 LO:43.34);ALT=T]chr2:45302937];VARTYPE=BND:INV-hh;JOINTYPE=hh
