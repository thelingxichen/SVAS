chr6	103737464	+	chr6	103762890	+	GCCA	0	19	2965285_1	55.0	.	EVDNC=ASSMB;INSERTION=GCCA;MAPQ=60;MATEID=2965285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_103757501_103782501_9C;SPAN=25426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:27 GQ:9.2 PL:[55.4, 0.0, 9.2] SR:19 DR:0 LR:-57.18 LO:57.18);ALT=T[chr6:103762890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
