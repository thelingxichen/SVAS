chr7	83251681	+	chr7	83253881	-	.	8	0	5010138_1	23.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5010138_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:83251681(+)-7:83253881(+)__7_83226501_83251501D;SPAN=2200;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:8 DP:0 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=C]chr7:83253881];VARTYPE=BND:INV-hh;JOINTYPE=hh
