chr3	26767297	+	chr3	26759838	+	.	54	56	1905481_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1905481_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_26754001_26779001_136C;SPAN=7459;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:87 DP:123 GQ:42.8 PL:[254.0, 0.0, 42.8] SR:56 DR:54 LR:-262.2 LO:262.2);ALT=]chr3:26767297]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	27111741	+	chr20	53286216	+	.	6	18	1906506_1	56.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=AATAATAATAATAATAATAAT;MAPQ=44;MATEID=1906506_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_27097001_27122001_260C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:35 GQ:26.9 PL:[56.6, 0.0, 26.9] SR:18 DR:6 LR:-57.04 LO:57.04);ALT=T[chr20:53286216[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
