chr17	13972967	+	chr17	13977638	+	.	8	3	6321985_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=6321985_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_13965001_13990001_156C;SPAN=4671;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:3 DR:8 LR:-11.02 LO:18.56);ALT=T[chr17:13977638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	14189911	+	chr17	14191556	+	.	58	38	6322347_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=6322347_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_17_14185501_14210501_94C;SPAN=1645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:40 GQ:21 PL:[231.0, 21.0, 0.0] SR:38 DR:58 LR:-231.1 LO:231.1);ALT=A[chr17:14191556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	14659428	+	chr17	14662387	-	.	13	0	6323867_1	26.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=6323867_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:14659428(+)-17:14662387(+)__17_14651001_14676001D;SPAN=2959;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:63 GQ:26 PL:[26.0, 0.0, 125.0] SR:0 DR:13 LR:-25.84 LO:29.66);ALT=G]chr17:14662387];VARTYPE=BND:INV-hh;JOINTYPE=hh
