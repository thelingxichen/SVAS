chr20	35679167	+	chr20	35683050	+	.	10	0	10513182_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=10513182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35679167(+)-20:35683050(-)__20_35672001_35697001D;SPAN=3883;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:238 GQ:31.3 PL:[0.0, 31.3, 640.3] SR:0 DR:10 LR:31.47 LO:15.5);ALT=G[chr20:35683050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
