chr9	84324363	+	chr9	84326927	+	.	73	28	5907089_1	49.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TAAAATGGCTCTAGC;MAPQ=60;MATEID=5907089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_84304501_84329501_229C;SPAN=2564;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:87 DP:878 GQ:49.5 PL:[49.5, 0.0, 2083.0] SR:28 DR:73 LR:-49.32 LO:168.3);ALT=C[chr9:84326927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	84930646	+	chr9	84932455	+	.	60	49	5908097_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5908097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_84917001_84942001_206C;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:17 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:49 DR:60 LR:-260.8 LO:260.8);ALT=T[chr9:84932455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
