chr6	132793514	+	chr6	132824585	+	AACTGTTGCCTCAATTCAGGTGAATCTTGAGGTGTTCCAAGTTGATTCAGAGTTCTTTGTATTTCCACAG	0	21	3031668_1	58.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AACTGTTGCCTCAATTCAGGTGAATCTTGAGGTGTTCCAAGTTGATTCAGAGTTCTTTGTATTTCCACAG;MAPQ=60;MATEID=3031668_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_132814501_132839501_41C;SPAN=31071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:42 GQ:41.6 PL:[58.1, 0.0, 41.6] SR:21 DR:0 LR:-58.04 LO:58.04);ALT=C[chr6:132824585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	132796844	+	chr6	132834143	+	.	12	0	3031671_1	26.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3031671_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:132796844(+)-6:132834143(-)__6_132814501_132839501D;SPAN=37299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:49 GQ:26.3 PL:[26.3, 0.0, 92.3] SR:0 DR:12 LR:-26.34 LO:28.41);ALT=A[chr6:132834143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	132824729	+	chr6	132834144	+	.	16	6	3031697_1	41.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=3031697_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_132814501_132839501_6C;SPAN=9415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:89 GQ:41.9 PL:[41.9, 0.0, 173.9] SR:6 DR:16 LR:-41.91 LO:46.48);ALT=T[chr6:132834144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	133341834	+	chr6	133347886	+	.	66	22	3033172_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTGTGATGTTTT;MAPQ=60;MATEID=3033172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_133329001_133354001_39C;SPAN=6052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:289 GQ:99 PL:[251.8, 0.0, 449.9] SR:22 DR:66 LR:-251.8 LO:254.9);ALT=T[chr6:133347886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
