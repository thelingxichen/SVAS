chr10	32257895	+	chr10	32260613	+	.	53	47	6180422_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAGATATTAGTTG;MAPQ=60;MATEID=6180422_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_32242001_32267001_174C;SPAN=2718;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:96 GQ:15.9 PL:[264.0, 15.9, 0.0] SR:47 DR:53 LR:-267.7 LO:267.7);ALT=G[chr10:32260613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
