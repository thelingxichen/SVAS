chr15	41571293	-	chr15	41572739	+	.	9	0	8871143_1	2.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=8871143_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:41571293(-)-15:41572739(-)__15_41552001_41577001D;SPAN=1446;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=[chr15:41572739[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
