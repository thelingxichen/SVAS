chr3	106894706	-	chr3	106897160	+	.	8	0	1575047_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1575047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:106894706(-)-3:106897160(-)__3_106893501_106918501D;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:0 DR:8 LR:0.6845 LO:14.7);ALT=[chr3:106897160[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	107037949	+	chr3	107040333	+	AAAAT	0	52	1575449_1	99.0	.	EVDNC=ASSMB;INSERTION=AAAAT;MAPQ=60;MATEID=1575449_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107016001_107041001_373C;SPAN=2384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:83 GQ:50.3 PL:[149.3, 0.0, 50.3] SR:52 DR:0 LR:-151.7 LO:151.7);ALT=G[chr3:107040333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107766140	+	chr3	107776324	+	CTAGGAGGTTGTATAGTCTTCTGATTGGAAG	2	22	1578060_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTAGGAGGTTGTATAGTCTTCTGATTGGAAG;MAPQ=60;MATEID=1578060_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107775501_107800501_170C;SPAN=10184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:47 GQ:50 PL:[63.2, 0.0, 50.0] SR:22 DR:2 LR:-63.26 LO:63.26);ALT=C[chr3:107776324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107799192	+	chr3	107809709	+	.	95	52	1578139_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1578139_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107775501_107800501_182C;SPAN=10517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:114 DP:56 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:52 DR:95 LR:-336.7 LO:336.7);ALT=C[chr3:107809709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107881503	+	chr3	107882510	+	.	0	7	1577903_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1577903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107873501_107898501_172C;SPAN=1007;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:114 GQ:7.5 PL:[0.0, 7.5, 290.4] SR:7 DR:0 LR:7.778 LO:12.03);ALT=C[chr3:107882510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107938422	+	chr3	107940958	+	.	4	14	1578342_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=1578342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_107922501_107947501_162C;SPAN=2536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:139 GQ:18.5 PL:[18.5, 0.0, 318.8] SR:14 DR:4 LR:-18.46 LO:34.54);ALT=G[chr3:107940958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	107976829	-	chr4	160636435	+	.	11	0	2300703_1	18.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2300703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:107976829(-)-4:160636435(-)__4_160622001_160647001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:0 DR:11 LR:-18.7 LO:24.04);ALT=[chr4:160636435[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	159642637	+	chr4	159644356	+	.	0	13	2297069_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2297069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_159642001_159667001_175C;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:99 GQ:16.1 PL:[16.1, 0.0, 224.0] SR:13 DR:0 LR:-16.09 LO:26.85);ALT=T[chr4:159644356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	160534324	+	chr4	160453026	+	.	17	0	2300181_1	46.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2300181_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:160453026(-)-4:160534324(+)__4_160524001_160549001D;SPAN=81298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:37 GQ:42.8 PL:[46.1, 0.0, 42.8] SR:0 DR:17 LR:-46.1 LO:46.1);ALT=]chr4:160534324]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	160453252	+	chr4	160534622	+	.	24	0	2300182_1	69.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=2300182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:160453252(+)-4:160534622(-)__4_160524001_160549001D;SPAN=81370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:22 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=T[chr4:160534622[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
