chr6	100537906	+	chr6	100539259	+	ATGAAAA	56	44	4336342_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=ATGAAAA;MAPQ=60;MATEID=4336342_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_100523501_100548501_78C;SPAN=1353;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:18 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:44 DR:56 LR:-247.6 LO:247.6);ALT=C[chr6:100539259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
