chrX	142798602	+	chrX	142600095	+	.	17	0	11409717_1	47.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=11409717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:142600095(-)-23:142798602(+)__23_142786001_142811001D;SPAN=198507;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:31 GQ:24.8 PL:[47.9, 0.0, 24.8] SR:0 DR:17 LR:-48.01 LO:48.01);ALT=]chrX:142798602]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	142600335	+	chrX	142798848	+	.	22	0	11409718_1	69.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=11409718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:142600335(+)-23:142798848(-)__23_142786001_142811001D;SPAN=198513;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:22 DP:26 GQ:3.6 PL:[69.3, 3.6, 0.0] SR:0 DR:22 LR:-70.32 LO:70.32);ALT=T[chrX:142798848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	142803366	+	chrX	144329491	-	.	12	0	11412678_1	28.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=11412678_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:142803366(+)-23:144329491(+)__23_144305001_144330001D;SPAN=1526125;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:41 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:0 DR:12 LR:-28.5 LO:29.51);ALT=T]chrX:144329491];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	142803642	-	chrX	144329202	+	.	23	0	11412679_1	62.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=11412679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:142803642(-)-23:144329202(-)__23_144305001_144330001D;SPAN=1525560;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:48 GQ:53 PL:[62.9, 0.0, 53.0] SR:0 DR:23 LR:-62.96 LO:62.96);ALT=[chrX:144329202[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	143406976	+	chrX	143409979	+	TAC	72	37	11411087_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TAC;MAPQ=60;MATEID=11411087_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_23_143398501_143423501_1C;SPAN=3003;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:19 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:37 DR:72 LR:-274.0 LO:274.0);ALT=A[chrX:143409979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	144422077	+	chrX	144424506	+	.	62	55	11412649_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=11412649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_144403001_144428001_160C;SPAN=2429;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:20 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:55 DR:62 LR:-283.9 LO:283.9);ALT=G[chrX:144424506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
