chr2	143635305	+	chr2	143642917	+	.	32	4	1025011_1	88.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1025011_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_143619001_143644001_247C;SPAN=7612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:76 GQ:88.4 PL:[88.4, 0.0, 95.0] SR:4 DR:32 LR:-88.34 LO:88.36);ALT=G[chr2:143642917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143635332	+	chr2	143676173	+	.	9	0	1025012_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1025012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:143635332(+)-2:143676173(-)__2_143619001_143644001D;SPAN=40841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=C[chr2:143676173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143643105	+	chr2	143676175	+	.	0	14	1025029_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1025029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_143619001_143644001_131C;SPAN=33070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:42 GQ:35 PL:[35.0, 0.0, 64.7] SR:14 DR:0 LR:-34.84 LO:35.4);ALT=G[chr2:143676175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143676298	+	chr2	143685228	+	.	2	8	1024906_1	8.0	.	DISC_MAPQ=33;EVDNC=ASDIS;MAPQ=60;MATEID=1024906_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_143668001_143693001_177C;SPAN=8930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:77 GQ:8.9 PL:[8.9, 0.0, 177.2] SR:8 DR:2 LR:-8.848 LO:18.1);ALT=T[chr2:143685228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143798227	+	chr2	143799616	+	.	0	7	1025091_1	5.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1025091_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_143790501_143815501_53C;SPAN=1389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:64 GQ:5.9 PL:[5.9, 0.0, 147.8] SR:7 DR:0 LR:-5.768 LO:13.86);ALT=T[chr2:143799616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143887036	+	chr2	143913044	+	.	91	9	1025408_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1025408_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_143913001_143938001_40C;SPAN=26008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:37 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:9 DR:91 LR:-274.0 LO:274.0);ALT=G[chr2:143913044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	143887075	+	chr2	143959702	+	.	13	0	1025620_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1025620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:143887075(+)-2:143959702(-)__2_143937501_143962501D;SPAN=72627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:39 GQ:32.3 PL:[32.3, 0.0, 62.0] SR:0 DR:13 LR:-32.35 LO:32.87);ALT=G[chr2:143959702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	144194611	+	chr2	144244942	+	.	2	2	1026121_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1026121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_144182501_144207501_16C;SPAN=50331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:34 GQ:4.1 PL:[4.1, 0.0, 76.7] SR:2 DR:2 LR:-3.993 LO:8.056);ALT=A[chr2:144244942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	144245064	+	chr2	144276833	+	.	2	4	1026204_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1026204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_144256001_144281001_166C;SPAN=31769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:31 GQ:11.6 PL:[11.6, 0.0, 61.1] SR:4 DR:2 LR:-11.41 LO:13.5);ALT=G[chr2:144276833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	145147598	+	chr2	145153978	+	.	10	5	1028110_1	20.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=9;MATEID=1028110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_145138001_145163001_41C;SPAN=6380;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:85 GQ:20 PL:[20.0, 0.0, 185.0] SR:5 DR:10 LR:-19.88 LO:27.78);ALT=G[chr2:145153978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	145187594	+	chr2	145274845	+	.	0	20	1028510_1	55.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1028510_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_145260501_145285501_203C;SPAN=87251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:38 GQ:35.9 PL:[55.7, 0.0, 35.9] SR:20 DR:0 LR:-55.94 LO:55.94);ALT=C[chr2:145274845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	145187595	+	chr2	145277506	+	TTGAATAACTTTTCTTCATCTGGTTTT	14	5	1028511_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTGAATAACTTTTCTTCATCTGGTTTT;MAPQ=60;MATEID=1028511_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_145260501_145285501_7C;SPAN=89911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:5 DR:14 LR:-33.8 LO:35.92);ALT=T[chr2:145277506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	145274988	+	chr2	145277506	+	.	55	51	1028560_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1028560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_145260501_145285501_45C;SPAN=2518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:80 DP:103 GQ:11.9 PL:[236.3, 0.0, 11.9] SR:51 DR:55 LR:-248.0 LO:248.0);ALT=T[chr2:145277506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
