chr8	77896433	+	chr8	77898423	+	.	0	8	3926899_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3926899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_77885501_77910501_262C;SPAN=1990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-2.025 LO:15.08);ALT=T[chr8:77898423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	77896474	+	chr8	77912254	+	.	10	0	3926900_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3926900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:77896474(+)-8:77912254(-)__8_77885501_77910501D;SPAN=15780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=A[chr8:77912254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	77898589	+	chr8	77912253	+	.	13	0	3926939_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3926939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:77898589(+)-8:77912253(-)__8_77910001_77935001D;SPAN=13664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:28 GQ:32 PL:[35.3, 0.0, 32.0] SR:0 DR:13 LR:-35.33 LO:35.33);ALT=T[chr8:77912253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
