chr8	117657345	+	chr8	117658709	+	.	0	55	4038095_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=4038095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117649001_117674001_81C;SPAN=1364;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:147 GQ:99 PL:[141.8, 0.0, 214.4] SR:55 DR:0 LR:-141.7 LO:142.6);ALT=G[chr8:117658709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117658844	+	chr8	117661045	+	.	8	7	4038101_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4038101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117649001_117674001_36C;SPAN=2201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:84 GQ:20.3 PL:[20.3, 0.0, 182.0] SR:7 DR:8 LR:-20.16 LO:27.85);ALT=T[chr8:117661045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117661168	+	chr8	117668095	+	.	8	16	4038110_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=4038110_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_117649001_117674001_288C;SPAN=6927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:94 GQ:37.4 PL:[37.4, 0.0, 189.2] SR:16 DR:8 LR:-37.25 LO:43.16);ALT=G[chr8:117668095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117661168	+	chr8	117669454	+	CTGGCAAGGCTGAGCAATTCATGTTTATCTGCAACAGCTGACTTCTTTTCAAGTTCCCACATTAGGACATTGATCAGATGTGAATTTTTAATTACAATCGGCACTTCTTCAAACATGTACTCAAAGGTGATATTTGCTTTTTTCAAT	7	26	4038111_1	75.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTGGCAAGGCTGAGCAATTCATGTTTATCTGCAACAGCTGACTTCTTTTCAAGTTCCCACATTAGGACATTGATCAGATGTGAATTTTTAATTACAATCGGCACTTCTTCAAACATGTACTCAAAGGTGATATTTGCTTTTTTCAAT;MAPQ=60;MATEID=4038111_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_117649001_117674001_288C;SPAN=8286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:76 GQ:75.2 PL:[75.2, 0.0, 108.2] SR:26 DR:7 LR:-75.14 LO:75.49);ALT=G[chr8:117669454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117668244	+	chr8	117669454	+	.	11	13	4038124_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=4038124_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_117649001_117674001_288C;SPAN=1210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:76 GQ:52.1 PL:[52.1, 0.0, 131.3] SR:13 DR:11 LR:-52.03 LO:53.97);ALT=T[chr8:117669454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117668280	+	chr8	117671049	+	.	10	0	4038125_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4038125_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:117668280(+)-8:117671049(-)__8_117649001_117674001D;SPAN=2769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:77 GQ:12.2 PL:[12.2, 0.0, 173.9] SR:0 DR:10 LR:-12.15 LO:20.6);ALT=T[chr8:117671049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117669554	+	chr8	117671052	+	.	7	19	4038127_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4038127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117649001_117674001_321C;SPAN=1498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:77 GQ:51.8 PL:[51.8, 0.0, 134.3] SR:19 DR:7 LR:-51.76 LO:53.82);ALT=C[chr8:117671052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117671221	+	chr8	117738255	+	.	15	40	4038279_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4038279_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117722501_117747501_194C;SPAN=67034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:78 GQ:44.9 PL:[143.9, 0.0, 44.9] SR:40 DR:15 LR:-146.7 LO:146.7);ALT=T[chr8:117738255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117671271	+	chr8	117767979	+	.	37	0	4038342_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4038342_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:117671271(+)-8:117767979(-)__8_117747001_117772001D;SPAN=96708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:70 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.6 LO:103.6);ALT=C[chr8:117767979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117779030	+	chr8	117782429	+	.	0	8	4038583_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4038583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117771501_117796501_324C;SPAN=3399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:8 DR:0 LR:0.9554 LO:14.66);ALT=G[chr8:117782429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117859924	+	chr8	117862855	+	.	8	0	4038673_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4038673_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:117859924(+)-8:117862855(-)__8_117845001_117870001D;SPAN=2931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=G[chr8:117862855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117861270	+	chr8	117862856	+	.	2	3	4038678_1	0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4038678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117845001_117870001_5C;SPAN=1586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:87 GQ:10.2 PL:[0.0, 10.2, 231.0] SR:3 DR:2 LR:10.37 LO:6.36);ALT=T[chr8:117862856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117864949	+	chr8	117866484	+	.	6	9	4038691_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4038691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117845001_117870001_289C;SPAN=1535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:75 GQ:26 PL:[26.0, 0.0, 154.7] SR:9 DR:6 LR:-25.89 LO:31.26);ALT=T[chr8:117866484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	117879002	+	chr8	117886848	+	.	0	15	4038757_1	28.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4038757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_117869501_117894501_234C;SPAN=7846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:79 GQ:28.1 PL:[28.1, 0.0, 163.4] SR:15 DR:0 LR:-28.11 LO:33.61);ALT=T[chr8:117886848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	118533292	+	chr8	118540888	+	.	0	8	4040151_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4040151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_118531001_118556001_228C;SPAN=7596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:8 DR:0 LR:0.4135 LO:14.74);ALT=G[chr8:118540888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	118873738	+	chr8	118875337	-	GAGATAGAGTC	27	24	4041232_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=GAGATAGAGTC;MAPQ=60;MATEID=4041232_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=TTTTTTTTTTT;SCTG=c_8_118874001_118899001_225C;SPAN=1599;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:38 GQ:12.4 PL:[60.7, 12.4, 0.0] SR:24 DR:27 LR:-60.73 LO:60.73);ALT=T]chr8:118875337];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	118873791	+	chr8	118875593	+	.	30	0	4041234_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4041234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:118873791(+)-8:118875593(-)__8_118874001_118899001D;SPAN=1802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:27 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=T[chr8:118875593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
