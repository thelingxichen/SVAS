chr8	19682485	+	chr8	19683935	+	.	3	4	3770052_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3770052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_19673501_19698501_209C;SPAN=1450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:89 GQ:4.2 PL:[0.0, 4.2, 224.4] SR:4 DR:3 LR:4.306 LO:10.56);ALT=T[chr8:19683935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	19689622	+	chr8	19690678	+	.	0	5	3770081_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3770081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_19673501_19698501_133C;SPAN=1056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:89 GQ:7.5 PL:[0.0, 7.5, 231.0] SR:5 DR:0 LR:7.607 LO:8.395);ALT=G[chr8:19690678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
