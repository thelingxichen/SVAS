chr19	27961383	+	chr19	27963247	+	.	57	43	6776166_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CTTTTACACCATAGGCCTCA;MAPQ=60;MATEID=6776166_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_19_27954501_27979501_104C;SPAN=1864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:54 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:43 DR:57 LR:-267.4 LO:267.4);ALT=A[chr19:27963247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	27976052	+	chr19	27979426	+	.	22	13	6776270_1	92.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGTTTGGAAACAATGTTTTTGTAGAATCTGTGAAGGGATATTT;MAPQ=60;MATEID=6776270_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_19_27979001_28004001_68C;SPAN=3374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:31 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:13 DR:22 LR:-92.42 LO:92.42);ALT=T[chr19:27979426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	28284565	+	chr19	28288659	+	.	8	0	6777659_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6777659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:28284565(+)-19:28288659(-)__19_28273001_28298001D;SPAN=4094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=C[chr19:28288659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
