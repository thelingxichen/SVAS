chr10	124134328	+	chr10	124152694	+	.	8	0	4708576_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4708576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:124134328(+)-10:124152694(-)__10_124141501_124166501D;SPAN=18366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:22 GQ:20.6 PL:[20.6, 0.0, 30.5] SR:0 DR:8 LR:-20.45 LO:20.61);ALT=G[chr10:124152694[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	124615305	+	chr10	124639001	+	.	10	4	4709458_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4709458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_124607001_124632001_34C;SPAN=23696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:26 GQ:26 PL:[26.0, 0.0, 35.9] SR:4 DR:10 LR:-25.97 LO:26.07);ALT=G[chr10:124639001[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	124921931	+	chr10	124923336	+	TTGGGTTTTGTTTCTGCATCTGTCACTTGGCGAATGAAGATACCATCTTCAGGATGTTCTGTGTCATCCATTTCATACATATATGATGACGCTATTGCAAGCGTAGTCCCATCATTACTGAAGGCAAGTGATGCGATGCTCGTGGGGTACCGATGGAATTGGCACAGTCGCTTTTTGTTAAATGGATCCCAAATATTTACAAAGCCATCAGAACC	0	15	4709875_1	35.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=TTGGGTTTTGTTTCTGCATCTGTCACTTGGCGAATGAAGATACCATCTTCAGGATGTTCTGTGTCATCCATTTCATACATATATGATGACGCTATTGCAAGCGTAGTCCCATCATTACTGAAGGCAAGTGATGCGATGCTCGTGGGGTACCGATGGAATTGGCACAGTCGCTTTTTGTTAAATGGATCCCAAATATTTACAAAGCCATCAGAACC;MAPQ=60;MATEID=4709875_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_124901001_124926001_33C;SPAN=1405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:15 DR:0 LR:-34.89 LO:36.48);ALT=T[chr10:124923336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
