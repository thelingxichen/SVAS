chr19	24494240	+	chr19	24485418	+	.	27	42	10230812_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TATCTG;MAPQ=60;MATEID=10230812_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_24475501_24500501_285C;SPAN=8822;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:56 DP:102 GQ:88.1 PL:[157.4, 0.0, 88.1] SR:42 DR:27 LR:-158.2 LO:158.2);ALT=]chr19:24494240]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	24485532	+	chr19	24494320	+	.	17	30	10230815_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGTAGAATCTGCGAAGTGATATTTGGGA;MAPQ=60;MATEID=10230815_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_24475501_24500501_215C;SPAN=8788;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:100 GQ:99 PL:[118.1, 0.0, 124.7] SR:30 DR:17 LR:-118.2 LO:118.2);ALT=A[chr19:24494320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24546085	+	chr19	24539642	+	.	135	79	10231385_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAAACTGCTTTGTGATG;MAPQ=60;MATEID=10231385_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_24524501_24549501_326C;SPAN=6443;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:181 DP:305 GQ:99 PL:[515.0, 0.0, 224.5] SR:79 DR:135 LR:-521.0 LO:521.0);ALT=]chr19:24546085]G;VARTYPE=BND:DUP-th;JOINTYPE=th
