chr13	89110970	+	chr13	89112881	-	ATATAATATTATATATATA	7	8	5589150_1	37.0	.	DISC_MAPQ=16;EVDNC=ASDIS;INSERTION=ATATAATATTATATATATA;MAPQ=25;MATEID=5589150_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_89106501_89131501_106C;SPAN=1911;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:44 GQ:37.7 PL:[37.7, 0.0, 67.4] SR:8 DR:7 LR:-37.59 LO:38.11);ALT=A]chr13:89112881];VARTYPE=BND:INV-hh;JOINTYPE=hh
