chr9	214978	+	chr9	271624	+	.	10	0	4122699_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4122699_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:214978(+)-9:271624(-)__9_196001_221001D;SPAN=56646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:0 DR:10 LR:-20.55 LO:23.07);ALT=T[chr9:271624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	215032	+	chr9	286461	+	TTCTTCAGTGGAAATAAGGAAACAGTTTACTCTCCCACCAAACCTTGGCCAGTACCATCGACAGAGCATAAGTACCTCTGGCTTCCCCTCTCTTCAACTA	0	19	4122701_1	50.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGTA;INSERTION=TTCTTCAGTGGAAATAAGGAAACAGTTTACTCTCCCACCAAACCTTGGCCAGTACCATCGACAGAGCATAAGTACCTCTGGCTTCCCCTCTCTTCAACTA;MAPQ=60;MATEID=4122701_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_9_196001_221001_271C;SPAN=71429;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:45 GQ:50.6 PL:[50.6, 0.0, 57.2] SR:19 DR:0 LR:-50.53 LO:50.56);ALT=A[chr9:286461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	312167	+	chr9	317041	+	.	0	7	4122566_1	6.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4122566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_294001_319001_110C;SPAN=4874;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:63 GQ:6.2 PL:[6.2, 0.0, 144.8] SR:7 DR:0 LR:-6.039 LO:13.91);ALT=G[chr9:317041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
