chr3	24298445	+	chr3	24159667	+	.	14	0	1896150_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1896150_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:24159667(-)-3:24298445(+)__3_24279501_24304501D;SPAN=138778;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:70 GQ:27.2 PL:[27.2, 0.0, 142.7] SR:0 DR:14 LR:-27.25 LO:31.73);ALT=]chr3:24298445]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	25030887	+	chr3	25032250	+	GGTGTAC	61	34	1898895_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GGTGTAC;MAPQ=60;MATEID=1898895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_25014501_25039501_351C;SPAN=1363;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:77 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:34 DR:61 LR:-227.8 LO:227.8);ALT=A[chr3:25032250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
