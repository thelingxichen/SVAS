chr9	28031835	+	chr9	28059140	-	AATAGT	24	24	4161253_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AATAGT;MAPQ=60;MATEID=4161253_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_28028001_28053001_229C;SPAN=27305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:16 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:24 DR:24 LR:-95.72 LO:95.72);ALT=A]chr9:28059140];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	28031863	-	chr9	28034467	+	TTTTCGGAATT	18	13	4161254_1	85.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TTTTCGGAATT;MAPQ=60;MATEID=4161254_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_28028001_28053001_57C;SPAN=2604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:34 GQ:2.4 PL:[85.8, 2.4, 0.0] SR:13 DR:18 LR:-88.56 LO:88.56);ALT=[chr9:28034467[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	28034286	+	chr9	28157692	+	TGACTATTTCAC	25	14	4161303_1	89.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TGACTATTTCAC;MAPQ=60;MATEID=4161303_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_28150501_28175501_135C;SPAN=123406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:19 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:14 DR:25 LR:-89.12 LO:89.12);ALT=C[chr9:28157692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
