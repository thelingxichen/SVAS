chr1	232708423	+	chr2	106986732	-	TATATATATAC	2	26	602590_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TATATATATAC;MAPQ=60;MATEID=602590_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_232701001_232726001_357C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:8 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:26 DR:2 LR:-82.52 LO:82.52);ALT=A]chr2:106986732];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	232896557	+	chr1	232891500	+	.	8	0	603253_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=603253_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:232891500(-)-1:232896557(+)__1_232872501_232897501D;SPAN=5057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:131 GQ:8.7 PL:[0.0, 8.7, 333.3] SR:0 DR:8 LR:9.083 LO:13.73);ALT=]chr1:232896557]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	233086491	+	chr1	233091301	+	.	23	12	603759_1	67.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=603759_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_233068501_233093501_241C;SPAN=4810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:105 GQ:67.4 PL:[67.4, 0.0, 186.2] SR:12 DR:23 LR:-67.28 LO:70.43);ALT=G[chr1:233091301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	233105866	+	chr1	233113909	+	.	3	7	603817_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=603817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_233093001_233118001_232C;SPAN=8043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:105 GQ:4.7 PL:[4.7, 0.0, 248.9] SR:7 DR:3 LR:-4.563 LO:19.17);ALT=T[chr1:233113909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	233707697	-	chr5	163685082	+	.	3	2	2631921_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCTTTTAT;MAPQ=60;MATEID=2631921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_163684501_163709501_50C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:17 GQ:11.9 PL:[11.9, 0.0, 28.4] SR:2 DR:3 LR:-11.9 LO:12.31);ALT=[chr5:163685082[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	106879557	+	chr2	106885916	+	GCCCAG	31	32	929748_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;INSERTION=GCCCAG;MAPQ=60;MATEID=929748_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_106869001_106894001_35C;SPAN=6359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:44 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:32 DR:31 LR:-148.5 LO:148.5);ALT=C[chr2:106885916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	162864810	+	chr5	162866261	+	.	0	11	2630745_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2630745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_162851501_162876501_124C;SPAN=1451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:59 GQ:20.3 PL:[20.3, 0.0, 122.6] SR:11 DR:0 LR:-20.33 LO:24.55);ALT=G[chr5:162866261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	162884088	+	chr5	162886868	+	.	10	2	2630873_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2630873_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_162876001_162901001_228C;SPAN=2780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:72 GQ:20.3 PL:[20.3, 0.0, 152.3] SR:2 DR:10 LR:-20.11 LO:26.14);ALT=T[chr5:162886868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	162930443	+	chr5	162939005	+	.	8	0	2630961_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2630961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:162930443(+)-5:162939005(-)__5_162925001_162950001D;SPAN=8562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=A[chr5:162939005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	162932756	+	chr5	162939006	+	.	23	7	2630966_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2630966_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_162925001_162950001_185C;SPAN=6250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:52 GQ:52.1 PL:[71.9, 0.0, 52.1] SR:7 DR:23 LR:-71.86 LO:71.86);ALT=G[chr5:162939006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	162939202	+	chr5	162940559	+	.	4	7	2630979_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2630979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_162925001_162950001_35C;SPAN=1357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:7 DR:4 LR:-17.52 LO:20.4);ALT=G[chr5:162940559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	163579919	+	chr5	163604217	-	.	15	9	2631975_1	62.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GGAGCTAAATGATGAGAACTTATGAACACAAAGAAGGAAACAACAG;MAPQ=60;MATEID=2631975_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_163586501_163611501_228C;SPAN=24298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:37 GQ:26.3 PL:[62.6, 0.0, 26.3] SR:9 DR:15 LR:-63.36 LO:63.36);ALT=G]chr5:163604217];VARTYPE=BND:INV-hh;JOINTYPE=hh
