chr17	51852805	+	chr17	51860708	+	.	24	0	6434238_1	68.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=6434238_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:51852805(+)-17:51860708(-)__17_51842001_51867001D;SPAN=7903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:42 GQ:31.7 PL:[68.0, 0.0, 31.7] SR:0 DR:24 LR:-68.45 LO:68.45);ALT=T[chr17:51860708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
