chr10	81787050	+	chr10	81793402	+	.	9	0	6388938_1	0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6388938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:81787050(+)-10:81793402(-)__10_81781001_81806001D;SPAN=6352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:113 GQ:0.6 PL:[0.0, 0.6, 273.9] SR:0 DR:9 LR:0.9055 LO:16.52);ALT=G[chr10:81793402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	82295404	+	chr16	75503315	+	.	35	0	9423482_1	99.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=9423482_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:82295404(+)-16:75503315(-)__16_75484501_75509501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:23 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:35 LR:-102.3 LO:102.3);ALT=G[chr16:75503315[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	82750298	+	chr10	82752650	+	.	65	52	6393535_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=6393535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_82736501_82761501_303C;SPAN=2352;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:107 GQ:28.8 PL:[316.8, 28.8, 0.0] SR:52 DR:65 LR:-316.0 LO:316.0);ALT=G[chr10:82752650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	73392080	-	chr16	73393283	+	.	2	2	9410751_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCCCCAG;MAPQ=60;MATEID=9410751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_73377501_73402501_274C;SPAN=1203;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:166 GQ:31.6 PL:[0.0, 31.6, 465.4] SR:2 DR:2 LR:31.77 LO:5.232);ALT=[chr16:73393283[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	73868574	+	chr16	73869693	-	.	8	0	9413091_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9413091_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:73868574(+)-16:73869693(+)__16_73843001_73868001D;SPAN=1119;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:8 DP:0 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=G]chr16:73869693];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	75190857	+	chr16	74698063	+	.	96	29	9422046_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=9422046_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75166001_75191001_65C;SPAN=492794;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:109 DP:72 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:29 DR:96 LR:-323.5 LO:323.5);ALT=]chr16:75190857]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	75523308	+	chr16	75418894	+	.	9	0	9423044_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=9423044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:75418894(-)-16:75523308(+)__16_75509001_75534001D;SPAN=104414;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-15.89 LO:19.85);ALT=]chr16:75523308]T;VARTYPE=BND:DUP-th;JOINTYPE=th
