chr1	243127797	+	chr1	243129216	+	.	48	62	638158_1	99.0	.	DISC_MAPQ=14;EVDNC=ASDIS;HOMSEQ=GCCTCCCAAAGTGCTGGGATTACAGG;MAPQ=60;MATEID=638158_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_1_243113501_243138501_253C;SPAN=1419;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:15 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:62 DR:48 LR:-287.2 LO:287.2);ALT=G[chr1:243129216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	243385118	+	chr1	243388478	+	.	4	9	638930_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=638930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_243383001_243408001_144C;SPAN=3360;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:103 GQ:5.3 PL:[5.3, 0.0, 242.9] SR:9 DR:4 LR:-5.105 LO:19.26);ALT=G[chr1:243388478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	243419544	+	chr1	243433393	+	.	26	6	639256_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=639256_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_243432001_243457001_190C;SPAN=13849;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:63 GQ:65.6 PL:[85.4, 0.0, 65.6] SR:6 DR:26 LR:-85.37 LO:85.37);ALT=T[chr1:243433393[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
