chr5	11438206	+	chr5	11445528	+	.	13	38	3210297_1	86.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3210297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_11441501_11466501_373C;SPAN=7322;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:170 GQ:86 PL:[86.0, 0.0, 326.9] SR:38 DR:13 LR:-85.98 LO:93.88);ALT=G[chr5:11445528[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
