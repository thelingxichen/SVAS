chr4	135433002	+	chr4	135435702	+	GTACA	85	44	2932787_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GTACA;MAPQ=60;MATEID=2932787_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_4_135436001_135461001_313C;SPAN=2700;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:0 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:44 DR:85 LR:-326.8 LO:326.8);ALT=A[chr4:135435702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
