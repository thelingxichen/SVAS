chr3	146251337	+	chr3	146262254	+	TTTGTTTGTCCATGATTAAAACAGTT	0	12	1707241_1	12.0	.	EVDNC=ASSMB;INSERTION=TTTGTTTGTCCATGATTAAAACAGTT;MAPQ=60;MATEID=1707241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_146240501_146265501_330C;SPAN=10917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:99 GQ:12.8 PL:[12.8, 0.0, 227.3] SR:12 DR:0 LR:-12.79 LO:24.33);ALT=T[chr3:146262254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	146385190	+	chr3	146394862	+	.	43	29	1707604_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=1707604_2;MATENM=2;NM=4;NUMPARTS=2;SCTG=c_3_146387501_146412501_217C;SPAN=9672;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:81 GQ:8 PL:[186.2, 0.0, 8.0] SR:29 DR:43 LR:-195.4 LO:195.4);ALT=A[chr3:146394862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	146395165	+	chr3	146390405	+	ATTGGGGAG	60	34	1707614_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=ATTGGGGAG;MAPQ=60;MATEID=1707614_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_3_146387501_146412501_195C;SPAN=4760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:85 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:34 DR:60 LR:-250.9 LO:250.9);ALT=]chr3:146395165]A;VARTYPE=BND:DUP-th;JOINTYPE=th
