chr9	45130257	+	chr9	45128907	+	.	55	0	5853670_1	99.0	.	DISC_MAPQ=7;EVDNC=DSCRD;IMPRECISE;MAPQ=7;MATEID=5853670_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:45128907(-)-9:45130257(+)__9_45129001_45154001D;SPAN=1350;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:55 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:55 LR:-161.7 LO:161.7);ALT=]chr9:45130257]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	45579542	+	chr11	101760182	+	.	6	19	5855020_1	59.0	.	DISC_MAPQ=8;EVDNC=ASDIS;HOMSEQ=AAAGAAAGAAAGAGAAAGAAAGAAAAAGAAAGAA;MAPQ=16;MATEID=5855020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_45570001_45595001_168C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:20 DP:25 GQ:0 PL:[59.4, 0.0, 0.0] SR:19 DR:6 LR:-62.61 LO:62.61);ALT=A[chr11:101760182[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	101977277	+	chr11	102078986	+	.	0	48	7162536_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AT;MAPQ=60;MATEID=7162536_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_11_102067001_102092001_47C;SPAN=101709;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:48 DP:10 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:48 DR:0 LR:-141.9 LO:141.9);ALT=T[chr11:102078986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	102608901	+	chr11	102610276	-	.	4	3	7163901_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTATATTTGGAAAAA;MAPQ=60;MATEID=7163901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_102606001_102631001_139C;SPAN=1375;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:6 DP:69 GQ:1.1 PL:[1.1, 0.0, 166.1] SR:3 DR:4 LR:-1.112 LO:11.25);ALT=A]chr11:102610276];VARTYPE=BND:INV-hh;JOINTYPE=hh
