chr11	7790354	+	chr11	7791978	+	.	40	0	6634503_1	99.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=6634503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:7790354(+)-11:7791978(-)__11_7791001_7816001D;SPAN=1624;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:40 DP:2 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:40 LR:-118.8 LO:118.8);ALT=C[chr11:7791978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
