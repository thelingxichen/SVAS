chr13	101894146	+	chr13	101896425	+	.	125	72	5623472_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CAT;MAPQ=60;MATEID=5623472_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_13_101871001_101896001_113C;SPAN=2279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:163 DP:14 GQ:43.9 PL:[481.9, 43.9, 0.0] SR:72 DR:125 LR:-481.9 LO:481.9);ALT=T[chr13:101896425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
