chr7	12251051	+	chr7	12254434	+	.	9	3	3171178_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3171178_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_12250001_12275001_61C;SPAN=3383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:3 DR:9 LR:-6.73 LO:19.53);ALT=G[chr7:12254434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
