chr18	48530709	+	chr18	48700866	+	.	82	66	10018307_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACTA;MAPQ=60;MATEID=10018307_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_48510001_48535001_59C;SPAN=170157;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:117 DP:8 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:66 DR:82 LR:-346.6 LO:346.6);ALT=A[chr18:48700866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	49196735	+	chr18	49198874	+	CG	85	66	10019406_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=CG;MAPQ=60;MATEID=10019406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_49196001_49221001_4C;SPAN=2139;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:138 DP:25 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:66 DR:85 LR:-409.3 LO:409.3);ALT=G[chr18:49198874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
