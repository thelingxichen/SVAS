chr10	58119939	+	chr10	58120955	+	.	19	0	4603923_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4603923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:58119939(+)-10:58120955(-)__10_58114001_58139001D;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:57 GQ:47.3 PL:[47.3, 0.0, 90.2] SR:0 DR:19 LR:-47.28 LO:48.04);ALT=A[chr10:58120955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
