chr3	25030887	+	chr3	25032250	+	GGTGTAC	0	23	1307653_1	22.0	.	EVDNC=ASSMB;INSERTION=GGTGTAC;MAPQ=60;MATEID=1307653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_25014501_25039501_664C;SPAN=1363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:196 GQ:22.9 PL:[22.9, 0.0, 452.0] SR:23 DR:0 LR:-22.82 LO:46.29);ALT=A[chr3:25032250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	25640003	+	chr3	25642596	+	.	10	0	1311878_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1311878_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:25640003(+)-3:25642596(-)__3_25627001_25652001D;SPAN=2593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:188 GQ:17.8 PL:[0.0, 17.8, 491.8] SR:0 DR:10 LR:17.92 LO:16.55);ALT=A[chr3:25642596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	25642717	+	chr3	25646250	+	.	3	6	1311902_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1311902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_25627001_25652001_14C;SPAN=3533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:223 GQ:33.7 PL:[0.0, 33.7, 607.3] SR:6 DR:3 LR:34.01 LO:11.85);ALT=C[chr3:25646250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	25657079	+	chr3	25659908	+	.	2	3	1312336_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1312336_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_25651501_25676501_130C;SPAN=2829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:183 GQ:36.1 PL:[0.0, 36.1, 514.9] SR:3 DR:2 LR:36.38 LO:5.063);ALT=T[chr3:25659908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	25820183	+	chr3	25824751	+	.	0	9	1313293_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CTGA;MAPQ=60;MATEID=1313293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_25823001_25848001_81C;SPAN=4568;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:9 DR:0 LR:-7.222 LO:17.79);ALT=A[chr3:25824751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	26450970	+	chr3	26452299	+	.	232	146	1317799_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1317799_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_26435501_26460501_389C;SPAN=1329;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:300 DP:114 GQ:81.2 PL:[891.2, 81.2, 0.0] SR:146 DR:232 LR:-891.2 LO:891.2);ALT=T[chr3:26452299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
