chr18	7146700	+	chr18	7144405	+	.	46	26	9881143_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=ACCTGTAATCCCAGCTACTAGGGAGGCTGAGGCAGGAGA;MAPQ=60;MATEID=9881143_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_18_7129501_7154501_77C;SPAN=2295;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:67 DP:141 GQ:99 PL:[183.2, 0.0, 156.8] SR:26 DR:46 LR:-183.1 LO:183.1);ALT=]chr18:7146700]A;VARTYPE=BND:DUP-th;JOINTYPE=th
