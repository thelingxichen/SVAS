chr4	144158629	-	chr4	144159712	+	.	8	0	2965089_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=2965089_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:144158629(-)-4:144159712(-)__4_144158001_144183001D;SPAN=1083;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:0 DR:8 LR:5.561 LO:14.1);ALT=[chr4:144159712[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
