chr13	70918113	-	chr13	70920284	+	.	3	2	8140112_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTTCTCAAAATAT;MAPQ=60;MATEID=8140112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_70903001_70928001_355C;SPAN=2171;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:132 GQ:22.2 PL:[0.0, 22.2, 363.0] SR:2 DR:3 LR:22.56 LO:5.629);ALT=[chr13:70920284[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
