chr7	148072866	+	chr7	148076324	+	.	40	37	3681957_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=ATC;MAPQ=60;MATEID=3681957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_148053501_148078501_338C;SPAN=3458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:72 GQ:0.5 PL:[172.1, 0.0, 0.5] SR:37 DR:40 LR:-182.0 LO:182.0);ALT=C[chr7:148076324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	148178646	+	chr13	98695060	-	.	17	42	3682597_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3682597_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_7_148176001_148201001_26C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:63 GQ:6.9 PL:[165.0, 6.9, 0.0] SR:42 DR:17 LR:-169.0 LO:169.0);ALT=G]chr13:98695060];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	148396117	+	chr7	148427062	+	.	10	0	3683278_1	20.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3683278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:148396117(+)-7:148427062(-)__7_148421001_148446001D;SPAN=30945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=T[chr7:148427062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	148670131	+	chr7	148676766	+	.	64	24	3684165_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CTCTACTAAAAATACAAAAATTAGCT;MAPQ=60;MATEID=3684165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_148666001_148691001_27C;SPAN=6635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:51 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:24 DR:64 LR:-247.6 LO:247.6);ALT=T[chr7:148676766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	148718240	+	chr7	148725413	+	.	14	10	3684468_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3684468_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_148715001_148740001_48C;SPAN=7173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:98 GQ:29.6 PL:[29.6, 0.0, 207.8] SR:10 DR:14 LR:-29.57 LO:37.35);ALT=C[chr7:148725413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	97627470	+	chr13	97632693	+	.	43	36	5610808_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGCT;MAPQ=60;MATEID=5610808_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_97632501_97657501_195C;SPAN=5223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:31 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:36 DR:43 LR:-194.7 LO:194.7);ALT=T[chr13:97632693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	98629041	+	chr13	98634755	+	.	5	5	5613399_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5613399_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_98612501_98637501_285C;SPAN=5714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:5 DR:5 LR:-10.15 LO:16.58);ALT=G[chr13:98634755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
