chr4	61330106	+	chr4	61333187	+	G	78	97	1992388_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=1992388_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_4_61323501_61348501_162C;SPAN=3081;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:164 DP:33 GQ:44.2 PL:[485.2, 44.2, 0.0] SR:97 DR:78 LR:-485.2 LO:485.2);ALT=T[chr4:61333187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	61939191	+	chr4	61942244	+	.	48	39	1993829_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=1993829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_61936001_61961001_16C;SPAN=3053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:61 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:39 DR:48 LR:-208.0 LO:208.0);ALT=A[chr4:61942244[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
