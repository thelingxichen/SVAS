chr7	51594312	+	chr7	51598690	+	CTGCA	139	55	4804747_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CTGCA;MAPQ=60;MATEID=4804747_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_51597001_51622001_299C;SPAN=4378;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:176 DP:59 GQ:47.5 PL:[521.5, 47.5, 0.0] SR:55 DR:139 LR:-521.5 LO:521.5);ALT=G[chr7:51598690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
