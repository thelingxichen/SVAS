chr1	105428616	+	chr18	68438274	+	.	2	14	257019_1	49.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=A;MAPQ=18;MATEID=257019_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_105423501_105448501_124C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:17 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:14 DR:2 LR:-49.51 LO:49.51);ALT=A[chr18:68438274[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr18	68383843	+	chr18	68405438	+	.	17	0	6666933_1	41.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6666933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:68383843(+)-18:68405438(-)__18_68404001_68429001D;SPAN=21595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:54 GQ:41.6 PL:[41.6, 0.0, 87.8] SR:0 DR:17 LR:-41.49 LO:42.46);ALT=A[chr18:68405438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	68405811	+	chr18	68387250	+	TATTCACG	45	42	6666935_1	99.0	.	DISC_MAPQ=28;EVDNC=ASDIS;INSERTION=TATTCACG;MAPQ=60;MATEID=6666935_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_68404001_68429001_274C;SPAN=18561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:47 GQ:21 PL:[231.0, 21.0, 0.0] SR:42 DR:45 LR:-231.1 LO:231.1);ALT=]chr18:68405811]A;VARTYPE=BND:DUP-th;JOINTYPE=th
