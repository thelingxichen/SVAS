chr2	122368979	+	chr2	122367896	+	.	19	0	1304184_1	27.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=1304184_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:122367896(-)-2:122368979(+)__2_122353001_122378001D;SPAN=1083;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:131 GQ:27.5 PL:[27.5, 0.0, 288.2] SR:0 DR:19 LR:-27.23 LO:40.13);ALT=]chr2:122368979]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	122483129	+	chr2	122484253	-	.	2	2	1304553_1	0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=TGGGCGTGGTGG;MAPQ=60;MATEID=1304553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_122475501_122500501_264C;SPAN=1124;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:123 GQ:19.8 PL:[0.0, 19.8, 336.6] SR:2 DR:2 LR:20.12 LO:5.753);ALT=G]chr2:122484253];VARTYPE=BND:INV-hh;JOINTYPE=hh
