chr8	59465906	+	chr8	59484762	+	.	23	0	3876928_1	48.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3876928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:59465906(+)-8:59484762(-)__8_59461501_59486501D;SPAN=18856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:100 GQ:48.8 PL:[48.8, 0.0, 194.0] SR:0 DR:23 LR:-48.83 LO:53.72);ALT=C[chr8:59484762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	59465906	+	chr8	59483440	+	.	19	0	3876927_1	37.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3876927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:59465906(+)-8:59483440(-)__8_59461501_59486501D;SPAN=17534;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:94 GQ:37.4 PL:[37.4, 0.0, 189.2] SR:0 DR:19 LR:-37.25 LO:43.16);ALT=C[chr8:59483440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	59483524	+	chr8	59484764	+	.	0	36	3876977_1	92.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3876977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_59461501_59486501_321C;SPAN=1240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:98 GQ:92.3 PL:[92.3, 0.0, 145.1] SR:36 DR:0 LR:-92.29 LO:92.94);ALT=A[chr8:59484764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	59484873	+	chr8	59488458	+	.	3	14	3876979_1	44.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3876979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_59461501_59486501_59C;SPAN=3585;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:14 DR:3 LR:-44.2 LO:44.37);ALT=G[chr8:59488458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	60136747	+	chr8	60135407	+	.	172	25	3878877_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCTACTTGGGAGGCTGAGGCAGGAGAATTGCTTGAACCCGGGAGGTAGAGGTTTCAGTGAGCCAAGATC;MAPQ=60;MATEID=3878877_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_8_60123001_60148001_335C;SPAN=1340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:189 DP:120 GQ:51.1 PL:[561.1, 51.1, 0.0] SR:25 DR:172 LR:-561.1 LO:561.1);ALT=]chr8:60136747]G;VARTYPE=BND:DUP-th;JOINTYPE=th
