chr2	39962238	+	chr2	39580021	+	.	67	48	970935_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=970935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_39959501_39984501_56C;SPAN=382217;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:96 DP:45 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:48 DR:67 LR:-283.9 LO:283.9);ALT=]chr2:39962238]A;VARTYPE=BND:DUP-th;JOINTYPE=th
