chr7	156752475	+	chr7	156630824	+	.	10	7	5353784_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=5353784_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_156751001_156776001_204C;SPAN=121651;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:50 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:7 DR:10 LR:-29.37 LO:31.17);ALT=]chr7:156752475]T;VARTYPE=BND:DUP-th;JOINTYPE=th
