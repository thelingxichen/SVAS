chr6	99850587	+	chr6	99852479	+	GAGTCCAGTGAGGGAAGCCAGTGCACTGGACTGTGCCAGCTGTTTTGCAGGAG	0	18	2957070_1	33.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTTT;INSERTION=GAGTCCAGTGAGGGAAGCCAGTGCACTGGACTGTGCCAGCTGTTTTGCAGGAG;MAPQ=60;MATEID=2957070_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_99837501_99862501_127C;SPAN=1892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:95 GQ:33.8 PL:[33.8, 0.0, 195.5] SR:18 DR:0 LR:-33.68 LO:40.32);ALT=C[chr6:99852479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99852579	+	chr6	99853907	+	.	0	14	2957076_1	26.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2957076_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99837501_99862501_149C;SPAN=1328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:14 DR:0 LR:-26.71 LO:31.54);ALT=C[chr6:99853907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99854044	+	chr6	99855956	+	.	14	9	2957081_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2957081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99837501_99862501_134C;SPAN=1912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:71 GQ:40.4 PL:[40.4, 0.0, 129.5] SR:9 DR:14 LR:-40.18 LO:42.93);ALT=C[chr6:99855956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99856148	+	chr6	99858617	+	AATTTGTGGAGGCTCCTGCTTCACAGGAAGTGCAATAGGTGAACGCTGACGATCCCTGAATGATGATGGCCTTTCTCTTCGATTCTGGGGAGGTGCTGGAGGTCCTGGAGGTCCTGGTTGCCAATAAGGAGGATGAAATCCACCTTGCGGTGGACCAAAAGCAGCCCCATG	0	44	2957087_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTGA;INSERTION=AATTTGTGGAGGCTCCTGCTTCACAGGAAGTGCAATAGGTGAACGCTGACGATCCCTGAATGATGATGGCCTTTCTCTTCGATTCTGGGGAGGTGCTGGAGGTCCTGGAGGTCCTGGTTGCCAATAAGGAGGATGAAATCCACCTTGCGGTGGACCAAAAGCAGCCCCATG;MAPQ=60;MATEID=2957087_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_99837501_99862501_210C;SPAN=2469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:87 GQ:88.7 PL:[121.7, 0.0, 88.7] SR:44 DR:0 LR:-121.9 LO:121.9);ALT=C[chr6:99858617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99857224	+	chr6	99858617	+	.	6	24	2957088_1	71.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTGA;MAPQ=60;MATEID=2957088_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_99837501_99862501_210C;SPAN=1393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:88 GQ:71.9 PL:[71.9, 0.0, 141.2] SR:24 DR:6 LR:-71.89 LO:73.14);ALT=A[chr6:99858617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99858842	+	chr6	99860427	+	.	8	7	2957089_1	17.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2957089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99837501_99862501_141C;SPAN=1585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:84 GQ:17 PL:[17.0, 0.0, 185.3] SR:7 DR:8 LR:-16.85 LO:25.26);ALT=T[chr6:99860427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99860615	+	chr6	99862447	+	.	0	61	2957100_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2957100_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99837501_99862501_292C;SPAN=1832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:112 GQ:98.6 PL:[171.2, 0.0, 98.6] SR:61 DR:0 LR:-172.0 LO:172.0);ALT=C[chr6:99862447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99860664	+	chr6	99873089	+	.	36	0	2957101_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2957101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:99860664(+)-6:99873089(-)__6_99837501_99862501D;SPAN=12425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:36 LR:-118.8 LO:118.8);ALT=A[chr6:99873089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99862568	+	chr6	99864225	+	.	0	52	2956951_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2956951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99862001_99887001_37C;SPAN=1657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:97 GQ:89.3 PL:[145.4, 0.0, 89.3] SR:52 DR:0 LR:-146.1 LO:146.1);ALT=T[chr6:99864225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99862600	+	chr6	99873089	+	.	94	0	2957107_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2957107_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:99862600(+)-6:99873089(-)__6_99837501_99862501D;SPAN=10489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:0 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:0 DR:94 LR:-277.3 LO:277.3);ALT=G[chr6:99873089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	99864305	+	chr6	99873090	+	.	22	12	2956956_1	57.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2956956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_99862001_99887001_129C;SPAN=8785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:93 GQ:57.5 PL:[57.5, 0.0, 166.4] SR:12 DR:22 LR:-57.33 LO:60.37);ALT=C[chr6:99873090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	100010872	+	chr6	100016435	+	.	9	0	2957481_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2957481_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:100010872(+)-6:100016435(-)__6_100009001_100034001D;SPAN=5563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:0 DR:9 LR:-9.661 LO:18.26);ALT=C[chr6:100016435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
