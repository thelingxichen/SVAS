chr6	16788869	+	chr1	167076422	+	.	9	0	4048793_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4048793_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167076422(-)-6:16788869(+)__6_16782501_16807501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=]chr6:16788869]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	167866793	+	chr21	28927095	-	.	15	0	617433_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=617433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167866793(+)-21:28927095(+)__1_167849501_167874501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:0 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=A]chr21:28927095];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	168186186	-	chr1	182274316	+	AAAAAAAAAAAA	49	32	678072_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=AAAAAAAAAAAA;MAPQ=60;MATEID=678072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_182255501_182280501_276C;SPAN=14088130;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:42 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:32 DR:49 LR:-184.8 LO:184.8);ALT=[chr1:182274316[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	168186489	+	chr3	53175885	+	T	28	43	2024289_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=2024289_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_53165001_53190001_86C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:82 GQ:47.3 PL:[149.6, 0.0, 47.3] SR:43 DR:28 LR:-152.2 LO:152.2);ALT=T[chr3:53175885[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	168427011	+	chr1	168428843	+	CTTTCTCTTCTTT	48	34	619349_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=CTTTCTCTTCTTT;MAPQ=60;MATEID=619349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_168413001_168438001_40C;SPAN=1832;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:68 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:34 DR:48 LR:-201.3 LO:201.3);ALT=T[chr1:168428843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168546426	+	chr1	168548123	+	.	16	0	619861_1	5.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=619861_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:168546426(+)-1:168548123(-)__1_168535501_168560501D;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:174 GQ:5.8 PL:[5.8, 0.0, 415.1] SR:0 DR:16 LR:-5.675 LO:30.41);ALT=T[chr1:168548123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169249699	+	chr1	169243686	+	.	16	0	624015_1	32.0	.	DISC_MAPQ=11;EVDNC=DSCRD;IMPRECISE;MAPQ=11;MATEID=624015_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169243686(-)-1:169249699(+)__1_169221501_169246501D;SPAN=6013;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:77 GQ:32 PL:[32.0, 0.0, 154.1] SR:0 DR:16 LR:-31.96 LO:36.56);ALT=]chr1:169249699]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr21	23626258	+	chr21	29293614	-	.	33	0	10738679_1	89.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=10738679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:23626258(+)-21:29293614(+)__21_29277501_29302501D;SPAN=5667356;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:33 DP:72 GQ:83 PL:[89.6, 0.0, 83.0] SR:0 DR:33 LR:-89.43 LO:89.43);ALT=T]chr21:29293614];VARTYPE=BND:INV-hh;JOINTYPE=hh
