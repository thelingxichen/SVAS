chr5	20557824	+	chr5	20536718	+	.	69	28	3268302_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=3268302_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_20555501_20580501_13C;SPAN=21106;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:86 GQ:16.5 PL:[240.9, 16.5, 0.0] SR:28 DR:69 LR:-242.9 LO:242.9);ALT=]chr5:20557824]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	21431000	+	chr5	21432223	+	GCTG	0	52	3274354_1	99.0	.	EVDNC=ASSMB;INSERTION=GCTG;MAPQ=60;MATEID=3274354_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_21413001_21438001_220C;SPAN=1223;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:157 GQ:99 PL:[129.2, 0.0, 251.3] SR:52 DR:0 LR:-129.1 LO:131.3);ALT=G[chr5:21432223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
