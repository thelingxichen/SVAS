chr9	26935207	+	chr9	26946895	+	.	0	7	4159599_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4159599_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_26925501_26950501_97C;SPAN=11688;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:7 DR:0 LR:-2.246 LO:13.27);ALT=G[chr9:26946895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	26962085	+	chr9	26978126	+	.	2	9	4159751_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4159751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_26950001_26975001_70C;SPAN=16041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:9 DR:2 LR:-22.39 LO:22.75);ALT=A[chr9:26978126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
