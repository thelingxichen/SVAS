chr4	120263656	+	chr4	120264670	+	.	12	0	2875101_1	14.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2875101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:120263656(+)-4:120264670(-)__4_120246001_120271001D;SPAN=1014;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:95 GQ:14 PL:[14.0, 0.0, 215.3] SR:0 DR:12 LR:-13.87 LO:24.56);ALT=A[chr4:120264670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	120602312	-	chr22	42181904	+	TAAATA	7	24	10896387_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TAAATA;MAPQ=60;MATEID=10896387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42164501_42189501_207C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:49 GQ:42.8 PL:[75.8, 0.0, 42.8] SR:24 DR:7 LR:-76.34 LO:76.34);ALT=[chr22:42181904[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	120963567	+	chr4	120965120	+	.	78	49	2878014_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=AGTT;MAPQ=0;MATEID=2878014_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_4_120956501_120981501_8C;SECONDARY;SPAN=1553;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:103 DP:86 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:49 DR:78 LR:-303.7 LO:303.7);ALT=T[chr4:120965120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
