chr16	82183010	+	chr16	82197686	+	CAACCTCAGGATTAAATCCTCTGAATGACATTCTTCCATAGAGAAGATCTTCACATAGTAAGAAACTCTGCTCTTCTATTATGAAACT	2	14	6262698_1	28.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CAACCTCAGGATTAAATCCTCTGAATGACATTCTTCCATAGAGAAGATCTTCACATAGTAAGAAACTCTGCTCTTCTATTATGAAACT;MAPQ=60;MATEID=6262698_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_82173001_82198001_126C;SPAN=14676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:14 DR:2 LR:-28.06 LO:32.03);ALT=T[chr16:82197686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	82185167	+	chr16	82203729	+	.	9	0	6262700_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6262700_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:82185167(+)-16:82203729(-)__16_82173001_82198001D;SPAN=18562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:20 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.29 LO:24.29);ALT=A[chr16:82203729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	82197812	+	chr16	82203729	+	.	10	0	6262715_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6262715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:82197812(+)-16:82203729(-)__16_82173001_82198001D;SPAN=5917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:0 DR:10 LR:-26.24 LO:26.3);ALT=A[chr16:82203729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
