chr2	158290989	+	chr2	158300450	+	.	10	0	1057480_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1057480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:158290989(+)-2:158300450(-)__2_158270001_158295001D;SPAN=9461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=T[chr2:158300450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	158291310	+	chr2	158300436	+	.	22	0	1057483_1	64.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1057483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:158291310(+)-2:158300436(-)__2_158270001_158295001D;SPAN=9126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:29 GQ:5.3 PL:[64.7, 0.0, 5.3] SR:0 DR:22 LR:-67.69 LO:67.69);ALT=G[chr2:158300436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
