chr12	4398157	+	chr12	4409025	+	.	3	7	5074526_1	8.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5074526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_4385501_4410501_115C;SPAN=10868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:7 DR:3 LR:-8.035 LO:17.94);ALT=G[chr12:4409025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4648156	+	chr12	4652927	+	.	11	0	5075225_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5075225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:4648156(+)-12:4652927(-)__12_4630501_4655501D;SPAN=4771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:79 GQ:14.9 PL:[14.9, 0.0, 176.6] SR:0 DR:11 LR:-14.91 LO:23.02);ALT=G[chr12:4652927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4714252	+	chr12	4719319	+	.	25	9	5075377_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5075377_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_4704001_4729001_30C;SPAN=5067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:99 GQ:55.7 PL:[55.7, 0.0, 184.4] SR:9 DR:25 LR:-55.7 LO:59.57);ALT=G[chr12:4719319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4719450	+	chr12	4721709	+	.	0	11	5075388_1	13.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5075388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_4704001_4729001_326C;SPAN=2259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:11 DR:0 LR:-13.28 LO:22.64);ALT=T[chr12:4721709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4758343	+	chr12	4763458	+	.	40	4	5076596_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=5076596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_4753001_4778001_227C;SPAN=5115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:81 GQ:80.6 PL:[113.6, 0.0, 80.6] SR:4 DR:40 LR:-113.6 LO:113.6);ALT=T[chr12:4763458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4758368	+	chr12	4763989	+	.	8	0	5076598_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5076598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:4758368(+)-12:4763989(-)__12_4753001_4778001D;SPAN=5621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=C[chr12:4763989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4763629	+	chr12	4766913	+	ACGCATGGGGTCACAGGTAATCATACCCTATCGGTGTGATAAATATGACATCATGCACCTTCGTCCCATGGGTGACCTGGGCCAGCTTCTGTTTCT	0	54	5076617_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ACGCATGGGGTCACAGGTAATCATACCCTATCGGTGTGATAAATATGACATCATGCACCTTCGTCCCATGGGTGACCTGGGCCAGCTTCTGTTTCT;MAPQ=60;MATEID=5076617_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_4753001_4778001_586C;SPAN=3284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:83 GQ:43.7 PL:[155.9, 0.0, 43.7] SR:54 DR:0 LR:-159.1 LO:159.1);ALT=G[chr12:4766913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	4764089	+	chr12	4766913	+	.	0	13	5076618_1	22.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=5076618_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_12_4753001_4778001_586C;SPAN=2824;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:13 DR:0 LR:-22.32 LO:28.48);ALT=G[chr12:4766913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
