chr13	61781604	+	chr13	61665128	+	.	9	0	8107684_1	15.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=8107684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:61665128(-)-13:61781604(+)__13_61642001_61667001D;SPAN=116476;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:0 DR:9 LR:-15.08 LO:19.6);ALT=]chr13:61781604]C;VARTYPE=BND:DUP-th;JOINTYPE=th
