chr11	128564172	+	chr11	128628008	+	.	17	19	5047122_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5047122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_128625001_128650001_323C;SPAN=63836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:37 GQ:3.2 PL:[85.7, 0.0, 3.2] SR:19 DR:17 LR:-90.16 LO:90.16);ALT=G[chr11:128628008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
