chr14	77787526	+	chr14	77791211	+	.	14	12	5809180_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5809180_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_14_77763001_77788001_332C;SPAN=3685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:39 GQ:38.9 PL:[38.9, 0.0, 55.4] SR:12 DR:14 LR:-38.95 LO:39.11);ALT=G[chr14:77791211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	77787526	+	chr14	77793180	+	CCCATCCTCTATTCCTATTTCCGAAGCTCCTGCTCATGGAGAGTTCGAATT	14	23	5809181_1	88.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CCCATCCTCTATTCCTATTTCCGAAGCTCCTGCTCATGGAGAGTTCGAATT;MAPQ=60;MATEID=5809181_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_77763001_77788001_332C;SPAN=5654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:39 GQ:5.9 PL:[88.4, 0.0, 5.9] SR:23 DR:14 LR:-92.71 LO:92.71);ALT=G[chr14:77793180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	77924613	+	chr14	77925958	+	.	0	28	5809605_1	62.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5809605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_77910001_77935001_145C;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:109 GQ:62.9 PL:[62.9, 0.0, 201.5] SR:28 DR:0 LR:-62.9 LO:66.96);ALT=G[chr14:77925958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	77926152	+	chr14	77928498	+	.	2	5	5809610_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GACAGGTA;MAPQ=60;MATEID=5809610_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_77910001_77935001_69C;SPAN=2346;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:90 GQ:4.5 PL:[0.0, 4.5, 227.7] SR:5 DR:2 LR:4.577 LO:10.53);ALT=A[chr14:77928498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	77978746	+	chr14	77984380	+	.	2	7	5809826_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5809826_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_77983501_78008501_120C;SPAN=5634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:7 DR:2 LR:-15.84 LO:18.23);ALT=C[chr14:77984380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	77984511	+	chr14	77987789	+	.	3	3	5809830_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5809830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_77983501_78008501_390C;SPAN=3278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:3 DR:3 LR:1.055 LO:10.95);ALT=C[chr14:77987789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78021864	+	chr14	78023384	+	.	13	5	5809961_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5809961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_78008001_78033001_265C;SPAN=1520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:87 GQ:29.3 PL:[29.3, 0.0, 181.1] SR:5 DR:13 LR:-29.25 LO:35.61);ALT=T[chr14:78023384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78063725	+	chr14	78082791	+	.	0	36	5810103_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5810103_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_78081501_78106501_39C;SPAN=19066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:53 GQ:22.1 PL:[104.6, 0.0, 22.1] SR:36 DR:0 LR:-107.3 LO:107.3);ALT=T[chr14:78082791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78174532	+	chr14	78182114	+	.	35	0	5810545_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5810545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:78174532(+)-14:78182114(-)__14_78179501_78204501D;SPAN=7582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:49 GQ:16.4 PL:[102.2, 0.0, 16.4] SR:0 DR:35 LR:-105.8 LO:105.8);ALT=T[chr14:78182114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78174553	+	chr14	78177181	+	CAGCTGAAAGAACACTTTGCACAGTTCGGCCATGTCAGAAGGTGCATTTTACCTTTT	11	26	5810531_1	62.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GT;INSERTION=CAGCTGAAAGAACACTTTGCACAGTTCGGCCATGTCAGAAGGTGCATTTTACCTTTT;MAPQ=60;MATEID=5810531_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_78155001_78180001_144C;SECONDARY;SPAN=2628;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:98 GQ:62.6 PL:[62.6, 0.0, 174.8] SR:26 DR:11 LR:-62.58 LO:65.54);ALT=T[chr14:78177181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78174553	+	chr14	78183836	+	CAGCTGAAAGAACACTTTGCACAGTTCGGCCATGTCAGAAGGTGCATTTTACCTTTTGACAAGGAGACTGGCTTTCACAGAGGTTTGGGTTGGGTTCAGTTTTCTTCAGAAGAAGGACTTCGGAATGCACTACAACAGGAAAATCATATTATAGATGGAGTA	4	78	5810547_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AAGGT;INSERTION=CAGCTGAAAGAACACTTTGCACAGTTCGGCCATGTCAGAAGGTGCATTTTACCTTTTGACAAGGAGACTGGCTTTCACAGAGGTTTGGGTTGGGTTCAGTTTTCTTCAGAAGAAGGACTTCGGAATGCACTACAACAGGAAAATCATATTATAGATGGAGTA;MAPQ=60;MATEID=5810547_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_14_78179501_78204501_101C;SPAN=9283;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:43 GQ:21 PL:[231.0, 21.0, 0.0] SR:78 DR:4 LR:-231.1 LO:231.1);ALT=T[chr14:78183836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78177240	+	chr14	78183836	+	ACAAGGAGACTGGCTTTCACAGAGGTTTGGGTTGGGTTCAGTTTTCTTCAGAAGAAGGACTTCGGAATGCACTACAACAGGAAAATCATATTATAGATGGAGTA	3	128	5810534_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AAGGT;INSERTION=ACAAGGAGACTGGCTTTCACAGAGGTTTGGGTTGGGTTCAGTTTTCTTCAGAAGAAGGACTTCGGAATGCACTACAACAGGAAAATCATATTATAGATGGAGTA;MAPQ=60;MATEID=5810534_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_78155001_78180001_106C;SPAN=6596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:60 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:128 DR:3 LR:-382.9 LO:382.9);ALT=G[chr14:78183836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78182224	+	chr14	78183836	+	.	0	43	5810555_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AAGGT;MAPQ=60;MATEID=5810555_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_14_78179501_78204501_101C;SPAN=1612;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:93 GQ:99 PL:[116.9, 0.0, 107.0] SR:43 DR:0 LR:-116.8 LO:116.8);ALT=T[chr14:78183836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78205406	+	chr14	78217660	+	.	2	4	5810630_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5810630_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_78204001_78229001_105C;SPAN=12254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:98 GQ:6.6 PL:[0.0, 6.6, 250.8] SR:4 DR:2 LR:6.745 LO:10.3);ALT=T[chr14:78217660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78217825	+	chr14	78221309	+	.	0	25	5810660_1	62.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5810660_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_78204001_78229001_102C;SPAN=3484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:74 GQ:62.6 PL:[62.6, 0.0, 115.4] SR:25 DR:0 LR:-62.48 LO:63.39);ALT=T[chr14:78221309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	78221456	+	chr14	78227456	+	.	14	0	5810672_1	15.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5810672_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:78221456(+)-14:78227456(-)__14_78204001_78229001D;SPAN=6000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:115 GQ:15.2 PL:[15.2, 0.0, 262.7] SR:0 DR:14 LR:-15.06 LO:28.42);ALT=G[chr14:78227456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
