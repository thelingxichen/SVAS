chr14	37769601	+	chr16	61079337	-	.	37	0	9356419_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=9356419_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:37769601(+)-16:61079337(+)__16_61078501_61103501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:37 DP:59 GQ:36.8 PL:[106.1, 0.0, 36.8] SR:0 DR:37 LR:-108.0 LO:108.0);ALT=T]chr16:61079337];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr16	60081112	+	chr16	60098562	+	.	123	115	9351739_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;MAPQ=29;MATEID=9351739_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_60098501_60123501_58C;SPAN=17450;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:185 DP:25 GQ:49.9 PL:[547.9, 49.9, 0.0] SR:115 DR:123 LR:-547.9 LO:547.9);ALT=G[chr16:60098562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
