chr2	130954939	+	chr2	130957404	+	.	54	43	1339805_1	99.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=CACACCTGTA;MAPQ=25;MATEID=1339805_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_130952501_130977501_272C;SPAN=2465;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:43 DR:54 LR:-237.7 LO:237.7);ALT=A[chr2:130957404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
