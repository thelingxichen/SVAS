chr2	220180587	+	chr2	208472402	+	CC	35	47	1697588_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CC;MAPQ=60;MATEID=1697588_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_220157001_220182001_265C;SPAN=11708185;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:71 DP:103 GQ:41.6 PL:[206.6, 0.0, 41.6] SR:47 DR:35 LR:-212.5 LO:212.5);ALT=]chr2:220180587]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	208474495	+	chr2	208476785	+	.	89	44	1650729_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAAACCTATTC;MAPQ=60;MATEID=1650729_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_208470501_208495501_355C;SPAN=2290;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:120 DP:31 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:44 DR:89 LR:-356.5 LO:356.5);ALT=C[chr2:208476785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209033781	+	chr17	19995674	-	.	58	0	1654719_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1654719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:209033781(+)-17:19995674(+)__2_209009501_209034501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:58 DP:61 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:58 LR:-178.2 LO:178.2);ALT=A]chr17:19995674];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	231930032	-	chr19	54800810	+	.	9	0	10373895_1	19.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=10373895_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231930032(-)-19:54800810(-)__19_54782001_54807001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=[chr19:54800810[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	231930154	+	chr19	54800680	-	.	17	0	10373896_1	46.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=10373896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231930154(+)-19:54800680(+)__19_54782001_54807001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:17 DP:37 GQ:42.8 PL:[46.1, 0.0, 42.8] SR:0 DR:17 LR:-46.1 LO:46.1);ALT=C]chr19:54800680];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	232705543	+	chr2	232703709	+	.	53	0	1751501_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=1751501_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232703709(-)-2:232705543(+)__2_232701001_232726001D;SPAN=1834;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:118 GQ:99 PL:[143.0, 0.0, 143.0] SR:0 DR:53 LR:-143.0 LO:143.0);ALT=]chr2:232705543]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	232713985	+	chr2	232712304	+	.	68	0	1751533_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=1751533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232712304(-)-2:232713985(+)__2_232701001_232726001D;SPAN=1681;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:106 GQ:60.5 PL:[195.8, 0.0, 60.5] SR:0 DR:68 LR:-199.6 LO:199.6);ALT=]chr2:232713985]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	232847537	+	chr2	232848626	-	.	9	0	1750836_1	18.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1750836_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232847537(+)-2:232848626(+)__2_232848001_232873001D;SPAN=1089;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=C]chr2:232848626];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	116368767	+	chr9	6360629	-	TAGCTACAAAATTAGCCAGGCATGGTGTCACATGCTTGT	6	59	4365811_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=TAGCTACAAAATTAGCCAGGCATGGTGTCACATGCTTGT;MAPQ=60;MATEID=4365811_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_6_116350501_116375501_5C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:59 DP:26 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:59 DR:6 LR:-174.9 LO:174.9);ALT=T]chr9:6360629];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	6798901	+	chr10	6248506	+	.	11	0	6072090_1	29.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6072090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:6798901(+)-10:6248506(-)__10_6247501_6272501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=A[chr10:6248506[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr19	53773169	+	chr10	6248540	+	.	10	0	6072098_1	27.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6072098_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:6248540(-)-19:53773169(+)__10_6247501_6272501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:20 GQ:20.9 PL:[27.5, 0.0, 20.9] SR:0 DR:10 LR:-27.64 LO:27.64);ALT=]chr19:53773169]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	6411580	+	chr10	6417630	+	.	76	37	6071734_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGCAAATCATTTTCCT;MAPQ=60;MATEID=6071734_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_10_6394501_6419501_61C;SPAN=6050;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:48 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:37 DR:76 LR:-287.2 LO:287.2);ALT=T[chr10:6417630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	106044581	+	chr19	49290023	+	.	14	37	10343319_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCCATAAAGAAATAGCACTTGA;MAPQ=60;MATEID=10343319_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_49269501_49294501_155C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:73 GQ:66.2 PL:[109.1, 0.0, 66.2] SR:37 DR:14 LR:-109.5 LO:109.5);ALT=A[chr19:49290023[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr19	54819659	+	chr14	97671207	+	.	4	37	10374132_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATATATATATATATATATATATATATAT;MAPQ=60;MATEID=10374132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54806501_54831501_305C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:26 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:37 DR:4 LR:-118.8 LO:118.8);ALT=]chr19:54819659]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	20492232	+	chr19	47922793	-	.	22	0	10335123_1	63.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=10335123_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:20492232(+)-19:47922793(+)__19_47922001_47947001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:35 GQ:20.3 PL:[63.2, 0.0, 20.3] SR:0 DR:22 LR:-64.24 LO:64.24);ALT=C]chr19:47922793];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr17	20616861	-	chr17	20617869	+	.	6	2	9562825_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCTCACTGCAACCTC;MAPQ=60;MATEID=9562825_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_20604501_20629501_251C;SPAN=1008;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:7 DP:154 GQ:18.4 PL:[0.0, 18.4, 409.3] SR:2 DR:6 LR:18.62 LO:11.1);ALT=[chr17:20617869[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	21345304	+	chr17	21443258	+	.	43	33	9566675_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=9566675_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_21437501_21462501_106C;SPAN=97954;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:38 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:33 DR:43 LR:-184.8 LO:184.8);ALT=T[chr17:21443258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	21556719	+	chr17	21558069	+	.	0	135	9568003_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CA;MAPQ=27;MATEID=9568003_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_17_21535501_21560501_370C;SPAN=1350;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:135 DP:176 GQ:28.3 PL:[398.0, 0.0, 28.3] SR:135 DR:0 LR:-416.8 LO:416.8);ALT=A[chr17:21558069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48583806	-	chr19	48586142	+	.	9	0	10338522_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=10338522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48583806(-)-19:48586142(-)__19_48583501_48608501D;SPAN=2336;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:173 GQ:16.9 PL:[0.0, 16.9, 452.2] SR:0 DR:9 LR:17.16 LO:14.8);ALT=[chr19:48586142[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	49670789	+	chr19	49669581	+	.	23	0	10345572_1	39.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=10345572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49669581(-)-19:49670789(+)__19_49661501_49686501D;SPAN=1208;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:135 GQ:39.5 PL:[39.5, 0.0, 287.0] SR:0 DR:23 LR:-39.35 LO:50.34);ALT=]chr19:49670789]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	50272479	+	chr19	52935944	-	.	9	58	10363339_1	99.0	.	DISC_MAPQ=19;EVDNC=ASDIS;HOMSEQ=CTGGAGTGCAATG;MAPQ=54;MATEID=10363339_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52920001_52945001_198C;SPAN=2663465;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:63 DP:59 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:58 DR:9 LR:-184.8 LO:184.8);ALT=G]chr19:52935944];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	52888816	+	chr19	52891387	+	A	64	57	10363034_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=10363034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52871001_52896001_380C;SPAN=2571;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:95 DP:101 GQ:27 PL:[297.0, 27.0, 0.0] SR:57 DR:64 LR:-297.1 LO:297.1);ALT=A[chr19:52891387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53041673	+	chr19	53225285	-	.	6	9	10364021_1	24.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=TCATTAGCCAAGATTGTGCCATTGCACTCCAGCCTGGGCAACA;MAPQ=60;MATEID=10364021_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_19_53018001_53043001_300C;SPAN=183612;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:79 GQ:24.8 PL:[24.8, 0.0, 166.7] SR:9 DR:6 LR:-24.81 LO:30.91);ALT=A]chr19:53225285];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	53096022	+	chr19	53097609	+	.	64	38	10363602_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTAATTTTGTATTTTT;MAPQ=60;MATEID=10363602_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_53091501_53116501_159C;SPAN=1587;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:78 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:38 DR:64 LR:-267.4 LO:267.4);ALT=T[chr19:53097609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53135358	+	chr19	54339143	+	.	15	0	10371815_1	35.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=10371815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53135358(+)-19:54339143(-)__19_54316501_54341501D;SPAN=1203785;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:51 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.7 LO:36.92);ALT=G[chr19:54339143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53193323	+	chr19	53869417	-	.	34	0	10368348_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=10368348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53193323(+)-19:53869417(+)__19_53851001_53876001D;SPAN=676094;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:34 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:34 LR:-102.3 LO:102.3);ALT=G]chr19:53869417];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	53356862	+	chr19	53320000	+	TCCCGAGTAGCTGGGATTACAGGCGTGCACCACCACGCCCAGCTAATTTTGTATTTTTAGTAGAGACGGGGTTTCTCCATGTTGGTCAGACTGGTCTCAAACTCCAGACCTCACGTGATTTGCCCACCTTGGCCTCCTAAAGTGCTAGGATTACAGGCATCAGTCACTGTGCCCGGCCTATTCCTTCATTATTTTAAGAATAGGAAATCAACGTAAATCATAGCAGGAGATTCATTCAACCATTCTTAGCACATTAAGCTGATGGAGACAGGGTGTTACTGTGGAGAGGCTTGTGAAACAGGCTTTTGGTAAAAATGGTTACAATTTTTCTCAAATATGGGAGCAGTACTTCTTTTTTATCCTAGAGGAGAAAGCCGTATTCTCATTCCACC	41	59	10366159_1	99.0	.	DISC_MAPQ=20;EVDNC=TSI_L;HOMSEQ=AAG;INSERTION=TCCCGAGTAGCTGGGATTACAGGCGTGCACCACCACGCCCAGCTAATTTTGTATTTTTAGTAGAGACGGGGTTTCTCCATGTTGGTCAGACTGGTCTCAAACTCCAGACCTCACGTGATTTGCCCACCTTGGCCTCCTAAAGTGCTAGGATTACAGGCATCAGTCACTGTGCCCGGCCTATTCCTTCATTATTTTAAGAATAGGAAATCAACGTAAATCATAGCAGGAGATTCATTCAACCATTCTTAGCACATTAAGCTGATGGAGACAGGGTGTTACTGTGGAGAGGCTTGTGAAACAGGCTTTTGGTAAAAATGGTTACAATTTTTCTCAAATATGGGAGCAGTACTTCTTTTTTATCCTAGAGGAGAAAGCCGTATTCTCATTCCACC;MAPQ=60;MATEID=10366159_2;MATENM=0;NM=4;NUMPARTS=3;SCTG=c_19_53336501_53361501_240C;SPAN=36862;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:71 GQ:21 PL:[231.0, 21.0, 0.0] SR:59 DR:41 LR:-231.1 LO:231.1);ALT=]chr19:53356862]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	53422214	+	chr19	53424208	+	.	72	15	10365958_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAATCT;MAPQ=60;MATEID=10365958_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_53410001_53435001_366C;SPAN=1994;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:83 DP:144 GQ:99 PL:[235.1, 0.0, 113.0] SR:15 DR:72 LR:-237.2 LO:237.2);ALT=T[chr19:53424208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54540315	+	chr19	53435123	+	.	27	0	10372611_1	79.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=10372611_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53435123(-)-19:54540315(+)__19_54537001_54562001D;SPAN=1105192;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:27 DP:22 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:0 DR:27 LR:-79.22 LO:79.22);ALT=]chr19:54540315]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	53435459	+	chr19	54540595	+	.	25	0	10372612_1	71.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=10372612_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53435459(+)-19:54540595(-)__19_54537001_54562001D;SPAN=1105136;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:25 DP:41 GQ:25.4 PL:[71.6, 0.0, 25.4] SR:0 DR:25 LR:-72.45 LO:72.45);ALT=G[chr19:54540595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53689177	+	chr19	53691952	+	.	48	28	10367996_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GGGTTTTT;MAPQ=60;MATEID=10367996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_53679501_53704501_442C;SPAN=2775;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:134 GQ:99 PL:[175.1, 0.0, 148.7] SR:28 DR:48 LR:-175.1 LO:175.1);ALT=T[chr19:53691952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53788567	+	chr19	53801887	-	.	10	0	10367447_1	4.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=10367447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53788567(+)-19:53801887(+)__19_53777501_53802501D;SPAN=13320;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:107 GQ:4.1 PL:[4.1, 0.0, 254.9] SR:0 DR:10 LR:-4.021 LO:19.08);ALT=A]chr19:53801887];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	54384950	+	chr19	54383882	+	.	10	0	10371137_1	0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=10371137_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54383882(-)-19:54384950(+)__19_54365501_54390501D;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:222 GQ:26.8 PL:[0.0, 26.8, 590.8] SR:0 DR:10 LR:27.14 LO:15.81);ALT=]chr19:54384950]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54428571	+	chr19	54425402	+	.	153	0	10372330_1	99.0	.	DISC_MAPQ=19;EVDNC=ASDIS;HOMSEQ=CCCCAGGTCTGGTCATTGGTGGAGTTGTCCCAGGTCTGGTCATTGGTGGAGTTG;MAPQ=0;MATEID=10372330_2;MATENM=0;NM=3;NUMPARTS=2;REPSEQ=CCC;SCTG=c_19_54414501_54439501_436C;SECONDARY;SPAN=3169;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:153 DP:182 GQ:16 PL:[472.0, 16.0, 0.0] SR:0 DR:153 LR:-487.7 LO:487.7);ALT=]chr19:54428571]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54800910	+	chr19	54807620	+	.	23	0	10374136_1	65.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=10374136_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54800910(+)-19:54807620(-)__19_54806501_54831501D;SPAN=6710;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:23 DP:39 GQ:29 PL:[65.3, 0.0, 29.0] SR:0 DR:23 LR:-66.1 LO:66.1);ALT=G[chr19:54807620[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
