chr6	146865258	+	chr6	146870599	+	.	9	13	3063619_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3063619_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_146853001_146878001_106C;SPAN=5341;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:87 GQ:39.2 PL:[39.2, 0.0, 171.2] SR:13 DR:9 LR:-39.15 LO:43.89);ALT=G[chr6:146870599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
