chr11	54885354	+	chr11	54892206	+	.	51	15	4863067_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GGCCTATGGTGAAAAAGGAAATATCTTC;MAPQ=60;MATEID=4863067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_54880001_54905001_87C;SPAN=6852;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:22 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:15 DR:51 LR:-181.5 LO:181.5);ALT=C[chr11:54892206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	55016471	+	chr11	55014914	+	.	70	25	4863538_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=TTTGCAGATTCTACAAAGAGA;MAPQ=60;MATEID=4863538_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_55002501_55027501_292C;SPAN=1557;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:97 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:25 DR:70 LR:-287.2 LO:287.2);ALT=]chr11:55016471]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	55196437	+	chr11	55084689	+	.	11	0	4863395_1	27.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=4863395_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:55084689(-)-11:55196437(+)__11_55076001_55101001D;SPAN=111748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:33 GQ:27.5 PL:[27.5, 0.0, 50.6] SR:0 DR:11 LR:-27.37 LO:27.81);ALT=]chr11:55196437]G;VARTYPE=BND:DUP-th;JOINTYPE=th
