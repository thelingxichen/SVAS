chr4	21161002	+	chr4	21167098	+	.	13	15	1918696_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGAAAATTATACTAAA;MAPQ=60;MATEID=1918696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_21143501_21168501_67C;SPAN=6096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:28 GQ:5.6 PL:[61.7, 0.0, 5.6] SR:15 DR:13 LR:-64.39 LO:64.39);ALT=A[chr4:21167098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
