chr1	196601824	-	chr1	196603253	+	.	8	0	477820_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=477820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:196601824(-)-1:196603253(-)__1_196588001_196613001D;SPAN=1429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:0 DR:8 LR:2.581 LO:14.46);ALT=[chr1:196603253[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	197500520	+	chr1	197503272	+	.	122	85	480839_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AACAAATCTTTT;MAPQ=60;MATEID=480839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_197494501_197519501_334C;SPAN=2752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:157 DP:61 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:85 DR:122 LR:-465.4 LO:465.4);ALT=T[chr1:197503272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	197742108	+	chr1	197744337	+	.	9	0	481041_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=481041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:197742108(+)-1:197744337(-)__1_197739501_197764501D;SPAN=2229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:0 DR:9 LR:-4.242 LO:17.27);ALT=C[chr1:197744337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198608472	+	chr1	198665840	+	GCAAAGCCCAACACCTTCCCCCACT	33	30	483817_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GCAAAGCCCAACACCTTCCCCCACT;MAPQ=60;MATEID=483817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198646001_198671001_263C;SPAN=57368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:67 GQ:31.4 PL:[130.4, 0.0, 31.4] SR:30 DR:33 LR:-133.7 LO:133.7);ALT=G[chr1:198665840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198608472	+	chr1	198661473	+	.	11	7	483816_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=483816_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198646001_198671001_266C;SPAN=53001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:7 DR:11 LR:-21.68 LO:25.03);ALT=G[chr1:198661473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198608472	+	chr1	198668692	+	GCAAAGCCCAACACCTTCCCCCACT	0	14	483818_1	26.0	.	EVDNC=ASSMB;INSERTION=GCAAAGCCCAACACCTTCCCCCACT;MAPQ=60;MATEID=483818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198646001_198671001_38C;SPAN=60220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:14 DR:0 LR:-26.17 LO:31.35);ALT=G[chr1:198668692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198666040	+	chr1	198668691	+	.	0	10	483882_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=483882_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198646001_198671001_359C;SPAN=2651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:129 GQ:1.8 PL:[0.0, 1.8, 316.8] SR:10 DR:0 LR:1.939 LO:18.23);ALT=T[chr1:198668691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198668833	+	chr1	198671513	+	.	0	13	483900_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=483900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198670501_198695501_168C;SPAN=2680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:97 GQ:16.7 PL:[16.7, 0.0, 218.0] SR:13 DR:0 LR:-16.63 LO:26.97);ALT=G[chr1:198671513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198676082	+	chr1	198677259	+	.	0	6	483918_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=483918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198670501_198695501_311C;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:102 GQ:7.5 PL:[0.0, 7.5, 260.7] SR:6 DR:0 LR:7.828 LO:10.2);ALT=G[chr1:198677259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198701686	+	chr1	198704255	+	GTTTCAAAGAACCCAGGAAATACATTGCTGCACAAGGTCCCAGGGATGAAACTGTTGATGATTTCTGGAGGATGATTTGGGAACAGAAAGCCACAGTTATTGTCATGGTCACTCGATGTGAAGAAGGAAACAG	2	15	483982_1	23.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GTTTCAAAGAACCCAGGAAATACATTGCTGCACAAGGTCCCAGGGATGAAACTGTTGATGATTTCTGGAGGATGATTTGGGAACAGAAAGCCACAGTTATTGTCATGGTCACTCGATGTGAAGAAGGAAACAG;MAPQ=60;MATEID=483982_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_198695001_198720001_123C;SPAN=2569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:96 GQ:23.6 PL:[23.6, 0.0, 208.4] SR:15 DR:2 LR:-23.51 LO:32.21);ALT=G[chr1:198704255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198704381	+	chr1	198710998	+	.	5	5	483990_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=483990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198695001_198720001_310C;SPAN=6617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:5 DR:5 LR:-5.326 LO:17.45);ALT=T[chr1:198710998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198711497	+	chr1	198713181	+	.	0	11	484007_1	3.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=484007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198695001_198720001_89C;SPAN=1684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:122 GQ:3.5 PL:[3.5, 0.0, 290.6] SR:11 DR:0 LR:-3.258 LO:20.81);ALT=G[chr1:198713181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198721902	+	chr1	198723396	+	.	6	6	484052_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=484052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198719501_198744501_39C;SPAN=1494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:89 GQ:12.2 PL:[12.2, 0.0, 203.6] SR:6 DR:6 LR:-12.2 LO:22.41);ALT=G[chr1:198723396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198723534	+	chr1	198725035	+	.	10	6	484055_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=484055_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198719501_198744501_15C;SPAN=1501;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:109 GQ:16.7 PL:[16.7, 0.0, 247.7] SR:6 DR:10 LR:-16.68 LO:28.77);ALT=G[chr1:198725035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198869698	+	chr1	198906355	+	.	0	16	484493_1	39.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=484493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198891001_198916001_343C;SPAN=36657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:16 DR:0 LR:-39.54 LO:40.27);ALT=T[chr1:198906355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	198875870	+	chr1	198906355	+	.	0	15	484495_1	36.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=484495_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_198891001_198916001_16C;SPAN=30485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:49 GQ:36.2 PL:[36.2, 0.0, 82.4] SR:15 DR:0 LR:-36.24 LO:37.24);ALT=T[chr1:198906355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	199589210	-	chr1	199590390	+	.	5	2	486416_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=486416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_199577001_199602001_131C;SPAN=1180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:90 GQ:4.5 PL:[0.0, 4.5, 227.7] SR:2 DR:5 LR:4.577 LO:10.53);ALT=[chr1:199590390[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	200067552	-	chr2	23698253	+	.	17	41	716886_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=716886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_23691501_23716501_356C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:43 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:41 DR:17 LR:-148.5 LO:148.5);ALT=[chr2:23698253[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	200067673	+	chr2	23698254	-	.	23	44	716888_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=716888_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_23691501_23716501_54C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:42 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:44 DR:23 LR:-181.5 LO:181.5);ALT=C]chr2:23698254];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	24291329	+	chr2	24296945	+	.	5	122	718834_1	99.0	.	DISC_MAPQ=35;EVDNC=TSI_L;HOMSEQ=C;MAPQ=15;MATEID=718834_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CCCC;SCTG=c_2_24279501_24304501_172C;SPAN=5616;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:127 DP:113 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:122 DR:5 LR:-376.3 LO:376.3);ALT=C[chr2:24296945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24291356	+	chr2	24299069	+	.	53	0	718835_1	99.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=718835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:24291356(+)-2:24299069(-)__2_24279501_24304501D;SPAN=7713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:83 GQ:47 PL:[152.6, 0.0, 47.0] SR:0 DR:53 LR:-155.4 LO:155.4);ALT=A[chr2:24299069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24297064	+	chr2	24299070	+	.	123	44	718855_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=CACTCTGATTTGACGAATAGGTCCATATTTCCCAAATATATCATACATTTCTTCAGCTGTGATTTTGTATGGCAAATTTCTTATATACAATATCCGATTTACTTCAGGTGGAAGTCGAATGTTCGCCCTCTTGGCCGCTTGCA;MAPQ=60;MATEID=718855_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_2_24279501_24304501_172C;SPAN=2006;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:157 DP:79 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:44 DR:123 LR:-465.4 LO:465.4);ALT=T[chr2:24299070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24303825	+	chr2	24318010	+	.	2	6	719021_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=719021_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_24304001_24329001_381C;SPAN=14185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:6 DR:2 LR:-18.01 LO:19.15);ALT=G[chr2:24318010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24306027	+	chr2	24307059	+	.	0	11	719031_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CTGCA;MAPQ=60;MATEID=719031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_24304001_24329001_194C;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:106 GQ:7.7 PL:[7.7, 0.0, 248.6] SR:11 DR:0 LR:-7.593 LO:21.52);ALT=A[chr2:24307059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24538094	+	chr2	24583173	+	ATTCATAGCTGTGGGAAACTGAGCCATCATGGTCCTGAGTTTTCCTTGCTAGCTCTCAGCCAT	0	22	720021_1	65.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATTCATAGCTGTGGGAAACTGAGCCATCATGGTCCTGAGTTTTCCTTGCTAGCTCTCAGCCAT;MAPQ=60;MATEID=720021_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_2_24573501_24598501_100C;SPAN=45079;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:28 GQ:2.3 PL:[65.0, 0.0, 2.3] SR:22 DR:0 LR:-68.45 LO:68.45);ALT=C[chr2:24583173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	24550987	+	chr2	24583173	+	.	15	15	720023_1	69.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=720023_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_2_24573501_24598501_100C;SPAN=32186;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:28 GQ:0.9 PL:[69.3, 0.9, 0.0] SR:15 DR:15 LR:-72.68 LO:72.68);ALT=G[chr2:24583173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
