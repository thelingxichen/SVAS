chr1	120578314	-	chr1	145242756	+	.	4	2	281121_1	0	.	DISC_MAPQ=5;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=281121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_120564501_120589501_131C;SPAN=24664442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:112 GQ:13.5 PL:[0.0, 13.5, 297.0] SR:2 DR:4 LR:13.84 LO:7.886);ALT=[chr1:145242756[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	144896297	+	chr1	144901047	+	GTAACAGG	37	42	296991_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;INSERTION=GTAACAGG;MAPQ=60;MATEID=296991_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_1_144893001_144918001_148C;SPAN=4750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:112 GQ:75.5 PL:[194.3, 0.0, 75.5] SR:42 DR:37 LR:-196.8 LO:196.8);ALT=G[chr1:144901047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	144896297	+	chr1	144906810	+	GTAACAGGATTTATCCTGCTATCAATTTACTCTTGCTGGAGGTTGACAGAAGTAGGAGTGATTATTAACATAAACTGTAATCACTATGAGCCATTAGAAACGAAGAATCACCCAGAGCTGAATCTTACTAGCGATTCAGAAG	17	89	296992_1	99.0	.	DISC_MAPQ=47;EVDNC=TSI_G;INSERTION=GTAACAGGATTTATCCTGCTATCAATTTACTCTTGCTGGAGGTTGACAGAAGTAGGAGTGATTATTAACATAAACTGTAATCACTATGAGCCATTAGAAACGAAGAATCACCCAGAGCTGAATCTTACTAGCGATTCAGAAG;MAPQ=60;MATEID=296992_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_144893001_144918001_148C;SPAN=10513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:96 DP:122 GQ:10.1 PL:[284.0, 0.0, 10.1] SR:89 DR:17 LR:-298.9 LO:298.9);ALT=G[chr1:144906810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	144901180	+	chr1	144906810	+	GTAACAGG	41	61	297002_1	99.0	.	DISC_MAPQ=32;EVDNC=TSI_L;INSERTION=GTAACAGG;MAPQ=60;MATEID=297002_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_1_144893001_144918001_148C;SPAN=5630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:124 GQ:45.8 PL:[253.7, 0.0, 45.8] SR:61 DR:41 LR:-261.6 LO:261.6);ALT=G[chr1:144906810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145096621	+	chr1	145103905	+	.	9	9	298779_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=298779_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_145089001_145114001_363C;SPAN=7284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:170 GQ:3.4 PL:[3.4, 0.0, 409.4] SR:9 DR:9 LR:-3.458 LO:28.23);ALT=G[chr1:145103905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145104017	+	chr1	145109524	+	.	0	7	298840_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=298840_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_1_145089001_145114001_752C;SPAN=5507;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:257 GQ:46.3 PL:[0.0, 46.3, 716.2] SR:7 DR:0 LR:46.52 LO:9.527);ALT=A[chr1:145109524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145459827	+	chr1	145470319	+	.	25	0	301603_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=301603_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:145459827(+)-1:145470319(-)__1_145456501_145481501D;SPAN=10492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:123 GQ:49.4 PL:[49.4, 0.0, 247.4] SR:0 DR:25 LR:-49.2 LO:56.86);ALT=A[chr1:145470319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145460265	+	chr1	145470320	+	.	53	4	301604_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=301604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_145456501_145481501_272C;SPAN=10055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:118 GQ:99 PL:[149.6, 0.0, 136.4] SR:4 DR:53 LR:-149.6 LO:149.6);ALT=T[chr1:145470320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145516470	+	chr1	145518070	+	.	10	0	302545_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=302545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:145516470(+)-1:145518070(-)__1_145505501_145530501D;SPAN=1600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:109 GQ:3.5 PL:[3.5, 0.0, 260.9] SR:0 DR:10 LR:-3.479 LO:19.0);ALT=A[chr1:145518070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145592771	+	chr1	145594037	+	.	0	7	303089_1	0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=303089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_145579001_145604001_157C;SPAN=1266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:114 GQ:7.5 PL:[0.0, 7.5, 290.4] SR:7 DR:0 LR:7.778 LO:12.03);ALT=C[chr1:145594037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	145609388	+	chr1	145610817	+	.	9	0	303727_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=303727_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:145609388(+)-1:145610817(-)__1_145603501_145628501D;SPAN=1429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:96 GQ:3.8 PL:[3.8, 0.0, 228.2] SR:0 DR:9 LR:-3.7 LO:17.19);ALT=A[chr1:145610817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
