chr12	100288344	+	chr12	100291788	+	TA	14	11	5308096_1	53.0	.	DISC_MAPQ=50;EVDNC=ASDIS;INSERTION=TA;MAPQ=60;MATEID=5308096_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_100278501_100303501_302C;SPAN=3444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:59 GQ:53.3 PL:[53.3, 0.0, 89.6] SR:11 DR:14 LR:-53.34 LO:53.85);ALT=A[chr12:100291788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	100594689	+	chr12	100598717	+	.	14	0	5308955_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5308955_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:100594689(+)-12:100598717(-)__12_100597001_100622001D;SPAN=4028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:43 GQ:34.7 PL:[34.7, 0.0, 67.7] SR:0 DR:14 LR:-34.56 LO:35.22);ALT=A[chr12:100598717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
