chr14	99929915	+	chr14	99932040	+	.	0	8	5863755_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5863755_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_99911001_99936001_81C;SPAN=2125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:8 DR:0 LR:-1.483 LO:15.0);ALT=T[chr14:99932040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	99932177	+	chr14	99947080	+	.	11	0	5863764_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5863764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:99932177(+)-14:99947080(-)__14_99911001_99936001D;SPAN=14903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:33 GQ:27.5 PL:[27.5, 0.0, 50.6] SR:0 DR:11 LR:-27.37 LO:27.81);ALT=A[chr14:99947080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	99947863	+	chr14	99958987	+	.	10	0	5863605_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5863605_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:99947863(+)-14:99958987(-)__14_99935501_99960501D;SPAN=11124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:78 GQ:11.9 PL:[11.9, 0.0, 176.9] SR:0 DR:10 LR:-11.88 LO:20.54);ALT=T[chr14:99958987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100531848	+	chr14	100551022	+	.	32	4	5865388_1	94.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5865388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_100523501_100548501_121C;SPAN=19174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:42 GQ:5.3 PL:[94.4, 0.0, 5.3] SR:4 DR:32 LR:-98.59 LO:98.59);ALT=G[chr14:100551022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100531859	+	chr14	100563814	+	.	12	0	5865389_1	28.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5865389_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:100531859(+)-14:100563814(-)__14_100523501_100548501D;SPAN=31955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:42 GQ:28.4 PL:[28.4, 0.0, 71.3] SR:0 DR:12 LR:-28.23 LO:29.36);ALT=G[chr14:100563814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100551194	+	chr14	100563815	+	.	2	16	5865310_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=5865310_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_100548001_100573001_308C;SPAN=12621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:87 GQ:35.9 PL:[35.9, 0.0, 174.5] SR:16 DR:2 LR:-35.85 LO:41.09);ALT=T[chr14:100563815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100706260	+	chr14	100728637	+	.	2	7	5865757_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=5865757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_100719501_100744501_3C;SPAN=22377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:7 DR:2 LR:-16.11 LO:18.33);ALT=G[chr14:100728637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100828260	+	chr14	100835423	+	.	4	5	5866596_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5866596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_100817501_100842501_71C;SPAN=7163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:5 DR:4 LR:1.005 LO:12.81);ALT=T[chr14:100835423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	100828287	+	chr14	100842595	+	.	9	0	5866641_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5866641_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:100828287(+)-14:100842595(-)__14_100842001_100867001D;SPAN=14308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=A[chr14:100842595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
