chr3	83853128	+	chr3	83855350	+	.	70	43	1515025_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATATGGCCTTTT;MAPQ=60;MATEID=1515025_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_83839001_83864001_309C;SPAN=2222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:34 GQ:24 PL:[264.0, 24.0, 0.0] SR:43 DR:70 LR:-264.1 LO:264.1);ALT=T[chr3:83855350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	84104942	+	chr3	84107385	+	.	109	76	1515550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=1515550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_84084001_84109001_235C;SPAN=2443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:34 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:76 DR:109 LR:-429.1 LO:429.1);ALT=C[chr3:84107385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	84699513	+	chr3	84702893	+	.	16	0	1517389_1	28.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=1517389_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:84699513(+)-3:84702893(-)__3_84696501_84721501D;SPAN=3380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:91 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:0 DR:16 LR:-28.16 LO:35.26);ALT=T[chr3:84702893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
