chr4	19354467	-	chr5	13827595	+	CGTGGCTGTACCCTGAAAAGCCACAGGCGTGGAGCTGCCCAAGGCTTTAGGAGCCCACCTCTTGCATCAGCAGGTCTGGATGTGAGACATGGAGTCAAAGCAGATCATTTTGGAAATTTAAGGTTTAATTACTGCCTTATTGAATTTTGGACTTGCATGAGGCCTGTAGCCTCTTTGTTTTGGCCAATTTCTCCCATTTGGAACAGGTATATTTACC	12	145	3225448_1	99.0	.	DISC_MAPQ=24;EVDNC=TSI_G;HOMSEQ=CAATGCCTGTACCCCCATTGTATCTAGGGAGTAACTAACTT;INSERTION=CGTGGCTGTACCCTGAAAAGCCACAGGCGTGGAGCTGCCCAAGGCTTTAGGAGCCCACCTCTTGCATCAGCAGGTCTGGATGTGAGACATGGAGTCAAAGCAGATCATTTTGGAAATTTAAGGTTTAATTACTGCCTTATTGAATTTTGGACTTGCATGAGGCCTGTAGCCTCTTTGTTTTGGCCAATTTCTCCCATTTGGAACAGGTATATTTACC;MAPQ=60;MATEID=3225448_2;MATENM=0;NM=2;NUMPARTS=6;SCTG=c_5_13818001_13843001_787C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:147 DP:77 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:145 DR:12 LR:-435.7 LO:435.7);ALT=[chr5:13827595[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	13416607	+	chr5	13422854	+	.	161	93	3221588_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATCACGTCAACC;MAPQ=60;MATEID=3221588_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_13401501_13426501_468C;SPAN=6247;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:204 DP:115 GQ:55 PL:[604.0, 55.0, 0.0] SR:93 DR:161 LR:-604.0 LO:604.0);ALT=C[chr5:13422854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
