chr4	183836260	+	chr4	183838440	+	.	22	0	2371850_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2371850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:183836260(+)-4:183838440(-)__4_183823501_183848501D;SPAN=2180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:81 GQ:50.9 PL:[50.9, 0.0, 143.3] SR:0 DR:22 LR:-50.68 LO:53.24);ALT=G[chr4:183838440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	183836729	+	chr4	183838464	+	.	19	2	2371853_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2371853_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_183823501_183848501_244C;SPAN=1735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:78 GQ:44.9 PL:[44.9, 0.0, 143.9] SR:2 DR:19 LR:-44.89 LO:47.81);ALT=C[chr4:183838464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	184630709	+	chr4	184631729	-	.	9	0	2374752_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2374752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:184630709(+)-4:184631729(+)__4_184607501_184632501D;SPAN=1020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:110 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.0927 LO:16.63);ALT=A]chr4:184631729];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	185178528	+	chr4	185181485	+	.	0	29	2376868_1	74.0	.	EVDNC=ASSMB;HOMSEQ=GGAA;MAPQ=36;MATEID=2376868_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_4_185171001_185196001_110C;SPAN=2957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:78 GQ:74.6 PL:[74.6, 0.0, 114.2] SR:29 DR:0 LR:-74.6 LO:75.06);ALT=A[chr4:185181485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	185350272	+	chr4	185395622	+	.	11	0	2377776_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2377776_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:185350272(+)-4:185395622(-)__4_185391501_185416501D;SPAN=45350;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:43 GQ:24.8 PL:[24.8, 0.0, 77.6] SR:0 DR:11 LR:-24.66 LO:26.28);ALT=G[chr4:185395622[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	185570998	+	chr4	185573175	+	.	8	0	2378541_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2378541_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:185570998(+)-4:185573175(-)__4_185563001_185588001D;SPAN=2177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=C[chr4:185573175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	185612867	+	chr4	185615674	+	.	4	3	2378425_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2378425_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_185612001_185637001_219C;SPAN=2807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:107 GQ:9 PL:[0.0, 9.0, 277.2] SR:3 DR:4 LR:9.183 LO:10.07);ALT=G[chr4:185615674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	185646217	+	chr4	185650072	+	.	0	9	2378731_1	3.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2378731_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_185636501_185661501_7C;SPAN=3855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:9 DR:0 LR:-3.158 LO:17.1);ALT=C[chr4:185650072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	185650236	+	chr4	185655169	+	.	13	0	2378753_1	17.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=2378753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:185650236(+)-4:185655169(-)__4_185636501_185661501D;SPAN=4933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:95 GQ:17.3 PL:[17.3, 0.0, 212.0] SR:0 DR:13 LR:-17.18 LO:27.1);ALT=C[chr4:185655169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	186112367	+	chr4	186124939	+	.	16	2	2380468_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2380468_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_186102001_186127001_159C;SPAN=12572;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:109 GQ:26.6 PL:[26.6, 0.0, 237.8] SR:2 DR:16 LR:-26.59 LO:36.49);ALT=C[chr4:186124939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	186339925	+	chr4	186347016	+	ATTAGGAGTAGCTAGCTGAAAAGCCAAATCAAGGCCTCCTCTTATTCTGAAGAGTATATCCATACTTTCTGAAA	10	8	2381525_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TCACC;INSERTION=ATTAGGAGTAGCTAGCTGAAAAGCCAAATCAAGGCCTCCTCTTATTCTGAAGAGTATATCCATACTTTCTGAAA;MAPQ=60;MATEID=2381525_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_186347001_186372001_455C;SPAN=7091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:58 GQ:37.1 PL:[37.1, 0.0, 103.1] SR:8 DR:10 LR:-37.1 LO:38.85);ALT=C[chr4:186347016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	186339925	+	chr4	186343639	+	.	2	6	2381151_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2381151_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_4_186322501_186347501_333C;SPAN=3714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:6 DR:2 LR:0.4135 LO:14.74);ALT=C[chr4:186343639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	186343718	+	chr4	186347016	+	.	4	4	2381165_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TCACC;MAPQ=60;MATEID=2381165_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_4_186322501_186347501_333C;SPAN=3298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:105 GQ:11.7 PL:[0.0, 11.7, 277.2] SR:4 DR:4 LR:11.94 LO:8.028);ALT=C[chr4:186347016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	186441692	+	chr4	186444073	+	.	114	0	2381239_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2381239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:186441692(+)-4:186444073(-)__4_186420501_186445501D;SPAN=2381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:114 DP:19 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:0 DR:114 LR:-336.7 LO:336.7);ALT=A[chr4:186444073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	187093527	+	chr4	187098241	+	.	12	0	2384115_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2384115_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:187093527(+)-4:187098241(-)__4_187082001_187107001D;SPAN=4714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:57 GQ:24.2 PL:[24.2, 0.0, 113.3] SR:0 DR:12 LR:-24.17 LO:27.5);ALT=T[chr4:187098241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	187353484	+	chr4	187357165	+	.	46	35	2385581_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GCACACACGGCATTACCCAC;MAPQ=60;MATEID=2385581_2;MATENM=5;NM=3;NUMPARTS=2;SCTG=c_4_187351501_187376501_124C;SPAN=3681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:82 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:35 DR:46 LR:-241.0 LO:241.0);ALT=C[chr4:187357165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	187400707	-	chr4	187401712	+	.	8	0	2384968_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2384968_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:187400707(-)-4:187401712(-)__4_187400501_187425501D;SPAN=1005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr4:187401712[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	187503660	+	chr4	190110405	-	.	10	0	2394124_1	16.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2394124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:187503660(+)-4:190110405(+)__4_190095501_190120501D;SPAN=2606745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:63 GQ:16.1 PL:[16.1, 0.0, 134.9] SR:0 DR:10 LR:-15.94 LO:21.55);ALT=T]chr4:190110405];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	189659676	-	chr6	153323771	+	.	8	0	3079884_1	14.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3079884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:189659676(-)-6:153323771(-)__6_153321001_153346001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=[chr6:153323771[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	190058014	+	chr4	190064273	+	.	99	78	2394515_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ATAAATTACCCAGTCT;MAPQ=60;MATEID=2394515_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_190046501_190071501_297C;SPAN=6259;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:162 DP:41 GQ:43.6 PL:[478.6, 43.6, 0.0] SR:78 DR:99 LR:-478.6 LO:478.6);ALT=T[chr4:190064273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	190191603	+	chr4	190200463	+	.	71	59	2394545_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=GTT;MAPQ=60;MATEID=2394545_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_190193501_190218501_10C;SPAN=8860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:42 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:59 DR:71 LR:-307.0 LO:307.0);ALT=T[chr4:190200463[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	190862226	+	chr4	190864355	+	.	18	16	2396926_1	49.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2396926_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_190855001_190880001_200C;SPAN=2129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:85 GQ:49.7 PL:[49.7, 0.0, 155.3] SR:16 DR:18 LR:-49.59 LO:52.7);ALT=G[chr4:190864355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	153029990	+	chr6	153033790	+	.	42	25	3079342_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTGAAAGAGTATTTATTT;MAPQ=60;MATEID=3079342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_153027001_153052001_82C;SPAN=3800;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:47 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:25 DR:42 LR:-151.8 LO:151.8);ALT=T[chr6:153033790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
