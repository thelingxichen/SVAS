chr12	110252097	+	chr12	110250648	+	.	9	0	7828282_1	6.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7828282_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110250648(-)-12:110252097(+)__12_110250001_110275001D;SPAN=1449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:0 DR:9 LR:-6.139 LO:17.59);ALT=]chr12:110252097]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	110616588	-	chr12	110617822	+	.	12	0	7829743_1	23.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7829743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:110616588(-)-12:110617822(-)__12_110593001_110618001D;SPAN=1234;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:61 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:0 DR:12 LR:-23.09 LO:27.1);ALT=[chr12:110617822[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
