chr1	161342533	-	chr1	161343608	+	.	8	0	588285_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=588285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161342533(-)-1:161343608(-)__1_161332501_161357501D;SPAN=1075;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:122 GQ:6.3 PL:[0.0, 6.3, 306.9] SR:0 DR:8 LR:6.645 LO:13.98);ALT=[chr1:161343608[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	161667711	+	chr1	161800339	+	.	27	0	592513_1	70.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=592513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161667711(+)-1:161800339(-)__1_161798001_161823001D;SPAN=132628;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:70 GQ:70.1 PL:[70.1, 0.0, 99.8] SR:0 DR:27 LR:-70.16 LO:70.45);ALT=C[chr1:161800339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
