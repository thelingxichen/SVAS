chrX	132819582	-	chrX	132820811	+	.	2	2	11389064_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTGTGTGTGTGTGTGT;MAPQ=60;MATEID=11389064_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_132814501_132839501_295C;SPAN=1229;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:2 DR:2 LR:6.844 LO:6.647);ALT=[chrX:132820811[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
