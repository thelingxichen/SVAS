chr5	49695124	+	chr5	49699012	+	ATTTTTTCTATGCCTGGGGACATTATTTTCTATACCATTGCTATCATCTGATTTCAGCTGTTCAATCTGCTCAAATTCTTTCCCCTCAT	3	22	2467381_1	60.0	.	DISC_MAPQ=3;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATTTTTTCTATGCCTGGGGACATTATTTTCTATACCATTGCTATCATCTGATTTCAGCTGTTCAATCTGCTCAAATTCTTTCCCCTCAT;MAPQ=60;MATEID=2467381_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_49686001_49711001_215C;SECONDARY;SPAN=3888;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:58 GQ:60.2 PL:[60.2, 0.0, 80.0] SR:22 DR:3 LR:-60.21 LO:60.37);ALT=C[chr5:49699012[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49699325	+	chr5	49706710	+	.	9	0	2467388_1	17.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=2467388_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:49699325(+)-5:49706710(-)__5_49686001_49711001D;SPAN=7385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=A[chr5:49706710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49706801	+	chr5	49723978	+	GTATTGGGTATACAAGGTGCTTCCTGTTGCACTGACAAGATAATTATTCTCAAGTTGTTCACCATCTTTTTTCCAAGTCACATTTACTGCATTCAAATCCCCAGATGTTGTGAACTGGCATGTGAGATTTACATTAGAAGGCCTTTCTAAAGTGATATTTTTTTCTACTGGCATACTAGAATGTT	0	56	2467398_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTATTGGGTATACAAGGTGCTTCCTGTTGCACTGACAAGATAATTATTCTCAAGTTGTTCACCATCTTTTTTCCAAGTCACATTTACTGCATTCAAATCCCCAGATGTTGTGAACTGGCATGTGAGATTTACATTAGAAGGCCTTTCTAAAGTGATATTTTTTTCTACTGGCATACTAGAATGTT;MAPQ=60;MATEID=2467398_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_49686001_49711001_296C;SPAN=17177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:30 GQ:15 PL:[165.0, 15.0, 0.0] SR:56 DR:0 LR:-165.0 LO:165.0);ALT=T[chr5:49723978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49707218	+	chr5	49723978	+	.	5	40	2467298_1	99.0	.	DISC_MAPQ=30;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2467298_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_49710501_49735501_252C;SPAN=16760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:40 GQ:12 PL:[132.0, 12.0, 0.0] SR:40 DR:5 LR:-132.0 LO:132.0);ALT=C[chr5:49723978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49707267	+	chr5	49736873	+	.	12	0	2467447_1	28.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=2467447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:49707267(+)-5:49736873(-)__5_49735001_49760001D;SPAN=29606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:40 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:0 DR:12 LR:-28.78 LO:29.66);ALT=T[chr5:49736873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49724063	+	chr5	49736874	+	.	60	84	2467449_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2467449_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_49735001_49760001_256C;SPAN=12811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:42 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:84 DR:60 LR:-326.8 LO:326.8);ALT=T[chr5:49736874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49822803	+	chr5	49949875	+	.	8	0	2467839_1	16.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2467839_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:49822803(+)-5:49949875(-)__5_49931001_49956001D;SPAN=127072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:0 DR:8 LR:-16.11 LO:18.33);ALT=G[chr5:49949875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49935251	+	chr5	49949853	+	.	10	0	2467853_1	20.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=2467853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:49935251(+)-5:49949853(-)__5_49931001_49956001D;SPAN=14602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=C[chr5:49949853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49963020	+	chr5	50055474	+	ATTTCAGATACTCTGACTCCACCTTTACTTTTACCTACGTTGGCGGCCCCAGAAGTGTATCCTACTCAGTACATGTATCTGAAGATTACC	2	16	2467792_1	44.0	.	DISC_MAPQ=25;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=ATTTCAGATACTCTGACTCCACCTTTACTTTTACCTACGTTGGCGGCCCCAGAAGTGTATCCTACTCAGTACATGTATCTGAAGATTACC;MAPQ=60;MATEID=2467792_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_49955501_49980501_156C;SECONDARY;SPAN=92454;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:30 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:16 DR:2 LR:-44.89 LO:44.89);ALT=G[chr5:50055474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	49963020	+	chr5	50045983	+	ATTTCAGATACTCTGACTCCACCTTTACTTTTACCTACGTTGGCGGCCCCAGA	2	15	2467895_1	41.0	.	DISC_MAPQ=46;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATTTCAGATACTCTGACTCCACCTTTACTTTTACCTACGTTGGCGGCCCCAGA;MAPQ=60;MATEID=2467895_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_50029001_50054001_171C;SPAN=82963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:28 GQ:25.4 PL:[41.9, 0.0, 25.4] SR:15 DR:2 LR:-42.13 LO:42.13);ALT=G[chr5:50045983[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	50093067	+	chr5	50111265	+	.	2	2	2468305_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2468305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_50102501_50127501_235C;SPAN=18198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:24 GQ:6.8 PL:[6.8, 0.0, 49.7] SR:2 DR:2 LR:-6.702 LO:8.712);ALT=G[chr5:50111265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	50129882	+	chr5	50137800	+	TGATCACCTCATCTGACCTGCACAAACATGGAGAGATATGGGTTGTCCCCAATACTGACCATGTCTGCACACGATTCTTTTTCGT	3	13	2467943_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGATCACCTCATCTGACCTGCACAAACATGGAGAGATATGGGTTGTCCCCAATACTGACCATGTCTGCACACGATTCTTTTTCGT;MAPQ=60;MATEID=2467943_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_50127001_50152001_42C;SPAN=7918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:13 DR:3 LR:-34.89 LO:36.48);ALT=G[chr5:50137800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	50130849	+	chr5	50137800	+	.	4	7	2467945_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2467945_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_50127001_50152001_42C;SPAN=6951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:7 DR:4 LR:-21.68 LO:25.03);ALT=T[chr5:50137800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
