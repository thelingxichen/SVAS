chr22	49425468	+	chr2	85714118	+	G	8	28	1136534_1	75.0	.	DISC_MAPQ=11;EVDNC=ASDIS;INSERTION=G;MAPQ=11;MATEID=1136534_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_85701001_85726001_257C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:31 DP:98 GQ:75.8 PL:[75.8, 0.0, 161.6] SR:28 DR:8 LR:-75.78 LO:77.5);ALT=]chr22:49425468]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	86137592	+	chr2	86138755	-	.	8	0	1137985_1	0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=1137985_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:86137592(+)-2:86138755(+)__2_86117501_86142501D;SPAN=1163;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:142 GQ:11.7 PL:[0.0, 11.7, 366.3] SR:0 DR:8 LR:12.06 LO:13.44);ALT=A]chr2:86138755];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	86283455	-	chr2	86323000	+	GCATGCCTGTA	18	52	1139281_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=ATCCCAGCTACTCGGGAGGCTGAGGCAGGAGAATTGCTT;INSERTION=GCATGCCTGTA;MAPQ=60;MATEID=1139281_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_2_86264501_86289501_597C;SPAN=39545;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:73 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:52 DR:18 LR:-214.6 LO:214.6);ALT=[chr2:86323000[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	49715779	+	chr22	49717444	+	.	0	71	10914155_1	99.0	.	EVDNC=ASSMB;HOMSEQ=T;MAPQ=60;MATEID=10914155_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_49710501_49735501_145C;SPAN=1665;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:24 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:71 DR:0 LR:-208.0 LO:208.0);ALT=T[chr22:49717444[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
