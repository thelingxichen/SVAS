chr16	65551833	+	chr16	65553090	+	.	65	52	9371810_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=60;MATEID=9371810_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_65537501_65562501_354C;SPAN=1257;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:98 DP:82 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:52 DR:65 LR:-290.5 LO:290.5);ALT=C[chr16:65553090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
