chr6	666376	+	chr6	667822	+	.	0	126	3979689_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3979689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_661501_686501_382C;SPAN=1446;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:126 DP:52 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:126 DR:0 LR:-373.0 LO:373.0);ALT=A[chr6:667822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	736236	+	chr20	61823936	-	.	18	0	3980540_1	52.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3980540_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:736236(+)-20:61823936(+)__6_735001_760001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:18 DP:15 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=G]chr20:61823936];VARTYPE=BND:TRX-hh;JOINTYPE=hh
