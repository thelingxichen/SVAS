chr11	30344750	+	chr11	30352431	+	.	19	4	4808097_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4808097_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_11_30331001_30356001_149C;SPAN=7681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:94 GQ:44 PL:[44.0, 0.0, 182.6] SR:4 DR:19 LR:-43.85 LO:48.74);ALT=G[chr11:30352431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
