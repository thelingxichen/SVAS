chr11	69982555	+	chr11	69984488	+	.	96	59	4906428_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTC;MAPQ=60;MATEID=4906428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_69972001_69997001_240C;SPAN=1933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:29 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:59 DR:96 LR:-399.4 LO:399.4);ALT=C[chr11:69984488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
