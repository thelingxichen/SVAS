chr12	123668122	+	chr12	123669280	-	.	8	0	7881755_1	0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=7881755_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123668122(+)-12:123669280(+)__12_123651501_123676501D;SPAN=1158;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:142 GQ:11.7 PL:[0.0, 11.7, 366.3] SR:0 DR:8 LR:12.06 LO:13.44);ALT=A]chr12:123669280];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	124368288	-	chr12	124369368	+	.	3	4	7886019_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATGCAGAA;MAPQ=60;MATEID=7886019_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124362001_124387001_14C;SPAN=1080;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:138 GQ:17.4 PL:[0.0, 17.4, 369.6] SR:4 DR:3 LR:17.58 LO:9.393);ALT=[chr12:124369368[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
