chr2	79253983	+	chr2	79385800	-	.	22	0	1110891_1	59.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1110891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:79253983(+)-2:79385800(+)__2_79233001_79258001D;SPAN=131817;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:49 GQ:59.3 PL:[59.3, 0.0, 59.3] SR:0 DR:22 LR:-59.35 LO:59.35);ALT=G]chr2:79385800];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	79254085	-	chr2	79385657	+	.	16	0	1110892_1	36.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1110892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:79254085(-)-2:79385657(-)__2_79233001_79258001D;SPAN=131572;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:0 DR:16 LR:-36.83 LO:38.71);ALT=[chr2:79385657[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
