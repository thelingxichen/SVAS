chr5	169064373	+	chr5	169081406	+	.	6	3	2639476_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2639476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_169050001_169075001_53C;SPAN=17033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:31 GQ:14.9 PL:[14.9, 0.0, 57.8] SR:3 DR:6 LR:-14.71 LO:16.28);ALT=G[chr5:169081406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	169081490	+	chr5	169101300	+	ACTGGTATAGGGGATACCTCATAAAGCACAAAATGTTACAGGGCATTTTTCCTAAGTCATTTATCCACATCAAGGAAGTGACAGTTGAGAAAAGAAGAAATACTGAGAACATCATTCCTGCAGAAATTCCTCTGGCACAAGAAGTGACAACGACACTTTGGGAATGGGGAAGCATCTGGAAACAACTCTATGT	0	13	2639357_1	33.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ACTGGTATAGGGGATACCTCATAAAGCACAAAATGTTACAGGGCATTTTTCCTAAGTCATTTATCCACATCAAGGAAGTGACAGTTGAGAAAAGAAGAAATACTGAGAACATCATTCCTGCAGAAATTCCTCTGGCACAAGAAGTGACAACGACACTTTGGGAATGGGGAAGCATCTGGAAACAACTCTATGT;MAPQ=60;MATEID=2639357_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_5_169074501_169099501_119C;SPAN=19810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:13 DR:0 LR:-33.7 LO:33.85);ALT=G[chr5:169101300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	169675825	+	chr5	169677733	+	.	4	2	2640543_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2640543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_169662501_169687501_253C;SPAN=1908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:59 GQ:3.8 PL:[3.8, 0.0, 139.1] SR:2 DR:4 LR:-3.821 LO:11.68);ALT=T[chr5:169677733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
