chr15	48623989	+	chr15	48626611	+	.	22	0	5945796_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5945796_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:48623989(+)-15:48626611(-)__15_48608001_48633001D;SPAN=2622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:77 GQ:51.8 PL:[51.8, 0.0, 134.3] SR:0 DR:22 LR:-51.76 LO:53.82);ALT=C[chr15:48626611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	48624603	+	chr15	48626612	+	CTCCACGGTCA	50	125	5945802_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;INSERTION=CTCCACGGTCA;MAPQ=60;MATEID=5945802_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_48608001_48633001_62C;SPAN=2009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:130 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:125 DR:50 LR:-448.9 LO:448.9);ALT=G[chr15:48626612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49330011	+	chr15	49338593	+	.	8	0	5946743_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5946743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:49330011(+)-15:49338593(-)__15_49318501_49343501D;SPAN=8582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:0 DR:8 LR:-9.611 LO:16.46);ALT=A[chr15:49338593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49431851	+	chr15	49437158	+	AACTTGAAGTTAATCTTAATCATTTGTTTCAGTGCTTTAAATCCCCATTCTCCTTTTTCACCTTCAAGTTCCA	0	49	5946782_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AAACCT;INSERTION=AACTTGAAGTTAATCTTAATCATTTGTTTCAGTGCTTTAAATCCCCATTCTCCTTTTTCACCTTCAAGTTCCA;MAPQ=60;MATEID=5946782_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_49416501_49441501_244C;SPAN=5307;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:59 GQ:2.7 PL:[148.5, 2.7, 0.0] SR:49 DR:0 LR:-155.5 LO:155.5);ALT=C[chr15:49437158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49431894	+	chr15	49447727	+	.	11	0	5946888_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5946888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:49431894(+)-15:49447727(-)__15_49441001_49466001D;SPAN=15833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:30 GQ:28.1 PL:[28.1, 0.0, 44.6] SR:0 DR:11 LR:-28.18 LO:28.39);ALT=C[chr15:49447727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49436548	+	chr15	49447720	+	.	23	0	5946890_1	69.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5946890_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:49436548(+)-15:49447720(-)__15_49441001_49466001D;SPAN=11172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:24 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:23 LR:-69.32 LO:69.32);ALT=A[chr15:49447720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49437304	+	chr15	49447726	+	.	22	0	5946891_1	64.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5946891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:49437304(+)-15:49447726(-)__15_49441001_49466001D;SPAN=10422;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:29 GQ:5.3 PL:[64.7, 0.0, 5.3] SR:0 DR:22 LR:-67.69 LO:67.69);ALT=G[chr15:49447726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	49913345	+	chr15	49917306	+	.	16	0	5947461_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5947461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:49913345(+)-15:49917306(-)__15_49906501_49931501D;SPAN=3961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:52 GQ:38.9 PL:[38.9, 0.0, 85.1] SR:0 DR:16 LR:-38.73 LO:39.77);ALT=T[chr15:49917306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50211148	+	chr15	50212443	+	.	2	3	5947789_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5947789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_50200501_50225501_190C;SPAN=1295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:55 GQ:1.5 PL:[0.0, 1.5, 135.3] SR:3 DR:2 LR:1.697 LO:7.178);ALT=C[chr15:50212443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50331026	+	chr15	50339548	+	ATAGTCATCTGTGGCATCTTTGACAGCTGTCATAGTTATCACCAGGACCAAAGGCACAATGGTGGTAAACCAGGTCAAGGAGGAAATTTCTGGAATTAG	3	20	5947979_1	55.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATAGTCATCTGTGGCATCTTTGACAGCTGTCATAGTTATCACCAGGACCAAAGGCACAATGGTGGTAAACCAGGTCAAGGAGGAAATTTCTGGAATTAG;MAPQ=60;MATEID=5947979_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_50323001_50348001_280C;SPAN=8522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:53 GQ:55.1 PL:[55.1, 0.0, 71.6] SR:20 DR:3 LR:-54.96 LO:55.11);ALT=A[chr15:50339548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50336892	+	chr15	50339548	+	.	4	9	5947983_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5947983_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_15_50323001_50348001_280C;SPAN=2656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:44 GQ:27.8 PL:[27.8, 0.0, 77.3] SR:9 DR:4 LR:-27.69 LO:29.07);ALT=G[chr15:50339548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50339662	+	chr15	50366323	+	.	0	23	5947987_1	69.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5947987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_50323001_50348001_97C;SPAN=26661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:24 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:23 DR:0 LR:-69.32 LO:69.32);ALT=C[chr15:50366323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50366383	+	chr15	50399136	+	.	0	32	5948118_1	95.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5948118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_50396501_50421501_44C;SPAN=32753;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:33 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:32 DR:0 LR:-95.72 LO:95.72);ALT=C[chr15:50399136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50366431	+	chr15	50411358	+	.	25	0	5948119_1	71.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5948119_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:50366431(+)-15:50411358(-)__15_50396501_50421501D;SPAN=44927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:40 GQ:25.4 PL:[71.6, 0.0, 25.4] SR:0 DR:25 LR:-72.9 LO:72.9);ALT=A[chr15:50411358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	50399207	+	chr15	50411318	+	.	22	18	5948125_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5948125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_50396501_50421501_203C;SPAN=12111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:62 GQ:65.9 PL:[82.4, 0.0, 65.9] SR:18 DR:22 LR:-82.3 LO:82.3);ALT=T[chr15:50411318[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	51041944	+	chr15	51057665	+	.	0	10	5949356_1	16.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5949356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_51033501_51058501_145C;SPAN=15721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:10 DR:0 LR:-16.21 LO:21.62);ALT=C[chr15:51057665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
