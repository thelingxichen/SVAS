chr12	43977460	+	chr12	43979550	+	.	47	40	5168014_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGACATTCCA;MAPQ=60;MATEID=5168014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_43977501_44002501_97C;SPAN=2090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:19 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:40 DR:47 LR:-224.5 LO:224.5);ALT=A[chr12:43979550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	44142415	+	chr12	44148139	+	.	0	8	5168526_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5168526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_44124501_44149501_128C;SPAN=5724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:8 DR:0 LR:-8.798 LO:16.28);ALT=G[chr12:44148139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	44149036	+	chr12	44152502	+	.	10	0	5168535_1	21.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=5168535_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:44149036(+)-12:44152502(-)__12_44124501_44149501D;SPAN=3466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:0 DR:10 LR:-21.63 LO:23.53);ALT=T[chr12:44152502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	44152871	+	chr12	44161902	+	.	8	0	5168448_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5168448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:44152871(+)-12:44161902(-)__12_44149001_44174001D;SPAN=9031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:0 DR:8 LR:-7.985 LO:16.11);ALT=T[chr12:44161902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
