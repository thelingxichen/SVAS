chr16	89937987	+	chr16	89721211	+	.	45	26	9457368_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=C;MAPQ=48;MATEID=9457368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_89719001_89744001_389C;SPAN=216776;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:64 DP:29 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:26 DR:45 LR:-188.1 LO:188.1);ALT=]chr16:89937987]C;VARTYPE=BND:DUP-th;JOINTYPE=th
