chr1	68365458	-	chr1	68367758	+	.	8	0	328053_1	0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=328053_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:68365458(-)-1:68367758(-)__1_68355001_68380001D;SPAN=2300;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:124 GQ:6.9 PL:[0.0, 6.9, 313.5] SR:0 DR:8 LR:7.187 LO:13.93);ALT=[chr1:68367758[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
