chr12	95365397	+	chr12	95387945	+	.	0	35	5295595_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5295595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95378501_95403501_141C;SPAN=22548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:47 GQ:10.4 PL:[102.8, 0.0, 10.4] SR:35 DR:0 LR:-107.1 LO:107.1);ALT=C[chr12:95387945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95365451	+	chr12	95397369	+	.	14	0	5295597_1	36.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5295597_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:95365451(+)-12:95397369(-)__12_95378501_95403501D;SPAN=31918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:36 GQ:36.5 PL:[36.5, 0.0, 49.7] SR:0 DR:14 LR:-36.46 LO:36.59);ALT=A[chr12:95397369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95388034	+	chr12	95396514	+	.	0	49	5295625_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5295625_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95378501_95403501_377C;SPAN=8480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:94 GQ:90.2 PL:[136.4, 0.0, 90.2] SR:49 DR:0 LR:-136.7 LO:136.7);ALT=C[chr12:95396514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95388083	+	chr12	95397373	+	.	45	0	5295626_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5295626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:95388083(+)-12:95397373(-)__12_95378501_95403501D;SPAN=9290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:67 GQ:31.4 PL:[130.4, 0.0, 31.4] SR:0 DR:45 LR:-133.7 LO:133.7);ALT=A[chr12:95397373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95835595	-	chr12	95836670	+	.	9	0	5296832_1	8.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5296832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:95835595(-)-12:95836670(-)__12_95819501_95844501D;SPAN=1075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:0 DR:9 LR:-8.577 LO:18.05);ALT=[chr12:95836670[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	95868107	+	chr12	95869846	+	.	39	28	5297230_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCAGG;MAPQ=60;MATEID=5297230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95844001_95869001_374C;SPAN=1739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:43 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:28 DR:39 LR:-161.7 LO:161.7);ALT=G[chr12:95869846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95869954	+	chr12	95876989	+	.	0	19	5296979_1	37.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5296979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95868501_95893501_382C;SPAN=7035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:94 GQ:37.4 PL:[37.4, 0.0, 189.2] SR:19 DR:0 LR:-37.25 LO:43.16);ALT=G[chr12:95876989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95877094	+	chr12	95887830	+	.	9	0	5296992_1	3.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5296992_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:95877094(+)-12:95887830(-)__12_95868501_95893501D;SPAN=10736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:0 DR:9 LR:-3.429 LO:17.14);ALT=A[chr12:95887830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	95879758	+	chr12	95887831	+	.	0	7	5296999_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5296999_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_95868501_95893501_67C;SPAN=8073;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=G[chr12:95887831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96233592	+	chr12	96236328	+	.	30	15	5298503_1	15.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TCCACAGTTTT;MAPQ=60;MATEID=5298503_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96211501_96236501_143C;SPAN=2736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:455 GQ:15.6 PL:[15.6, 0.0, 1088.0] SR:15 DR:30 LR:-15.37 LO:79.9);ALT=T[chr12:96236328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96252854	+	chr12	96254945	+	.	76	50	5298284_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5298284_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96236001_96261001_57C;SPAN=2091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:121 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:50 DR:76 LR:-354.2 LO:354.2);ALT=G[chr12:96254945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96340355	+	chr12	96342955	+	.	98	54	5298847_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGAGACTGC;MAPQ=60;MATEID=5298847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96334001_96359001_43C;SPAN=2600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:120 DP:60 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:54 DR:98 LR:-356.5 LO:356.5);ALT=C[chr12:96342955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96394884	+	chr12	96396737	+	.	3	20	5298666_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5298666_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96383001_96408001_198C;SPAN=1853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:82 GQ:47.3 PL:[47.3, 0.0, 149.6] SR:20 DR:3 LR:-47.11 LO:50.19);ALT=C[chr12:96396737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96421342	+	chr12	96422833	+	.	2	4	5298616_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5298616_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96407501_96432501_229C;SPAN=1491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:72 GQ:2.7 PL:[0.0, 2.7, 178.2] SR:4 DR:2 LR:3.002 LO:8.869);ALT=T[chr12:96422833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96422964	+	chr12	96429137	+	.	0	28	5298620_1	70.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=5298620_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96407501_96432501_140C;SPAN=6173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:83 GQ:70.1 PL:[70.1, 0.0, 129.5] SR:28 DR:0 LR:-69.94 LO:70.97);ALT=C[chr12:96429137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	96588486	+	chr12	96617342	+	.	3	4	5299353_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTA;MAPQ=60;MATEID=5299353_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_96603501_96628501_289C;SPAN=28856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:34 GQ:7.4 PL:[7.4, 0.0, 73.4] SR:4 DR:3 LR:-7.294 LO:10.59);ALT=A[chr12:96617342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
