chr18	36709399	+	chr13	60002628	+	.	6	33	8101348_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACACACACACACACACAATGGAATACTACTCAGCCATAAAAAGGAATGAA;MAPQ=60;MATEID=8101348_2;MATENM=8;NM=2;NUMPARTS=2;SCTG=c_13_60000501_60025501_1C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:39 DP:60 GQ:33.2 PL:[112.4, 0.0, 33.2] SR:33 DR:6 LR:-114.9 LO:114.9);ALT=]chr18:36709399]A;VARTYPE=BND:TRX-th;JOINTYPE=th
