chr7	127214969	+	chr7	127217982	+	C	0	41	5276157_1	99.0	.	EVDNC=ASSMB;INSERTION=C;MAPQ=60;MATEID=5276157_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_127204001_127229001_219C;SPAN=3013;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:41 DP:15 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:41 DR:0 LR:-118.8 LO:118.8);ALT=A[chr7:127217982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
