chr2	179296983	+	chr2	179300872	+	.	3	2	1108688_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1108688_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_179291001_179316001_259C;SPAN=3889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:2 DR:3 LR:4.677 LO:6.851);ALT=T[chr2:179300872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	179402419	+	chr2	179403422	+	.	0	5	1109091_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=1109091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_179389001_179414001_281C;SPAN=1003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:75 GQ:3.6 PL:[0.0, 3.6, 188.1] SR:5 DR:0 LR:3.814 LO:8.777);ALT=G[chr2:179403422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
