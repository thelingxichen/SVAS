chr4	130066147	+	chr4	130068441	+	.	15	0	2914091_1	42.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2914091_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:130066147(+)-4:130068441(-)__4_130046001_130071001D;SPAN=2294;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:15 DP:11 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=A[chr4:130068441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	130216516	+	chr4	130219483	+	.	68	28	2914542_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CATAGCTGGCAATTTCT;MAPQ=60;MATEID=2914542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_130193001_130218001_239C;SPAN=2967;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:34 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:28 DR:68 LR:-247.6 LO:247.6);ALT=T[chr4:130219483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
