chr16	28096255	-	chr16	28097320	+	.	7	1	9246446_1	0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AGCCAGGCAT;MAPQ=60;MATEID=9246446_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_28077001_28102001_120C;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:114 GQ:4.2 PL:[0.0, 4.2, 283.8] SR:1 DR:7 LR:4.477 LO:14.23);ALT=[chr16:28097320[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	28284677	+	chr16	28285741	-	.	8	0	9247527_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=9247527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:28284677(+)-16:28285741(+)__16_28273001_28298001D;SPAN=1064;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:166 GQ:18.4 PL:[0.0, 18.4, 439.0] SR:0 DR:8 LR:18.57 LO:12.89);ALT=G]chr16:28285741];VARTYPE=BND:INV-hh;JOINTYPE=hh
