chr3	63147962	-	chr3	63149523	+	.	10	0	1449627_1	1.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=1449627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:63147962(-)-3:63149523(-)__3_63136501_63161501D;SPAN=1561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:117 GQ:1.4 PL:[1.4, 0.0, 281.9] SR:0 DR:10 LR:-1.312 LO:18.67);ALT=[chr3:63149523[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	63820901	+	chr3	63823652	+	TATCTTCAACACTTTCTTTAATGTGTGAAAGATGCTCTAATTCTTTTCCCAGAGCCTCTAGTTCCTTTAATGTCTCATGCCTGTCTGGATGGTGCTGAATCACTTTTGCCAAAGCATCATATT	4	17	1451739_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TATCTTCAACACTTTCTTTAATGTGTGAAAGATGCTCTAATTCTTTTCCCAGAGCCTCTAGTTCCTTTAATGTCTCATGCCTGTCTGGATGGTGCTGAATCACTTTTGCCAAAGCATCATATT;MAPQ=60;MATEID=1451739_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_63822501_63847501_408C;SPAN=2751;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:17 DR:4 LR:-45.01 LO:45.06);ALT=T[chr3:63823652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63823742	+	chr3	63825332	+	TTCCTTGTAAATTTTTTCATAATTTTCCATTTCTCTGAGATTCATATCATATACTAGTAAAGTTTTGCCCATTGAAAATTCACATTGAGACAGCGTGCTCAGCATACGTTGGTACTGGCTATAT	3	66	1451747_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTCCTTGTAAATTTTTTCATAATTTTCCATTTCTCTGAGATTCATATCATATACTAGTAAAGTTTTGCCCATTGAAAATTCACATTGAGACAGCGTGCTCAGCATACGTTGGTACTGGCTATAT;MAPQ=60;MATEID=1451747_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_63822501_63847501_136C;SPAN=1590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:100 GQ:48.8 PL:[194.0, 0.0, 48.8] SR:66 DR:3 LR:-198.9 LO:198.9);ALT=T[chr3:63825332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63823783	+	chr3	63849446	+	.	13	0	1451748_1	31.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1451748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:63823783(+)-3:63849446(-)__3_63822501_63847501D;SPAN=25663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:44 GQ:31.1 PL:[31.1, 0.0, 74.0] SR:0 DR:13 LR:-30.99 LO:32.03);ALT=A[chr3:63849446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63824176	+	chr3	63825332	+	.	0	35	1451848_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1451848_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_3_63847001_63872001_40C;SPAN=1156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:0 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:35 DR:0 LR:-102.3 LO:102.3);ALT=C[chr3:63825332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63824224	+	chr3	63849446	+	.	44	0	1451849_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1451849_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:63824224(+)-3:63849446(-)__3_63847001_63872001D;SPAN=25222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:35 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:0 DR:44 LR:-128.7 LO:128.7);ALT=A[chr3:63849446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63825472	+	chr3	63849446	+	.	28	0	1451850_1	83.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1451850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:63825472(+)-3:63849446(-)__3_63847001_63872001D;SPAN=23974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:35 GQ:0.5 PL:[83.0, 0.0, 0.5] SR:0 DR:28 LR:-87.65 LO:87.65);ALT=T[chr3:63849446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	63847469	-	chr3	63848566	+	.	8	0	1451855_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1451855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:63847469(-)-3:63848566(-)__3_63847001_63872001D;SPAN=1097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=[chr3:63848566[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	63996631	+	chr3	63999114	+	.	3	10	1452362_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1452362_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_63994001_64019001_61C;SPAN=2483;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:107 GQ:14 PL:[14.0, 0.0, 245.0] SR:10 DR:3 LR:-13.92 LO:26.38);ALT=C[chr3:63999114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
