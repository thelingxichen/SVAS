chr12	127579217	+	chr12	127585803	+	.	19	0	7900537_1	40.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7900537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:127579217(+)-12:127585803(-)__12_127571501_127596501D;SPAN=6586;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:19 DP:84 GQ:40.1 PL:[40.1, 0.0, 162.2] SR:0 DR:19 LR:-39.96 LO:44.22);ALT=A[chr12:127585803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
