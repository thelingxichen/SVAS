chr21	23275815	+	chr21	25180328	+	.	9	0	7134378_1	26.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=7134378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:23275815(+)-21:25180328(-)__21_23250501_23275501D;SPAN=1904513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:0 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=C[chr21:25180328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	23626258	+	chr21	29293617	-	.	45	0	7148592_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7148592_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:23626258(+)-21:29293617(+)__21_29277501_29302501D;SPAN=5667359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:32 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=T]chr21:29293617];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr21	25801154	+	chr21	25810564	+	.	11	0	7139926_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7139926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:25801154(+)-21:25810564(-)__21_25798501_25823501D;SPAN=9410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:78 GQ:15.2 PL:[15.2, 0.0, 173.6] SR:0 DR:11 LR:-15.18 LO:23.09);ALT=C[chr21:25810564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
