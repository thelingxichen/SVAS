chr15	29020454	-	chrX	139983587	+	.	2	5	8811698_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCCTGGCTAA;MAPQ=60;MATEID=8811698_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_29008001_29033001_459C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:81 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:5 DR:2 LR:5.44 LO:8.605);ALT=[chrX:139983587[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
