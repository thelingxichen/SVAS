chr6	119013928	+	chr6	119011719	+	.	56	49	4369985_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=4369985_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_118996501_119021501_80C;SPAN=2209;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:61 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:49 DR:56 LR:-237.7 LO:237.7);ALT=]chr6:119013928]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	119012288	+	chr6	119013928	+	TACATTGTCA	0	52	4369990_1	99.0	.	EVDNC=ASSMB;INSERTION=TACATTGTCA;MAPQ=60;MATEID=4369990_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_118996501_119021501_11C;SPAN=1640;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:66 GQ:5.3 PL:[153.8, 0.0, 5.3] SR:52 DR:0 LR:-161.9 LO:161.9);ALT=A[chr6:119013928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
