chr4	80888062	+	chr4	80894092	+	.	51	31	2052377_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAATAGGGCGTCCG;MAPQ=60;MATEID=2052377_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_80874501_80899501_66C;SPAN=6030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:64 GQ:18 PL:[198.0, 18.0, 0.0] SR:31 DR:51 LR:-198.0 LO:198.0);ALT=G[chr4:80894092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
