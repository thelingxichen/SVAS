chr12	84593114	+	chr12	84596012	+	.	83	57	7779365_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GCCTCA;MAPQ=60;MATEID=7779365_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_84574001_84599001_55C;SPAN=2898;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:112 DP:21 GQ:30 PL:[330.0, 30.0, 0.0] SR:57 DR:83 LR:-330.1 LO:330.1);ALT=A[chr12:84596012[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
