chrX	147382685	+	chrX	147408470	+	.	9	0	11418383_1	18.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=11418383_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:147382685(+)-23:147408470(-)__23_147367501_147392501D;SPAN=25785;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.6 LO:20.81);ALT=A[chrX:147408470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	147509696	+	chrX	147511236	+	TG	82	59	11418302_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TG;MAPQ=60;MATEID=11418302_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_147490001_147515001_219C;SPAN=1540;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:114 DP:22 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:59 DR:82 LR:-336.7 LO:336.7);ALT=G[chrX:147511236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
