chr1	53594139	+	chr1	53595603	+	.	30	0	264882_1	77.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=264882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53594139(+)-1:53595603(-)__1_53581501_53606501D;SPAN=1464;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:80 GQ:77.3 PL:[77.3, 0.0, 116.9] SR:0 DR:30 LR:-77.36 LO:77.8);ALT=A[chr1:53595603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53891506	+	chr1	55489956	+	.	9	0	266445_1	11.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=266445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:53891506(+)-1:55489956(-)__1_53875501_53900501D;SPAN=1598450;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:0 DR:9 LR:-11.83 LO:18.75);ALT=A[chr1:55489956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	53896738	-	chr1	53897790	+	.	6	3	266471_1	0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CACACACACACACACACACA;MAPQ=60;MATEID=266471_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_53875501_53900501_402C;SPAN=1052;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:7 DP:148 GQ:16.9 PL:[0.0, 16.9, 392.7] SR:3 DR:6 LR:16.99 LO:11.22);ALT=[chr1:53897790[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	55092274	+	chr1	55095967	+	.	81	54	271821_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=271821_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_55076001_55101001_155C;SPAN=3693;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:84 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:54 DR:81 LR:-326.8 LO:326.8);ALT=G[chr1:55095967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	55927721	+	chr1	55929226	+	.	56	43	275757_1	99.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=TCATAG;MAPQ=22;MATEID=275757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_55909001_55934001_440C;SPAN=1505;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:78 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:43 DR:56 LR:-237.7 LO:237.7);ALT=G[chr1:55929226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	56831124	+	chr1	56834962	+	.	42	41	279068_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAGAACCACTGCCTC;MAPQ=60;MATEID=279068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_56815501_56840501_118C;SPAN=3838;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:66 DP:89 GQ:22.1 PL:[193.7, 0.0, 22.1] SR:41 DR:42 LR:-201.7 LO:201.7);ALT=C[chr1:56834962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
