chr14	50540150	+	chr14	50541658	+	.	80	0	8493794_1	99.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=8493794_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:50540150(+)-14:50541658(-)__14_50519001_50544001D;SPAN=1508;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:10 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:0 DR:80 LR:-237.7 LO:237.7);ALT=A[chr14:50541658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
