chr4	178361583	+	chr4	178363403	+	.	15	5	2354984_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2354984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_178360001_178385001_100C;SPAN=1820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:122 GQ:26.6 PL:[26.6, 0.0, 267.5] SR:5 DR:15 LR:-26.37 LO:38.16);ALT=G[chr4:178363403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
