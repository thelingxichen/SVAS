chr3	15845173	+	chr3	15846737	+	.	99	61	1861459_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=ATG;MAPQ=60;MATEID=1861459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15827001_15852001_70C;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:130 DP:31 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:61 DR:99 LR:-386.2 LO:386.2);ALT=G[chr3:15846737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	16239409	+	chr3	16241210	+	.	77	44	1863434_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1863434_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_16219001_16244001_15C;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:105 DP:74 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:44 DR:77 LR:-310.3 LO:310.3);ALT=T[chr3:16241210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
