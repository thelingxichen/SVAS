chr2	152132380	+	chr2	152135342	+	.	5	6	1043302_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1043302_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_152120501_152145501_167C;SPAN=2962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:6 DR:5 LR:-14.05 LO:21.05);ALT=T[chr2:152135342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	152135506	+	chr2	152139381	+	GGAATTCTTTGGTAGCCTCTTGTAACTCCGTTTCAAGCTTTTGGATCTCCTTCTTTAGTTGAATATTTTTCTTTGTAATTTCATCAATTAGTC	4	32	1043311_1	94.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTTA;INSERTION=GGAATTCTTTGGTAGCCTCTTGTAACTCCGTTTCAAGCTTTTGGATCTCCTTCTTTAGTTGAATATTTTTCTTTGTAATTTCATCAATTAGTC;MAPQ=60;MATEID=1043311_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_152120501_152145501_62C;SPAN=3875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:65 GQ:61.7 PL:[94.7, 0.0, 61.7] SR:32 DR:4 LR:-94.96 LO:94.96);ALT=T[chr2:152139381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	152135554	+	chr2	152146102	+	.	16	0	1043435_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1043435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:152135554(+)-2:152146102(-)__2_152145001_152170001D;SPAN=10548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:46 GQ:40.4 PL:[40.4, 0.0, 70.1] SR:0 DR:16 LR:-40.35 LO:40.82);ALT=A[chr2:152146102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	152138596	+	chr2	152146105	+	.	14	0	1043437_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1043437_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:152138596(+)-2:152146105(-)__2_152145001_152170001D;SPAN=7509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:48 GQ:33.2 PL:[33.2, 0.0, 82.7] SR:0 DR:14 LR:-33.21 LO:34.4);ALT=C[chr2:152146105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
