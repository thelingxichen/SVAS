chr13	95900008	+	chr13	95953492	+	.	0	9	5606558_1	22.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=5606558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_95942001_95967001_13C;SPAN=53484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:9 DR:0 LR:-22.12 LO:22.58);ALT=C[chr13:95953492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	96329594	+	chr13	96361479	+	.	12	15	5607687_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=5607687_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_96358501_96383501_223C;SPAN=31885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:37 GQ:29.6 PL:[59.3, 0.0, 29.6] SR:15 DR:12 LR:-59.79 LO:59.79);ALT=G[chr13:96361479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
