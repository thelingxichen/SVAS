chr6	21252871	+	chr2	67416846	+	.	16	0	1061711_1	35.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1061711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:67416846(-)-6:21252871(+)__2_67399501_67424501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:64 GQ:35.6 PL:[35.6, 0.0, 118.1] SR:0 DR:16 LR:-35.48 LO:38.04);ALT=]chr6:21252871]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	22003245	+	chr6	22004796	-	.	8	0	4072529_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4072529_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:22003245(+)-6:22004796(+)__6_22001001_22026001D;SPAN=1551;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:132 GQ:9 PL:[0.0, 9.0, 336.6] SR:0 DR:8 LR:9.354 LO:13.7);ALT=T]chr6:22004796];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	22050976	+	chr6	22054308	+	.	129	0	4073036_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4073036_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:22050976(+)-6:22054308(-)__6_22025501_22050501D;SPAN=3332;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:129 DP:0 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:0 DR:129 LR:-382.9 LO:382.9);ALT=G[chr6:22054308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
