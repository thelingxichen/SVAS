chr11	1915274	+	chr11	1936956	+	ATG	97	26	6622465_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=ATG;MAPQ=47;MATEID=6622465_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_1935501_1960501_270C;SPAN=21682;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:116 DP:56 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:26 DR:97 LR:-343.3 LO:343.3);ALT=G[chr11:1936956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	2077974	+	chr11	2073453	+	.	10	0	6623059_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6623059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:2073453(-)-11:2077974(+)__11_2058001_2083001D;SPAN=4521;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=]chr11:2077974]T;VARTYPE=BND:DUP-th;JOINTYPE=th
