chr1	48850099	+	chr8	21879137	-	.	10	0	244976_1	18.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=244976_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:48850099(+)-8:21879137(+)__1_48828501_48853501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:0 DR:10 LR:-18.65 LO:22.38);ALT=G]chr8:21879137];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	21170008	+	chr8	21171566	+	.	12	0	5412706_1	26.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=5412706_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:21170008(+)-8:21171566(-)__8_21168001_21193001D;SPAN=1558;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:50 GQ:26 PL:[26.0, 0.0, 95.3] SR:0 DR:12 LR:-26.07 LO:28.28);ALT=G[chr8:21171566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	21835004	+	chr19	10825684	+	.	10	30	5413982_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCTACTCTGGAGGCTGAGGCAGGAGAATC;MAPQ=21;MATEID=5413982_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_8_21829501_21854501_79C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:39 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:30 DR:10 LR:-125.4 LO:125.4);ALT=C[chr19:10825684[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	21922163	+	chr8	21994207	+	.	65	54	5414118_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5414118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_21903001_21928001_87C;SPAN=72044;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:5 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:54 DR:65 LR:-307.0 LO:307.0);ALT=G[chr8:21994207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10309164	+	chr19	10285593	+	.	9	0	10152973_1	8.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=10152973_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10285593(-)-19:10309164(+)__19_10265501_10290501D;SPAN=23571;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:0 DR:9 LR:-8.577 LO:18.05);ALT=]chr19:10309164]T;VARTYPE=BND:DUP-th;JOINTYPE=th
