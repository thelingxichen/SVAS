chr5	130495322	+	chr5	130500854	+	.	18	0	2580428_1	0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2580428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:130495322(+)-5:130500854(-)__5_130487001_130512001D;SPAN=5532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:18 DP:227 GQ:1.9 PL:[0.0, 1.9, 554.5] SR:0 DR:18 LR:2.082 LO:33.0);ALT=G[chr5:130500854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	130498404	+	chr5	130500853	+	.	136	0	2580436_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=2580436_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:130498404(+)-5:130500853(-)__5_130487001_130512001D;SPAN=2449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:136 DP:217 GQ:99 PL:[390.2, 0.0, 136.0] SR:0 DR:136 LR:-396.9 LO:396.9);ALT=T[chr5:130500853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	130599859	+	chr5	130651668	+	.	10	4	2580875_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2580875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_130634001_130659001_91C;SPAN=51809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:26 GQ:29.3 PL:[32.6, 0.0, 29.3] SR:4 DR:10 LR:-32.57 LO:32.57);ALT=G[chr5:130651668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
