chrX	104589118	+	chrX	104595554	+	.	69	61	11337866_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TCTG;MAPQ=60;MATEID=11337866_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_104590501_104615501_211C;SPAN=6436;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:104 DP:9 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:61 DR:69 LR:-307.0 LO:307.0);ALT=G[chrX:104595554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	104778934	+	chrX	104781455	+	AAA	63	46	11338107_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AAA;MAPQ=60;MATEID=11338107_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_104762001_104787001_122C;SPAN=2521;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:18 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:46 DR:63 LR:-254.2 LO:254.2);ALT=A[chrX:104781455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
