chr2	162332271	+	chr2	162334042	+	.	175	120	1465572_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCCA;MAPQ=36;MATEID=1465572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_162312501_162337501_86C;SPAN=1771;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:246 DP:53 GQ:66.4 PL:[729.4, 66.4, 0.0] SR:120 DR:175 LR:-729.5 LO:729.5);ALT=A[chr2:162334042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
