chr4	117166276	-	chr4	117167369	+	.	9	0	2163906_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2163906_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:117166276(-)-4:117167369(-)__4_117159001_117184001D;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:110 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.0927 LO:16.63);ALT=[chr4:117167369[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
