chr4	93568525	+	chr4	93570341	-	.	9	0	2788567_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2788567_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:93568525(+)-4:93570341(+)__4_93565501_93590501D;SPAN=1816;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=T]chr4:93570341];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	93855558	+	chr4	93861562	+	.	29	0	2789213_1	85.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2789213_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:93855558(+)-4:93861562(-)__4_93859501_93884501D;SPAN=6004;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:6 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=T[chr4:93861562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
