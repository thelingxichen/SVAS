chr5	34304798	+	chr5	34307905	+	.	31	31	3357356_1	99.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=ATTTTTTTT;MAPQ=46;MATEID=3357356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_34300001_34325001_86C;SPAN=3107;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:132 GQ:99 PL:[139.4, 0.0, 179.0] SR:31 DR:31 LR:-139.2 LO:139.5);ALT=T[chr5:34307905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
