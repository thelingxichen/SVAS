chr13	108871006	+	chr13	108881546	+	.	8	0	5640565_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5640565_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:108871006(+)-13:108881546(-)__13_108878001_108903001D;SPAN=10540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=G[chr13:108881546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	108922772	+	chr13	108955599	+	TCACTCAAGACTGCTTGCAACTGATTGCAGACAGTGAAACACCAACTATACAAAA	17	21	5640670_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TCACTCAAGACTGCTTGCAACTGATTGCAGACAGTGAAACACCAACTATACAAAA;MAPQ=60;MATEID=5640670_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_108902501_108927501_0C;SPAN=32827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:53 GQ:15.5 PL:[111.2, 0.0, 15.5] SR:21 DR:17 LR:-115.0 LO:115.0);ALT=G[chr13:108955599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	108922772	+	chr13	108939149	+	.	0	35	5640669_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5640669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_108902501_108927501_232C;SPAN=16377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:53 GQ:25.4 PL:[101.3, 0.0, 25.4] SR:35 DR:0 LR:-103.5 LO:103.5);ALT=G[chr13:108939149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	108955953	+	chr13	108959173	+	.	9	59	5641010_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5641010_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_108951501_108976501_71C;SPAN=3220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:115 GQ:97.7 PL:[180.2, 0.0, 97.7] SR:59 DR:9 LR:-181.4 LO:181.4);ALT=G[chr13:108959173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
