chr9	78919501	+	chr9	78922041	+	.	22	0	5897075_1	62.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5897075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:78919501(+)-9:78922041(-)__9_78914501_78939501D;SPAN=2540;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:22 DP:37 GQ:26.3 PL:[62.6, 0.0, 26.3] SR:0 DR:22 LR:-63.36 LO:63.36);ALT=C[chr9:78922041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
