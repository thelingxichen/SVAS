chr5	70751916	+	chr5	70754403	+	.	3	4	2499445_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=2499445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_70731501_70756501_207C;SPAN=2487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:53 GQ:5.6 PL:[5.6, 0.0, 121.1] SR:4 DR:3 LR:-5.447 LO:11.98);ALT=G[chr5:70754403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	71591417	+	chr5	71609908	+	CGTGATATTGTTAAAGAACTAACAGGCAACTTTCTCTCAAATGTTTTATCCATTAAAGATGCAAGATCAG	0	26	2500832_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CGTGATATTGTTAAAGAACTAACAGGCAACTTTCTCTCAAATGTTTTATCCATTAAAGATGCAAGATCAG;MAPQ=60;MATEID=2500832_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_71589001_71614001_229C;SPAN=18491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:49 GQ:46.1 PL:[72.5, 0.0, 46.1] SR:26 DR:0 LR:-72.86 LO:72.86);ALT=C[chr5:71609908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	71591465	+	chr5	71615993	+	.	8	0	2501124_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2501124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:71591465(+)-5:71615993(-)__5_71613501_71638501D;SPAN=24528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:22 GQ:20.6 PL:[20.6, 0.0, 30.5] SR:0 DR:8 LR:-20.45 LO:20.61);ALT=T[chr5:71615993[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	71593578	+	chr5	71615996	+	.	11	0	2501126_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2501126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:71593578(+)-5:71615996(-)__5_71613501_71638501D;SPAN=22418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:23 GQ:23.6 PL:[30.2, 0.0, 23.6] SR:0 DR:11 LR:-30.1 LO:30.1);ALT=T[chr5:71615996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	71610033	+	chr5	71616005	+	.	8	0	2501127_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2501127_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:71610033(+)-5:71616005(-)__5_71613501_71638501D;SPAN=5972;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:30 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.28 LO:19.28);ALT=T[chr5:71616005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
