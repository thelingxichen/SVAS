chrX	191990	+	chr5	99388695	+	.	25	79	10919340_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=10919340_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_171501_196501_399C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:32 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:79 DR:25 LR:-257.5 LO:257.5);ALT=]chrX:191990]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	40872459	+	chrX	569127	-	.	4	37	4159070_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4159070_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_40866001_40891001_57C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:38 DP:31 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:37 DR:4 LR:-112.2 LO:112.2);ALT=A]chrX:569127];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	65278040	+	chr11	65279260	-	.	10	0	6859538_1	0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6859538_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65278040(+)-11:65279260(+)__11_65268001_65293001D;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:160 GQ:10.3 PL:[0.0, 10.3, 409.3] SR:0 DR:10 LR:10.34 LO:17.26);ALT=C]chr11:65279260];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	65290401	-	chrX	2019169	+	.	5	38	6859635_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CATGTTTCTGTGAGCACA;MAPQ=36;MATEID=6859635_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_11_65268001_65293001_0C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:40 DP:95 GQ:99 PL:[106.4, 0.0, 122.9] SR:38 DR:5 LR:-106.3 LO:106.4);ALT=[chrX:2019169[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	65642111	+	chr11	65643520	+	.	0	44	6861773_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTGT;MAPQ=60;MATEID=6861773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_65635501_65660501_240C;SPAN=1409;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:154 GQ:99 PL:[103.7, 0.0, 268.7] SR:44 DR:0 LR:-103.5 LO:107.6);ALT=T[chr11:65643520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65703332	+	chr11	65707195	+	GCG	0	9	6862146_1	0	.	EVDNC=ASSMB;INSERTION=GCG;MAPQ=60;MATEID=6862146_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_65684501_65709501_400C;SPAN=3863;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:167 GQ:15.4 PL:[0.0, 15.4, 435.7] SR:9 DR:0 LR:15.54 LO:14.94);ALT=G[chr11:65707195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	92195	+	chrX	91061	+	.	9	0	10918365_1	0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=10918365_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:91061(-)-23:92195(+)__23_73501_98501D;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:152 GQ:11.2 PL:[0.0, 11.2, 389.4] SR:0 DR:9 LR:11.47 LO:15.32);ALT=]chrX:92195]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	325893	+	chrX	327608	+	.	13	0	10918424_1	0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=10918424_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:325893(+)-23:327608(-)__23_318501_343501D;SPAN=1715;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:13 DP:156 GQ:0.7 PL:[0.7, 0.0, 377.0] SR:0 DR:13 LR:-0.6488 LO:24.13);ALT=A[chrX:327608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	518955	-	chrX	520346	+	.	10	0	10921711_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=10921711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:518955(-)-23:520346(-)__23_514501_539501D;SPAN=1391;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:150 GQ:7.6 PL:[0.0, 7.6, 379.5] SR:0 DR:10 LR:7.629 LO:17.55);ALT=[chrX:520346[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	710355	-	chrX	711561	+	.	9	0	10921164_1	16.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=10921164_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:710355(-)-23:711561(-)__23_686001_711001D;SPAN=1206;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-15.89 LO:19.85);ALT=[chrX:711561[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	741908	+	chrX	740426	+	.	44	0	10921904_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=10921904_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:740426(-)-23:741908(+)__23_735001_760001D;SPAN=1482;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:44 DP:91 GQ:97.7 PL:[120.8, 0.0, 97.7] SR:0 DR:44 LR:-120.7 LO:120.7);ALT=]chrX:741908]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	766724	-	chrX	767857	+	.	10	0	10921375_1	0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=10921375_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:766724(-)-23:767857(-)__23_759501_784501D;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:183 GQ:16.3 PL:[0.0, 16.3, 475.3] SR:0 DR:10 LR:16.57 LO:16.67);ALT=[chrX:767857[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	802863	+	chrX	804142	-	.	9	0	10921273_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=10921273_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:802863(+)-23:804142(+)__23_784001_809001D;SPAN=1279;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:139 GQ:7.8 PL:[0.0, 7.8, 353.1] SR:0 DR:9 LR:7.95 LO:15.68);ALT=T]chrX:804142];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	1044379	+	chrX	1107283	+	.	22	41	10923505_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=TAGGGTTGTGACCCAG;MAPQ=13;MATEID=10923505_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_23_1029001_1054001_46C;SPAN=62904;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:57 DP:15 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:41 DR:22 LR:-168.3 LO:168.3);ALT=G[chrX:1107283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1450155	+	chrX	1453316	+	.	6	26	10924955_1	60.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=TACTCGGGAGGCTGAGGCAGGAGAATC;MAPQ=42;MATEID=10924955_2;MATENM=0;NM=7;NUMPARTS=2;SCTG=c_23_1445501_1470501_45C;SPAN=3161;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:30 DP:143 GQ:60.5 PL:[60.5, 0.0, 284.9] SR:26 DR:6 LR:-60.29 LO:68.7);ALT=C[chrX:1453316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1756051	+	chrX	1760254	+	.	10	0	10927120_1	8.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=10927120_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1756051(+)-23:1760254(-)__23_1739501_1764501D;SPAN=4203;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:0 DR:10 LR:-8.085 LO:19.77);ALT=C[chrX:1760254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	1938903	+	chrX	1937760	+	.	50	0	10928873_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=10928873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:1937760(-)-23:1938903(+)__23_1935501_1960501D;SPAN=1143;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:50 DP:95 GQ:89.9 PL:[139.4, 0.0, 89.9] SR:0 DR:50 LR:-139.8 LO:139.8);ALT=]chrX:1938903]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	2195519	+	chrX	2200337	+	.	34	1	10929850_1	69.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=GAGAGAGATGGAGAGGGAACAGGGAGAGAGAGGGAGGGCAAAC;MAPQ=0;MATEID=10929850_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_2180501_2205501_229C;SECONDARY;SPAN=4818;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:172 GQ:69.2 PL:[69.2, 0.0, 346.4] SR:1 DR:34 LR:-68.94 LO:79.62);ALT=C[chrX:2200337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	2242782	+	chrX	2468198	-	.	11	0	10931595_1	14.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=10931595_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:2242782(+)-23:2468198(+)__23_2450001_2475001D;SPAN=225416;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:0 DR:11 LR:-13.82 LO:22.76);ALT=G]chrX:2468198];VARTYPE=BND:INV-hh;JOINTYPE=hh
