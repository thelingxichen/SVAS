chr11	123841181	+	chr11	123843930	-	.	2	4	7247108_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATAAAAACTCTCAA;MAPQ=60;MATEID=7247108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_123823001_123848001_310C;SPAN=2749;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:4 DP:192 GQ:38.5 PL:[0.0, 38.5, 541.3] SR:4 DR:2 LR:38.81 LO:4.981);ALT=T]chr11:123843930];VARTYPE=BND:INV-hh;JOINTYPE=hh
