chr12	121875519	+	chr12	120534913	+	.	10	6	7871482_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=7871482_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121863001_121888001_346C;SPAN=1340606;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:6 DR:10 LR:-32.72 LO:35.42);ALT=]chr12:121875519]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	120772163	+	chr12	120566061	+	AAGTGC	9	8	7865151_1	26.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=AAGTGC;MAPQ=60;MATEID=7865151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120760501_120785501_405C;SPAN=206102;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:12 DP:50 GQ:26 PL:[26.0, 0.0, 95.3] SR:8 DR:9 LR:-26.07 LO:28.28);ALT=]chr12:120772163]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	30711670	+	chr12	120742612	+	.	3	35	10475291_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATATATAT;MAPQ=60;MATEID=10475291_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30698501_30723501_558C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:37 DP:32 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:35 DR:3 LR:-108.9 LO:108.9);ALT=]chr20:30711670]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	122094517	-	chr12	122095682	+	.	4	2	7872852_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCAAGCGATTCT;MAPQ=60;MATEID=7872852_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122083501_122108501_141C;SPAN=1165;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:5 DP:152 GQ:24.4 PL:[0.0, 24.4, 415.9] SR:2 DR:4 LR:24.68 LO:7.216);ALT=[chr12:122095682[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	122471296	-	chr12	122472430	+	.	10	0	7875186_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7875186_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:122471296(-)-12:122472430(-)__12_122451001_122476001D;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:147 GQ:6.6 PL:[0.0, 6.6, 369.6] SR:0 DR:10 LR:6.816 LO:17.64);ALT=[chr12:122472430[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	29810864	+	chr20	29804531	+	.	9	0	10468126_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=10468126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:29804531(-)-20:29810864(+)__20_29792001_29817001D;SPAN=6333;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:271 GQ:43.3 PL:[0.0, 43.3, 742.6] SR:0 DR:9 LR:43.71 LO:13.03);ALT=]chr20:29810864]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	30199849	-	chr20	30325274	+	TA	47	24	10472253_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TA;MAPQ=60;MATEID=10472253_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30306501_30331501_133C;SPAN=125425;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:64 DP:125 GQ:99 PL:[177.5, 0.0, 124.7] SR:24 DR:47 LR:-177.9 LO:177.9);ALT=[chr20:30325274[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	30322130	+	chr20	30329757	-	.	9	53	10472425_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=10472425_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30306501_30331501_262C;SPAN=7627;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:54 DP:191 GQ:99 PL:[126.8, 0.0, 334.7] SR:53 DR:9 LR:-126.5 LO:131.8);ALT=T]chr20:30329757];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	31049372	+	chr20	31050645	-	.	8	0	10477743_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=10477743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31049372(+)-20:31050645(+)__20_31041501_31066501D;SPAN=1273;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:141 GQ:11.4 PL:[0.0, 11.4, 363.0] SR:0 DR:8 LR:11.79 LO:13.47);ALT=C]chr20:31050645];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	31310881	+	chr20	31312779	+	.	48	30	10480640_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AAAGACTTGTG;MAPQ=35;MATEID=10480640_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_31311001_31336001_1C;SPAN=1898;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:37 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:30 DR:48 LR:-201.3 LO:201.3);ALT=G[chr20:31312779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
