chr2	132670950	+	chrX	102408249	-	.	5	9	998922_1	46.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=AGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAAG;MAPQ=48;MATEID=998922_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_2_132667501_132692501_72C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:16 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:9 DR:5 LR:-45.42 LO:45.42);ALT=T]chrX:102408249];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	133001427	-	chr14	19000146	+	.	28	0	5657600_1	75.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5657600_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:133001427(-)-14:19000146(-)__14_18987501_19012501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:63 GQ:75.5 PL:[75.5, 0.0, 75.5] SR:0 DR:28 LR:-75.36 LO:75.36);ALT=[chr14:19000146[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	133027308	+	chr2	133024059	+	.	10	0	1000784_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=1000784_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:133024059(-)-2:133027308(+)__2_133010501_133035501D;SPAN=3249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:148 GQ:6.9 PL:[0.0, 6.9, 372.9] SR:0 DR:10 LR:7.087 LO:17.61);ALT=]chr2:133027308]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	102508981	+	chrX	102510004	+	.	30	0	7487002_1	86.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7487002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:102508981(+)-23:102510004(-)__23_102508001_102533001D;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:47 GQ:26.9 PL:[86.3, 0.0, 26.9] SR:0 DR:30 LR:-87.95 LO:87.95);ALT=G[chrX:102510004[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	102931979	+	chrX	102940097	+	ACAATCTTCCTTCTTTCCCTTCCAAGAACTCCTAGTGATTTCCCAGATGAAATCTTATAGATCTTCTGGGATGGTCTAGAAGGGTGAAGTGGGAGATACA	0	18	7487688_1	44.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=ACAATCTTCCTTCTTTCCCTTCCAAGAACTCCTAGTGATTTCCCAGATGAAATCTTATAGATCTTCTGGGATGGTCTAGAAGGGTGAAGTGGGAGATACA;MAPQ=60;MATEID=7487688_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_102924501_102949501_207C;SPAN=8118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:57 GQ:44 PL:[44.0, 0.0, 93.5] SR:18 DR:0 LR:-43.98 LO:44.99);ALT=A[chrX:102940097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	102931979	+	chrX	102933427	+	.	0	10	7487687_1	20.0	.	DISC_MAPQ=255;EVDNC=TSI_L;MAPQ=60;MATEID=7487687_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_102924501_102949501_207C;SPAN=1448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:10 DR:0 LR:-20.01 LO:22.86);ALT=A[chrX:102933427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	102933590	+	chrX	102941564	+	.	12	0	7487693_1	25.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7487693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:102933590(+)-23:102941564(-)__23_102924501_102949501D;SPAN=7974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=G[chrX:102941564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	103375920	+	chrX	103401594	+	.	8	0	7488376_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7488376_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:103375920(+)-23:103401594(-)__23_103390001_103415001D;SPAN=25674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=G[chrX:103401594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
