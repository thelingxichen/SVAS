chrX	78619097	+	chrX	78622697	+	.	20	0	7457199_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7457199_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:78619097(+)-23:78622697(-)__23_78620501_78645501D;SPAN=3600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:38 GQ:35.9 PL:[55.7, 0.0, 35.9] SR:0 DR:20 LR:-55.94 LO:55.94);ALT=T[chrX:78622697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	78946448	+	chrX	78948837	+	T	57	24	7457688_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TTCCTCTTCT;INSERTION=T;MAPQ=60;MATEID=7457688_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_23_78939001_78964001_200C;SPAN=2389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:13 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:24 DR:57 LR:-194.7 LO:194.7);ALT=T[chrX:78948837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
