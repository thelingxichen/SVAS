chr2	139569396	+	chr3	44742593	-	.	4	17	1982732_1	45.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTTCCTTCCTTCCTTCCTTCCT;MAPQ=60;MATEID=1982732_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_62C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:18 DP:52 GQ:45.5 PL:[45.5, 0.0, 78.5] SR:17 DR:4 LR:-45.33 LO:45.88);ALT=T]chr3:44742593];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	241012418	+	chr3	45344935	-	GCTCTGTCACCAGGCTGGAGTGCAGTGGTACGATCC	8	75	1785137_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=GCTCTGTCACCAGGCTGGAGTGCAGTGGTACGATCC;MAPQ=60;MATEID=1785137_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_2_241006501_241031501_349C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:81 DP:51 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:75 DR:8 LR:-237.7 LO:237.7);ALT=C]chr3:45344935];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	241012441	-	chr3	45344858	+	GCCACCACCACGCCCAGCTAATTTTTTGCATTTTAGTAT	4	66	1785142_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;INSERTION=GCCACCACCACGCCCAGCTAATTTTTTGCATTTTAGTAT;MAPQ=60;MATEID=1785142_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_2_241006501_241031501_349C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:69 DP:53 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:66 DR:4 LR:-204.7 LO:204.7);ALT=[chr3:45344858[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	241097563	+	chr2	241098579	+	.	14	0	1785451_1	24.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=1785451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:241097563(+)-2:241098579(-)__2_241080001_241105001D;SPAN=1016;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:82 GQ:24.2 PL:[24.2, 0.0, 172.7] SR:0 DR:14 LR:-24.0 LO:30.65);ALT=T[chr2:241098579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	44585058	+	chr3	44412869	+	.	83	29	1981168_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=1981168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44565501_44590501_141C;SPAN=172189;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:106 DP:74 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:29 DR:83 LR:-313.6 LO:313.6);ALT=]chr3:44585058]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	44740991	-	chr3	44742263	+	.	99	72	1982760_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=TCCCAAAGTGCTGGGATTACAGG;MAPQ=60;MATEID=1982760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_303C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:161 DP:127 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:72 DR:99 LR:-475.3 LO:475.3);ALT=[chr3:44742263[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
