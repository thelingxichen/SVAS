chr11	60754438	+	chr11	60758281	+	TATATATATATATAATTTATATATAAATTTATATAAATTGGACCC	27	79	6836020_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;INSERTION=TATATATATATATAATTTATATATAAATTTATATAAATTGGACCC;MAPQ=10;MATEID=6836020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_60735501_60760501_239C;SPAN=3843;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:107 GQ:18.9 PL:[297.0, 18.9, 0.0] SR:79 DR:27 LR:-300.7 LO:300.7);ALT=A[chr11:60758281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61843628	+	chr11	61731233	+	.	77	27	6841445_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6841445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61838001_61863001_499C;SPAN=112395;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:97 DP:65 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:27 DR:77 LR:-287.2 LO:287.2);ALT=]chr11:61843628]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	61841813	+	chr14	81786774	+	C	33	47	6841489_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=6841489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61838001_61863001_496C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:68 DP:118 GQ:93.5 PL:[192.5, 0.0, 93.5] SR:47 DR:33 LR:-194.3 LO:194.3);ALT=G[chr14:81786774[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr14	81269554	+	chr14	81222756	+	.	68	45	8635552_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=8635552_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_81266501_81291501_126C;SPAN=46798;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:88 DP:57 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:45 DR:68 LR:-260.8 LO:260.8);ALT=]chr14:81269554]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	81878211	+	chr14	81880613	+	TGCTTATCTTAACTCTG	58	75	8637654_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=CTATCTGG;INSERTION=TGCTTATCTTAACTCTG;MAPQ=60;MATEID=8637654_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_14_81854501_81879501_303C;SPAN=2402;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:113 DP:41 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:75 DR:58 LR:-333.4 LO:333.4);ALT=G[chr14:81880613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	82499110	+	chr14	82503331	+	AACATAAATC	58	48	8640208_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AACATAAATC;MAPQ=60;MATEID=8640208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_82491501_82516501_29C;SPAN=4221;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:80 GQ:24 PL:[264.0, 24.0, 0.0] SR:48 DR:58 LR:-264.1 LO:264.1);ALT=T[chr14:82503331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
