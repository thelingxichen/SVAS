chr15	26872523	+	chr1	204151126	+	.	3	36	765789_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=TTTATT;MAPQ=60;MATEID=765789_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_204134001_204159001_30C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:36 DP:55 GQ:28.1 PL:[104.0, 0.0, 28.1] SR:36 DR:3 LR:-106.2 LO:106.2);ALT=]chr15:26872523]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	57775044	+	chr2	57773380	+	.	8	0	1019822_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1019822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:57773380(-)-2:57775044(+)__2_57771001_57796001D;SPAN=1664;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=]chr2:57775044]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	58234476	-	chr2	58235527	+	.	10	0	1021572_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1021572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:58234476(-)-2:58235527(-)__2_58212001_58237001D;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:158 GQ:9.7 PL:[0.0, 9.7, 402.6] SR:0 DR:10 LR:9.796 LO:17.32);ALT=[chr2:58235527[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	59108044	+	chr10	8604000	-	.	8	0	6076896_1	12.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6076896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:59108044(+)-10:8604000(+)__10_8599501_8624501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=C]chr10:8604000];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	90317662	-	chr10	8595388	+	.	57	54	6076273_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AAGCTCTCT;MAPQ=60;MATEID=6076273_2;MATENM=3;NM=0;NUMPARTS=3;SCTG=c_10_8575001_8600001_241C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:36 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:54 DR:57 LR:-270.7 LO:270.7);ALT=[chr10:8595388[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	90545003	+	chr8	90553464	+	.	36	39	5534974_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=20;MATEID=5534974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_90527501_90552501_190C;SPAN=8461;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:66 DP:50 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:39 DR:36 LR:-194.7 LO:194.7);ALT=A[chr8:90553464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	91422350	-	chr15	27718778	+	.	10	0	8802579_1	0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=8802579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_27709501_27734501_9C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:337 GQ:58.1 PL:[0.0, 58.1, 934.1] SR:0 DR:10 LR:58.29 LO:13.98);ALT=[chr15:27718778[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
