chr11	107151543	-	chr11	107169657	+	.	20	0	7171619_1	59.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=7171619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:107151543(-)-11:107169657(-)__11_107163001_107188001D;SPAN=18114;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:20 DP:5 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:20 LR:-59.41 LO:59.41);ALT=[chr11:107169657[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
