chr16	53243725	+	chr16	53256555	+	.	3	14	6213916_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6213916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_53238501_53263501_145C;SPAN=12830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:44 GQ:41 PL:[41.0, 0.0, 64.1] SR:14 DR:3 LR:-40.9 LO:41.22);ALT=G[chr16:53256555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	53515747	+	chr16	53524040	+	.	5	3	6214441_1	7.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6214441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_53508001_53533001_292C;SPAN=8293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:45 GQ:7.7 PL:[7.7, 0.0, 100.1] SR:3 DR:5 LR:-7.614 LO:12.43);ALT=G[chr16:53524040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
