chr1	26291455	+	chr1	27550413	+	.	59	26	141165_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=141165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27538001_27563001_109C;SPAN=1258958;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:75 DP:44 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:26 DR:59 LR:-221.2 LO:221.2);ALT=A[chr1:27550413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27072358	+	chr1	26890603	+	.	44	37	139279_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=AAC;MAPQ=60;MATEID=139279_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_27048001_27073001_58C;SPAN=181755;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:47 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:37 DR:44 LR:-208.0 LO:208.0);ALT=]chr1:27072358]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	69772314	+	chr1	27157317	+	TGCTCTGTCGCCC	7	75	9393483_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=TGCTCTGTCGCCC;MAPQ=60;MATEID=9393483_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_16_69751501_69776501_255C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:80 DP:30 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:75 DR:7 LR:-237.7 LO:237.7);ALT=]chr16:69772314]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	69854331	+	chr16	69858806	+	T	89	102	9392948_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=9392948_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69849501_69874501_471C;SPAN=4475;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:163 DP:103 GQ:43.9 PL:[481.9, 43.9, 0.0] SR:102 DR:89 LR:-481.9 LO:481.9);ALT=G[chr16:69858806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69859021	+	chr16	69854686	+	CAAAAGTGAACA	129	95	9392949_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CAAAAGTGAACA;MAPQ=60;MATEID=9392949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69849501_69874501_360C;SPAN=4335;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:187 DP:140 GQ:50.5 PL:[554.5, 50.5, 0.0] SR:95 DR:129 LR:-554.5 LO:554.5);ALT=]chr16:69859021]A;VARTYPE=BND:DUP-th;JOINTYPE=th
