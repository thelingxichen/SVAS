chr1	205687610	+	chr1	205688655	+	.	32	22	509544_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=509544_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_205677501_205702501_198C;SPAN=1045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:101 GQ:91.7 PL:[151.1, 0.0, 91.7] SR:22 DR:32 LR:-151.6 LO:151.6);ALT=G[chr1:205688655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	205689785	+	chr1	205719085	+	TGAGTGAGAATCATCCTTCTTGGTCTTCACATCTTTGTCTTCTGAGTCCTCACTATCTTCCTGTGAATTCTTTCCAGATCGCCTCTTATTTTTAGCTTCTCGGGGAGATGATCGAATTTTCTTAGTGGGAGGGCCCGAATCTCTTCCATAATCTTCATCTGCATCATCAGATTCCTGAAACTGTGAGTAATCAACAACCTTCCTATTT	2	88	509552_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TGAGTGAGAATCATCCTTCTTGGTCTTCACATCTTTGTCTTCTGAGTCCTCACTATCTTCCTGTGAATTCTTTCCAGATCGCCTCTTATTTTTAGCTTCTCGGGGAGATGATCGAATTTTCTTAGTGGGAGGGCCCGAATCTCTTCCATAATCTTCATCTGCATCATCAGATTCCTGAAACTGTGAGTAATCAACAACCTTCCTATTT;MAPQ=60;MATEID=509552_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_1_205677501_205702501_83C;SPAN=29300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:60 GQ:24 PL:[264.0, 24.0, 0.0] SR:88 DR:2 LR:-264.1 LO:264.1);ALT=C[chr1:205719085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	205689808	+	chr1	205696827	+	.	8	0	509553_1	2.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=509553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:205689808(+)-1:205696827(-)__1_205677501_205702501D;SPAN=7019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=A[chr1:205696827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	205696969	+	chr1	205719084	+	.	16	0	509822_1	33.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=509822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:205696969(+)-1:205719084(-)__1_205702001_205727001D;SPAN=22115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:70 GQ:33.8 PL:[33.8, 0.0, 136.1] SR:0 DR:16 LR:-33.85 LO:37.32);ALT=T[chr1:205719084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	205698803	+	chr1	205719245	+	.	19	0	509824_1	46.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=509824_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:205698803(+)-1:205719245(-)__1_205702001_205727001D;SPAN=20442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:62 GQ:46.1 PL:[46.1, 0.0, 102.2] SR:0 DR:19 LR:-45.92 LO:47.18);ALT=G[chr1:205719245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206288352	+	chr1	206289366	+	.	3	37	511650_1	74.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=511650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_206265501_206290501_457C;SPAN=1014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:200 GQ:74.5 PL:[74.5, 0.0, 411.2] SR:37 DR:3 LR:-74.55 LO:87.9);ALT=G[chr1:206289366[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206288402	+	chr1	206306066	+	.	32	0	511651_1	77.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=511651_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:206288402(+)-1:206306066(-)__1_206265501_206290501D;SPAN=17664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:104 GQ:77.6 PL:[77.6, 0.0, 173.3] SR:0 DR:32 LR:-77.46 LO:79.53);ALT=A[chr1:206306066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206289682	+	chr1	206306066	+	.	111	0	511660_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=511660_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:206289682(+)-1:206306066(-)__1_206265501_206290501D;SPAN=16384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:60 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:111 LR:-326.8 LO:326.8);ALT=C[chr1:206306066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206299832	+	chr1	206306067	+	.	18	0	511497_1	16.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=511497_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:206299832(+)-1:206306067(-)__1_206290001_206315001D;SPAN=6235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:158 GQ:16.6 PL:[16.6, 0.0, 366.5] SR:0 DR:18 LR:-16.61 LO:35.98);ALT=G[chr1:206306067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206644041	+	chr1	206646538	+	CTCAGCTCCTGGACGTGCCACAGACAGAAAGCATAACATACACTCGCCAGGAAGAGCCTTTGCCTGACTCAGGGCAGCTCAGAGTGTGG	0	10	512574_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=CTCAGCTCCTGGACGTGCCACAGACAGAAAGCATAACATACACTCGCCAGGAAGAGCCTTTGCCTGACTCAGGGCAGCTCAGAGTGTGG;MAPQ=60;MATEID=512574_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_206633001_206658001_20C;SPAN=2497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:10 DR:0 LR:-7.814 LO:19.72);ALT=G[chr1:206646538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	206765178	+	chr1	206766968	+	.	0	19	512944_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=512944_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_206755501_206780501_162C;SPAN=1790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:125 GQ:29 PL:[29.0, 0.0, 273.2] SR:19 DR:0 LR:-28.85 LO:40.55);ALT=C[chr1:206766968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	207542035	+	chr1	207545565	+	.	96	4	515527_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCAACATTCACTTTTGAAAGGGCCATGGAGGAAAATGAACCAGGAAGATCCTCCCTGGGGCAGAGCTACCAC;MAPQ=60;MATEID=515527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_207539501_207564501_272C;SPAN=3530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:8 GQ:27 PL:[297.0, 27.0, 0.0] SR:4 DR:96 LR:-297.1 LO:297.1);ALT=C[chr1:207545565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	207925654	+	chr1	207930358	+	.	6	9	516886_1	7.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=516886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_207907001_207932001_163C;SPAN=4704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:107 GQ:7.4 PL:[7.4, 0.0, 251.6] SR:9 DR:6 LR:-7.322 LO:21.47);ALT=G[chr1:207930358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	207981233	+	chr1	208014818	+	.	15	14	517068_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GAGG;MAPQ=60;MATEID=517068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_208005001_208030001_84C;SPAN=33585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:35 GQ:13.7 PL:[69.8, 0.0, 13.7] SR:14 DR:15 LR:-71.71 LO:71.71);ALT=G[chr1:208014818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	208072617	+	chr1	208084365	+	.	11	0	517299_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=517299_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:208072617(+)-1:208084365(-)__1_208078501_208103501D;SPAN=11748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:0 DR:11 LR:-23.31 LO:25.67);ALT=A[chr1:208084365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	208073348	+	chr1	208084347	+	.	87	26	517300_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=517300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_208078501_208103501_101C;SPAN=10999;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:50 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:26 DR:87 LR:-287.2 LO:287.2);ALT=G[chr1:208084347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
