chr13	72807622	+	chr13	72812359	+	ATATA	64	63	5549486_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=ATATA;MAPQ=60;MATEID=5549486_2;MATENM=2;NM=3;NUMPARTS=2;SCTG=c_13_72789501_72814501_13C;SPAN=4737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:27 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:63 DR:64 LR:-290.5 LO:290.5);ALT=C[chr13:72812359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	72843037	+	chr13	72846925	+	AAATTGCAG	26	25	5549623_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;INSERTION=AAATTGCAG;MAPQ=22;MATEID=5549623_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_13_72838501_72863501_232C;SPAN=3888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:52 GQ:2.6 PL:[121.4, 0.0, 2.6] SR:25 DR:26 LR:-127.7 LO:127.7);ALT=T[chr13:72846925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	73284485	+	chr13	73293089	+	.	0	21	5550880_1	46.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5550880_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_73279501_73304501_347C;SPAN=8604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:85 GQ:46.4 PL:[46.4, 0.0, 158.6] SR:21 DR:0 LR:-46.29 LO:49.8);ALT=T[chr13:73293089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	73293236	+	chr13	73301662	+	.	19	6	5550909_1	55.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5550909_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_73279501_73304501_296C;SPAN=8426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:77 GQ:55.1 PL:[55.1, 0.0, 131.0] SR:6 DR:19 LR:-55.06 LO:56.8);ALT=C[chr13:73301662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
