chr21	37529241	+	chr21	37537005	+	.	7	3	7170183_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7170183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_37534001_37559001_117C;SPAN=7764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:3 DR:7 LR:-16.11 LO:18.33);ALT=G[chr21:37537005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	37692650	+	chr21	37709169	+	.	12	0	7170909_1	30.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7170909_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:37692650(+)-21:37709169(-)__21_37681001_37706001D;SPAN=16519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:0 DR:12 LR:-30.67 LO:30.91);ALT=G[chr21:37709169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	37706016	+	chr21	37709170	+	.	0	9	7170709_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7170709_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_37705501_37730501_158C;SPAN=3154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:9 DR:0 LR:-9.39 LO:18.21);ALT=G[chr21:37709170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	38439680	+	chr21	38441852	+	.	0	21	7173073_1	57.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7173073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_38440501_38465501_149C;SPAN=2172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:45 GQ:50.6 PL:[57.2, 0.0, 50.6] SR:21 DR:0 LR:-57.14 LO:57.14);ALT=T[chr21:38441852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	38441924	+	chr21	38444734	+	.	0	17	7173082_1	37.0	.	EVDNC=ASSMB;MAPQ=45;MATEID=7173082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_38440501_38465501_175C;SPAN=2810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:68 GQ:37.7 PL:[37.7, 0.0, 126.8] SR:17 DR:0 LR:-37.69 LO:40.42);ALT=A[chr21:38444734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	38536517	+	chr21	38537852	+	.	2	8	7173300_1	12.0	.	DISC_MAPQ=41;EVDNC=ASDIS;MAPQ=60;MATEID=7173300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_38514001_38539001_75C;SPAN=1335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:76 GQ:12.5 PL:[12.5, 0.0, 170.9] SR:8 DR:2 LR:-12.42 LO:20.66);ALT=A[chr21:38537852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	38634241	+	chr21	38639574	+	.	8	0	7173783_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7173783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:38634241(+)-21:38639574(-)__21_38636501_38661501D;SPAN=5333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=A[chr21:38639574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
