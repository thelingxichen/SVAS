chr12	17707806	-	chr13	69485718	+	.	10	79	7436454_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATATATATATATATACATATATATA;MAPQ=60;MATEID=7436454_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_17689001_17714001_55C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:80 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:79 DR:10 LR:-247.6 LO:247.6);ALT=[chr13:69485718[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr13	68811522	+	chr13	68931387	+	.	49	29	8132939_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8132939_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_68918501_68943501_276C;SPAN=119865;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:65 DP:35 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:29 DR:49 LR:-191.4 LO:191.4);ALT=T[chr13:68931387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	68945754	+	chr13	68952611	+	.	56	51	8132995_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=8132995_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_68943001_68968001_224C;SPAN=6857;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:86 DP:84 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:51 DR:56 LR:-254.2 LO:254.2);ALT=T[chr13:68952611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
