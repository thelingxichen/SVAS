chr5	72794363	+	chr5	72798311	+	.	54	0	2502870_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2502870_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:72794363(+)-5:72798311(-)__5_72789501_72814501D;SPAN=3948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:131 GQ:99 PL:[143.0, 0.0, 172.7] SR:0 DR:54 LR:-142.8 LO:142.9);ALT=C[chr5:72798311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	72794363	+	chr5	72798738	+	.	10	0	2502871_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2502871_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:72794363(+)-5:72798738(-)__5_72789501_72814501D;SPAN=4375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:101 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.647 LO:19.35);ALT=C[chr5:72798738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	72798974	+	chr5	72801036	+	.	8	0	2502884_1	0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2502884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:72798974(+)-5:72801036(-)__5_72789501_72814501D;SPAN=2062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:130 GQ:8.7 PL:[0.0, 8.7, 333.3] SR:0 DR:8 LR:8.812 LO:13.76);ALT=A[chr5:72801036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
