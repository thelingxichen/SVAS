chr16	32517916	+	chr16	32520797	+	.	99	70	9277190_1	99.0	.	DISC_MAPQ=15;EVDNC=ASDIS;HOMSEQ=GTGTTTCCAAATTGCTGAA;MAPQ=29;MATEID=9277190_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_32511501_32536501_434C;SPAN=2881;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:138 DP:44 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:70 DR:99 LR:-409.3 LO:409.3);ALT=A[chr16:32520797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	33075552	+	chr16	33074343	+	.	11	0	9281763_1	18.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=9281763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:33074343(-)-16:33075552(+)__16_33050501_33075501D;SPAN=1209;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:0 DR:11 LR:-18.7 LO:24.04);ALT=]chr16:33075552]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	33899045	+	chr16	33897814	+	.	28	0	9289186_1	0	.	DISC_MAPQ=44;EVDNC=TSI_L;HOMSEQ=ATTCCATT;MAPQ=22;MATEID=9289186_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCTTACCTTA;SCTG=c_16_33883501_33908501_104C;SPAN=1231;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:28 DP:255 GQ:28 PL:[0.0, 28.0, 221.2] SR:0 DR:28 LR:32.66 LO:2.743);ALT=]chr16:33899045]A;VARTYPE=BND:DUP-th;JOINTYPE=th
