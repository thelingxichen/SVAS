chr3	18433452	+	chr3	18054231	+	.	64	30	1872416_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GAA;MAPQ=60;MATEID=1872416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_18424001_18449001_300C;SPAN=379221;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:78 DP:83 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:30 DR:64 LR:-244.3 LO:244.3);ALT=]chr3:18433452]G;VARTYPE=BND:DUP-th;JOINTYPE=th
