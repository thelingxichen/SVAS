chr7	2290350	-	chr7	3094712	+	.	35	0	4498279_1	94.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4498279_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2290350(-)-7:3094712(-)__7_2278501_2303501D;SPAN=804362;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:78 GQ:94.4 PL:[94.4, 0.0, 94.4] SR:0 DR:35 LR:-94.4 LO:94.4);ALT=[chr7:3094712[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
