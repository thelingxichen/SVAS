chr4	47458748	+	chr4	47462161	+	.	0	14	1957408_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1957408_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_47456501_47481501_268C;SPAN=3413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:14 DR:0 LR:-28.06 LO:32.03);ALT=T[chr4:47462161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	47458796	+	chr4	47465602	+	.	12	0	1957409_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1957409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:47458796(+)-4:47465602(-)__4_47456501_47481501D;SPAN=6806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:0 DR:12 LR:-20.92 LO:26.38);ALT=A[chr4:47465602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	47462318	+	chr4	47465603	+	.	29	4	1957413_1	88.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1957413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_47456501_47481501_246C;SPAN=3285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:53 GQ:38.6 PL:[88.1, 0.0, 38.6] SR:4 DR:29 LR:-88.92 LO:88.92);ALT=T[chr4:47465603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
