chr2	202146658	+	chr2	202149441	+	.	129	31	1623365_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TCAAATTCTT;MAPQ=60;MATEID=1623365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_202149501_202174501_204C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:151 DP:14 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:31 DR:129 LR:-445.6 LO:445.6);ALT=T[chr2:202149441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
