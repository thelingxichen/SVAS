chr6	170380346	+	chr6	170381487	+	CCCCATCCCTCCATCCACCCCCATCCCTCCATCCATCCC	2	51	4487179_1	99.0	.	DISC_MAPQ=4;EVDNC=TSI_G;HOMSEQ=ATCCACCCCCATCCCTCCATCCACCCCCATCCCTCCAT;INSERTION=CCCCATCCCTCCATCCACCCCCATCCCTCCATCCATCCC;MAPQ=25;MATEID=4487179_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_6_170373001_170398001_193C;SECONDARY;SPAN=1141;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:53 DP:89 GQ:65 PL:[150.8, 0.0, 65.0] SR:51 DR:2 LR:-152.7 LO:152.7);ALT=C[chr6:170381487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
