chr18	75266998	+	chr18	75268160	+	.	137	113	10085023_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=10085023_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_75264001_75289001_255C;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:205 DP:41 GQ:55.3 PL:[607.3, 55.3, 0.0] SR:113 DR:137 LR:-607.3 LO:607.3);ALT=T[chr18:75268160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
