chr3	105794689	+	chrX	26922374	-	G	5	32	2219027_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;INSERTION=G;MAPQ=15;MATEID=2219027_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_105791001_105816001_245C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:35 DP:36 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:32 DR:5 LR:-105.6 LO:105.6);ALT=G]chrX:26922374];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	141379669	+	chr3	105828863	+	.	50	40	3805332_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=4;MATEID=3805332_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_5_141365001_141390001_45C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:39 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:40 DR:50 LR:-217.9 LO:217.9);ALT=]chr5:141379669]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	105831609	+	chr9	107606637	-	.	29	0	5952209_1	85.0	.	DISC_MAPQ=6;EVDNC=DSCRD;IMPRECISE;MAPQ=6;MATEID=5952209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:105831609(+)-9:107606637(+)__9_107604001_107629001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:27 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=G]chr9:107606637];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	141579321	+	chr5	141011684	+	.	16	0	3806225_1	41.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=3806225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:141011684(-)-5:141579321(+)__5_141561001_141586001D;SPAN=567637;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:16 DP:40 GQ:41.9 PL:[41.9, 0.0, 55.1] SR:0 DR:16 LR:-41.98 LO:42.08);ALT=]chr5:141579321]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	107362893	+	chr9	107369025	+	.	27	0	5951435_1	79.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5951435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:107362893(+)-9:107369025(-)__9_107359001_107384001D;SPAN=6132;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:27 DP:36 GQ:6.8 PL:[79.4, 0.0, 6.8] SR:0 DR:27 LR:-82.78 LO:82.78);ALT=C[chr9:107369025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	107369441	+	chr9	107363217	+	.	38	22	5951437_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCTAATTTCTTGAAATAAGAAGAAAAATTCTTATTTCCTCCT;MAPQ=60;MATEID=5951437_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_9_107359001_107384001_195C;SPAN=6224;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:54 DP:41 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:22 DR:38 LR:-158.4 LO:158.4);ALT=]chr9:107369441]T;VARTYPE=BND:DUP-th;JOINTYPE=th
