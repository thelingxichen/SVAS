chr2	108275311	+	chr2	108279109	+	.	56	49	1236188_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1236188_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_108265501_108290501_317C;SPAN=3798;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:70 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:49 DR:56 LR:-267.4 LO:267.4);ALT=A[chr2:108279109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
