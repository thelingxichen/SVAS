chr1	218182502	+	chr1	218188595	+	.	0	71	826134_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TATTTTGACTTCTT;MAPQ=60;MATEID=826134_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_218172501_218197501_198C;SPAN=6093;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:71 DP:38 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:71 DR:0 LR:-208.0 LO:208.0);ALT=T[chr1:218188595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
