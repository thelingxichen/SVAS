chr18	64959014	+	chr18	64967262	+	.	79	60	10047262_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=10047262_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_18_64949501_64974501_19C;SPAN=8248;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:118 DP:22 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:60 DR:79 LR:-349.9 LO:349.9);ALT=C[chr18:64967262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	65038232	+	chr18	65598803	+	.	17	0	10048609_1	49.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=10048609_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:65038232(+)-18:65598803(-)__18_65586501_65611501D;SPAN=560571;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:17 DP:12 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:17 LR:-49.51 LO:49.51);ALT=C[chr18:65598803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
