chr6	23743259	+	chr6	23745946	+	.	49	49	2744835_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=2744835_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_6_23740501_23765501_206C;SPAN=2687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:66 GQ:21 PL:[231.0, 21.0, 0.0] SR:49 DR:49 LR:-231.1 LO:231.1);ALT=T[chr6:23745946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24325366	+	chr6	24327808	+	.	61	39	2746771_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TCTCC;MAPQ=60;MATEID=2746771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24304001_24329001_354C;SPAN=2442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:56 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:39 DR:61 LR:-237.7 LO:237.7);ALT=C[chr6:24327808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24667572	+	chr6	24698109	+	.	0	10	2748731_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2748731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24647001_24672001_419C;SPAN=30537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=G[chr6:24698109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24714669	+	chr6	24716375	+	.	2	6	2748416_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2748416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24696001_24721001_182C;SPAN=1706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:6 DR:2 LR:-1.754 LO:15.04);ALT=C[chr6:24716375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24716554	+	chr6	24718768	+	.	3	5	2748424_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2748424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24696001_24721001_114C;SPAN=2214;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:5 DR:3 LR:-2.838 LO:15.21);ALT=T[chr6:24718768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	24811887	+	chr6	24817951	+	.	35	35	2749183_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CGTTTAGTACTT;MAPQ=60;MATEID=2749183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_24794001_24819001_414C;SPAN=6064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:72 GQ:6 PL:[184.8, 6.0, 0.0] SR:35 DR:35 LR:-190.6 LO:190.6);ALT=T[chr6:24817951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	25016063	+	chr6	25042077	+	.	8	7	2749685_1	29.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=2749685_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_25014501_25039501_180C;SPAN=26014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:51 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:7 DR:8 LR:-29.1 LO:31.04);ALT=C[chr6:25042077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	25016097	+	chr6	25036305	+	.	17	0	2749688_1	25.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2749688_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:25016097(+)-6:25036305(-)__6_25014501_25039501D;SPAN=20208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:113 GQ:25.7 PL:[25.7, 0.0, 246.8] SR:0 DR:17 LR:-25.5 LO:36.2);ALT=C[chr6:25036305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	25963512	+	chr6	25966562	+	.	5	3	2752858_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2752858_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_25945501_25970501_349C;SPAN=3050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:87 GQ:6.9 PL:[0.0, 6.9, 224.4] SR:3 DR:5 LR:7.065 LO:8.445);ALT=T[chr6:25966562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	26124979	+	chr6	26138280	+	.	7	6	2753347_1	11.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2753347_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_26117001_26142001_364C;SPAN=13301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:90 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:6 DR:7 LR:-11.93 LO:22.35);ALT=T[chr6:26138280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	26538729	+	chr6	26545354	+	.	62	22	2754921_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2754921_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_26533501_26558501_393C;SPAN=6625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:128 GQ:99 PL:[193.1, 0.0, 117.2] SR:22 DR:62 LR:-194.1 LO:194.1);ALT=G[chr6:26545354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
