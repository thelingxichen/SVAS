chr16	21594442	+	chr16	22710751	-	CAT	157	51	9221280_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CAT;MAPQ=60;MATEID=9221280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_22687001_22712001_375C;SPAN=1116309;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:197 DP:90 GQ:53.2 PL:[584.2, 53.2, 0.0] SR:51 DR:157 LR:-584.2 LO:584.2);ALT=C]chr16:22710751];VARTYPE=BND:INV-hh;JOINTYPE=hh
