chr7	115624568	+	chr7	115670685	+	.	27	7	3539054_1	77.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=3539054_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_115664501_115689501_303C;SPAN=46117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:56 GQ:57.5 PL:[77.3, 0.0, 57.5] SR:7 DR:27 LR:-77.39 LO:77.39);ALT=C[chr7:115670685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	115892533	+	chr7	115897347	+	.	4	3	3539790_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=3539790_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_115885001_115910001_133C;SPAN=4814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:124 GQ:16.8 PL:[0.0, 16.8, 333.3] SR:3 DR:4 LR:17.09 LO:7.662);ALT=G[chr7:115897347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	116502740	+	chr7	116538825	+	.	25	0	3541831_1	67.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3541831_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:116502740(+)-7:116538825(-)__7_116497501_116522501D;SPAN=36085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:57 GQ:67.1 PL:[67.1, 0.0, 70.4] SR:0 DR:25 LR:-67.08 LO:67.09);ALT=G[chr7:116538825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	116502740	+	chr7	116533046	+	.	22	0	3541830_1	57.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3541830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:116502740(+)-7:116533046(-)__7_116497501_116522501D;SPAN=30306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:57 GQ:57.2 PL:[57.2, 0.0, 80.3] SR:0 DR:22 LR:-57.18 LO:57.41);ALT=G[chr7:116533046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	116502740	+	chr7	116528178	+	.	15	0	3541829_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3541829_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:116502740(+)-7:116528178(-)__7_116497501_116522501D;SPAN=25438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:57 GQ:34.1 PL:[34.1, 0.0, 103.4] SR:0 DR:15 LR:-34.07 LO:36.06);ALT=G[chr7:116528178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	116502758	+	chr7	116544228	+	.	15	0	3541832_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3541832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:116502758(+)-7:116544228(-)__7_116497501_116522501D;SPAN=41470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:0 DR:15 LR:-33.8 LO:35.92);ALT=C[chr7:116544228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
