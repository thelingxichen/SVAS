chr16	46715461	+	chr16	46723042	+	.	11	0	6203951_1	27.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6203951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:46715461(+)-16:46723042(-)__16_46721501_46746501D;SPAN=7581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:32 GQ:27.8 PL:[27.8, 0.0, 47.6] SR:0 DR:11 LR:-27.64 LO:28.0);ALT=A[chr16:46723042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	46837016	+	chr16	46843514	+	.	11	0	6204028_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6204028_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:46837016(+)-16:46843514(-)__16_46819501_46844501D;SPAN=6498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:0 DR:11 LR:-23.31 LO:25.67);ALT=G[chr16:46843514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	46843702	+	chr16	46858298	+	.	0	18	6204043_1	53.0	.	EVDNC=ASSMB;HOMSEQ=CTGTA;MAPQ=60;MATEID=6204043_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_46844001_46869001_69C;SPAN=14596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:24 GQ:3.5 PL:[53.0, 0.0, 3.5] SR:18 DR:0 LR:-55.19 LO:55.19);ALT=A[chr16:46858298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	46843749	+	chr16	46864993	+	.	13	0	6204044_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6204044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:46843749(+)-16:46864993(-)__16_46844001_46869001D;SPAN=21244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:22 GQ:14 PL:[37.1, 0.0, 14.0] SR:0 DR:13 LR:-37.38 LO:37.38);ALT=G[chr16:46864993[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	46858398	+	chr16	46864994	+	.	25	10	6204064_1	80.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=ACCTGT;MAPQ=60;MATEID=6204064_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_46844001_46869001_26C;SPAN=6596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:43 GQ:21.5 PL:[80.9, 0.0, 21.5] SR:10 DR:25 LR:-82.52 LO:82.52);ALT=T[chr16:46864994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	47002076	+	chr16	47005261	+	.	0	15	6204464_1	32.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6204464_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_46991001_47016001_234C;SPAN=3185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:15 DR:0 LR:-32.72 LO:35.42);ALT=T[chr16:47005261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	47005484	+	chr16	47007405	+	TTTGTCTCCTGCATTTGGATTCTTATCAGGATGATATTCCTTGGCTAACTTTCTGTATG	25	57	6204470_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=CCTT;INSERTION=TTTGTCTCCTGCATTTGGATTCTTATCAGGATGATATTCCTTGGCTAACTTTCTGTATG;MAPQ=60;MATEID=6204470_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_46991001_47016001_76C;SPAN=1921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:60 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:57 DR:25 LR:-201.3 LO:201.3);ALT=A[chr16:47007405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	47005922	+	chr16	47007505	+	.	28	0	6204473_1	81.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6204473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:47005922(+)-16:47007505(-)__16_46991001_47016001D;SPAN=1583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:42 GQ:18.5 PL:[81.2, 0.0, 18.5] SR:0 DR:28 LR:-83.03 LO:83.03);ALT=T[chr16:47007505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	47488069	+	chr16	47494748	+	TTGAAAGATACCTTTACTTTGGGTTTAAAATAGGGTGCATTCTGGTCTGCCAAAAAGACGATTAAGTCATTT	0	26	6205137_1	71.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTGAAAGATACCTTTACTTTGGGTTTAAAATAGGGTGCATTCTGGTCTGCCAAAAAGACGATTAAGTCATTT;MAPQ=60;MATEID=6205137_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_47481001_47506001_206C;SPAN=6679;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:53 GQ:55.1 PL:[71.6, 0.0, 55.1] SR:26 DR:0 LR:-71.55 LO:71.55);ALT=C[chr16:47494748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	47493124	+	chr16	47494905	+	.	11	0	6205146_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6205146_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:47493124(+)-16:47494905(-)__16_47481001_47506001D;SPAN=1781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:61 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-19.78 LO:24.38);ALT=G[chr16:47494905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	48295498	+	chr16	48296687	+	.	2	5	6206185_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6206185_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_48289501_48314501_265C;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:52 GQ:2.6 PL:[2.6, 0.0, 121.4] SR:5 DR:2 LR:-2.417 LO:9.606);ALT=G[chr16:48296687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
