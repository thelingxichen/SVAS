chrom_5p	bkpos_5p	strand_5p	chrom_3p	bkpos_3p	strand_3p	junc_reads	span_reads	id	qual	filter	meta_info
chr3	169201745	+	chr1	6259596	+	.	36	0	1779497_1	94.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=1779497_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6259596(-)-3:169201745(+)__3_169197001_169222001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:89 GQ:94.7 PL:[94.7, 0.0, 121.1] SR:0 DR:36 LR:-94.72 LO:94.9);ALT=]chr3:169201745]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	6845683	+	chr1	6885148	+	.	47	0	19397_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=19397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6845683(+)-1:6885148(-)__1_6884501_6909501D;SPAN=39465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=G[chr1:6885148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8021854	+	chr1	8025383	+	CTTGTAAACATATAACATAAAAATGGCTTCCAAAAGAGCTCTGGTCATCCTGGCTAAAGGAGCAGAGGAAATGGAGACGGTCATCCCTGTAGATGTCATGAGGCGAGCTGG	61	131	22705_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTTGTAAACATATAACATAAAAATGGCTTCCAAAAGAGCTCTGGTCATCCTGGCTAAAGGAGCAGAGGAAATGGAGACGGTCATCCCTGTAGATGTCATGAGGCGAGCTGG;MAPQ=60;MATEID=22705_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_8011501_8036501_97C;SPAN=3529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:99 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:131 DR:61 LR:-458.8 LO:458.8);ALT=G[chr1:8025383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8924153	+	chr1	8925344	+	.	32	12	25213_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=9;MATEID=25213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8918001_8943001_29C;SPAN=1191;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:78 GQ:64.7 PL:[124.1, 0.0, 64.7] SR:12 DR:32 LR:-125.1 LO:125.1);ALT=T[chr1:8925344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8934978	+	chr1	8938639	+	.	122	58	25255_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=43;MATEID=25255_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8918001_8943001_205C;SPAN=3661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:108 GQ:36 PL:[396.0, 36.0, 0.0] SR:58 DR:122 LR:-396.1 LO:396.1);ALT=T[chr1:8938639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8938639	-	chr1	236646440	+	.	163	19	617066_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CTAGCCACTGGGTCTC;MAPQ=60;MATEID=617066_2;MATENM=12;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_1_236645501_236670501_12C;SPAN=227707801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:182 DP:79 GQ:49 PL:[538.0, 49.0, 0.0] SR:19 DR:163 LR:-538.0 LO:538.0);ALT=[chr1:236646440[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	11796295	+	chr1	11807496	+	ATTCTCCTAGGTCACTGGCTGCTGACAACCT	36	11	34432_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATTCTCCTAGGTCACTGGCTGCTGACAACCT;MAPQ=60;MATEID=34432_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_11784501_11809501_105C;SPAN=11201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:81 GQ:93.8 PL:[100.4, 0.0, 93.8] SR:11 DR:36 LR:-100.2 LO:100.2);ALT=G[chr1:11807496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16154742	-	chr19	39926488	+	.	72	47	47148_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=CCGCTGCAGTCGGTGCAGGTCTTCGGACGCAAG;MAPQ=55;MATEID=47148_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_1_16145501_16170501_79C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:92 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:47 DR:72 LR:-283.9 LO:283.9);ALT=[chr19:39926488[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	16693823	+	chr1	16719723	+	.	48	0	48680_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=48680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:16693823(+)-1:16719723(-)__1_16684501_16709501D;SPAN=25900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:49 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:48 LR:-145.2 LO:145.2);ALT=C[chr1:16719723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17051748	-	chr1	234912188	+	GCCCCATCCCGCCGGCTTCTGC	189	57	50768_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;INSERTION=GCCCCATCCCGCCGGCTTCTGC;MAPQ=60;MATEID=50768_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17027501_17052501_901C;SPAN=217860440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:229 DP:175 GQ:61.9 PL:[679.9, 61.9, 0.0] SR:57 DR:189 LR:-680.0 LO:680.0);ALT=[chr1:234912188[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	17371386	+	chr1	17380442	+	.	34	6	53672_1	95.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=53672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17370501_17395501_125C;SPAN=9056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:74 GQ:82.4 PL:[95.6, 0.0, 82.4] SR:6 DR:34 LR:-95.52 LO:95.52);ALT=G[chr1:17380442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17634809	+	chr1	17657461	+	.	37	10	54878_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=54878_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_17640001_17665001_160C;SPAN=22652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:53 GQ:5.6 PL:[121.1, 0.0, 5.6] SR:10 DR:37 LR:-126.9 LO:126.9);ALT=G[chr1:17657461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17676184	+	chr1	17677654	+	.	47	20	54994_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CTGCACTCCAGCCTGGGTGACAGA;MAPQ=60;MATEID=54994_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_17664501_17689501_17C;SPAN=1470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:33 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:20 DR:47 LR:-184.8 LO:184.8);ALT=A[chr1:17677654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21107034	+	chr1	21113005	+	.	33	6	64936_1	90.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=64936_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_27C;SPAN=5971;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:92 GQ:90.8 PL:[90.8, 0.0, 130.4] SR:6 DR:33 LR:-90.61 LO:91.04);ALT=C[chr1:21113005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21107035	+	chr1	21113686	+	.	34	8	64938_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=64938_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_122C;SPAN=6651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:67 GQ:57.8 PL:[104.0, 0.0, 57.8] SR:8 DR:34 LR:-104.7 LO:104.7);ALT=T[chr1:21113686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21822955	+	chr1	21828058	+	.	50	47	67085_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=67085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21805001_21830001_245C;SPAN=5103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:47 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:47 DR:50 LR:-211.3 LO:211.3);ALT=G[chr1:21828058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	22379323	+	chr4	22729560	-	.	33	0	1920745_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1920745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:22379323(+)-4:22729560(+)__4_22711501_22736501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:50 GQ:26 PL:[95.3, 0.0, 26.0] SR:0 DR:33 LR:-97.6 LO:97.6);ALT=C]chr4:22729560];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	24969839	+	chrX	136067839	-	.	62	19	7535206_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7535206_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_23_136048501_136073501_21C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:26 GQ:21 PL:[231.0, 21.0, 0.0] SR:19 DR:62 LR:-231.1 LO:231.1);ALT=G]chrX:136067839];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	24969882	+	chr1	24973155	+	.	56	0	76459_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=76459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24969882(+)-1:24973155(-)__1_24965501_24990501D;SPAN=3273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:84 GQ:40.1 PL:[162.2, 0.0, 40.1] SR:0 DR:56 LR:-166.1 LO:166.1);ALT=C[chr1:24973155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25158703	+	chr1	25161510	+	.	60	51	77252_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTGATTTTTTATTTTT;MAPQ=60;MATEID=77252_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_25137001_25162001_156C;SPAN=2807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:32 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:51 DR:60 LR:-260.8 LO:260.8);ALT=T[chr1:25161510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25555664	+	chr1	25558930	+	.	50	0	78382_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=78382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25555664(+)-1:25558930(-)__1_25553501_25578501D;SPAN=3266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:113 GQ:99 PL:[134.6, 0.0, 137.9] SR:0 DR:50 LR:-134.4 LO:134.4);ALT=C[chr1:25558930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25664911	+	chr1	25669451	+	.	39	0	78319_1	98.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=78319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25664911(+)-1:25669451(-)__1_25651501_25676501D;SPAN=4540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:110 GQ:98.9 PL:[98.9, 0.0, 168.2] SR:0 DR:39 LR:-98.94 LO:99.92);ALT=C[chr1:25669451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25664947	+	chr1	25666965	+	.	60	41	78320_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=78320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25651501_25676501_199C;SPAN=2018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:107 GQ:20.6 PL:[238.4, 0.0, 20.6] SR:41 DR:60 LR:-249.1 LO:249.1);ALT=C[chr1:25666965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26228230	+	chr1	26231153	+	.	52	0	79997_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=79997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26228230(+)-1:26231153(-)__1_26215001_26240001D;SPAN=2923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:83 GQ:50.3 PL:[149.3, 0.0, 50.3] SR:0 DR:52 LR:-151.7 LO:151.7);ALT=G[chr1:26231153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26230334	+	chr1	26232878	+	.	37	0	80001_1	72.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=80001_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26230334(+)-1:26232878(-)__1_26215001_26240001D;SPAN=2544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:183 GQ:72.7 PL:[72.7, 0.0, 369.8] SR:0 DR:37 LR:-72.56 LO:84.05);ALT=A[chr1:26232878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26460160	+	chr1	26464769	+	.	31	0	80780_1	92.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=80780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26460160(+)-1:26464769(-)__1_26435501_26460501D;SPAN=4609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:32 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:31 LR:-92.42 LO:92.42);ALT=G[chr1:26464769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26644562	+	chr1	26646657	+	.	96	39	81416_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TACAG;MAPQ=60;MATEID=81416_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_26631501_26656501_208C;SPAN=2095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:121 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:39 DR:96 LR:-356.5 LO:356.5);ALT=G[chr1:26646657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27668642	+	chr1	27671785	+	.	78	10	84847_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=84847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27660501_27685501_160C;SPAN=3143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:89 GQ:24 PL:[264.0, 24.0, 0.0] SR:10 DR:78 LR:-264.1 LO:264.1);ALT=G[chr1:27671785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27755454	+	chr1	27816503	+	.	32	0	85404_1	91.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=85404_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27755454(+)-1:27816503(-)__1_27807501_27832501D;SPAN=61049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:53 GQ:35.3 PL:[91.4, 0.0, 35.3] SR:0 DR:32 LR:-92.5 LO:92.5);ALT=A[chr1:27816503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27950441	+	chr1	27961574	+	CCTTAGGCCCCTACTCCTGGGTCAGTGGGGCTGCGGCATGATCCTTGGGAGGGGTCAGAG	31	21	85581_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=CCTTAGGCCCCTACTCCTGGGTCAGTGGGGCTGCGGCATGATCCTTGGGAGGGGTCAGAG;MAPQ=60;MATEID=85581_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_27954501_27979501_302C;SPAN=11133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:30 GQ:12 PL:[132.0, 12.0, 0.0] SR:21 DR:31 LR:-132.0 LO:132.0);ALT=C[chr1:27961574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48481808	+	chr1	27975966	+	.	31	0	1395853_1	86.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=1395853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27975966(-)-3:48481808(+)__3_48461001_48486001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:59 GQ:56.6 PL:[86.3, 0.0, 56.6] SR:0 DR:31 LR:-86.67 LO:86.67);ALT=]chr3:48481808]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	27995096	+	chr1	27998631	+	.	38	0	85776_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=85776_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27995096(+)-1:27998631(-)__1_27979001_28004001D;SPAN=3535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:78 GQ:84.5 PL:[104.3, 0.0, 84.5] SR:0 DR:38 LR:-104.4 LO:104.4);ALT=G[chr1:27998631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28555536	+	chr1	28559427	+	.	32	11	87658_1	98.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=TTCACCT;MAPQ=60;MATEID=87658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28542501_28567501_63C;SPAN=3891;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:75 GQ:82.1 PL:[98.6, 0.0, 82.1] SR:11 DR:32 LR:-98.58 LO:98.58);ALT=T[chr1:28559427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28559446	-	chr14	35899082	+	.	41	0	5702808_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5702808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28559446(-)-14:35899082(-)__14_35892501_35917501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=[chr14:35899082[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	28832645	+	chr1	28835338	+	.	128	0	88659_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=88659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28832645(+)-1:28835338(-)__1_28812001_28837001D;SPAN=2693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:74 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:0 DR:128 LR:-379.6 LO:379.6);ALT=G[chr1:28835338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28948676	+	chr1	28969502	+	.	34	0	89185_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=89185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28948676(+)-1:28969502(-)__1_28959001_28984001D;SPAN=20826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:0 DR:34 LR:-110.1 LO:110.1);ALT=A[chr1:28969502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	30738623	+	chr1	30739932	+	.	48	32	93508_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCA;MAPQ=60;MATEID=93508_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_30723001_30748001_14C;SPAN=1309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:36 GQ:18 PL:[198.0, 18.0, 0.0] SR:32 DR:48 LR:-198.0 LO:198.0);ALT=A[chr1:30739932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31214612	+	chr1	31230553	+	.	98	0	94531_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=94531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31214612(+)-1:31230553(-)__1_31213001_31238001D;SPAN=15941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:118 GQ:5.4 PL:[297.0, 5.4, 0.0] SR:0 DR:98 LR:-310.9 LO:310.9);ALT=C[chr1:31230553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31215397	+	chr1	31230506	+	.	102	28	94534_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=94534_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_31213001_31238001_235C;SPAN=15109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:127 GQ:14.4 PL:[336.6, 14.4, 0.0] SR:28 DR:102 LR:-345.9 LO:345.9);ALT=C[chr1:31230506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31568380	+	chr19	48282071	-	CGCCA	84	30	6842369_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;INSERTION=CGCCA;MAPQ=60;MATEID=6842369_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48265001_48290001_363C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:47 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:30 DR:84 LR:-310.3 LO:310.3);ALT=G]chr19:48282071];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	32688221	+	chr1	32690009	+	.	52	0	99289_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=99289_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32688221(+)-1:32690009(-)__1_32683001_32708001D;SPAN=1788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:102 GQ:99 PL:[144.2, 0.0, 101.3] SR:0 DR:52 LR:-144.4 LO:144.4);ALT=C[chr1:32690009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32688231	+	chr1	32689635	+	.	47	46	99292_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=99292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32683001_32708001_238C;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:86 GQ:23 PL:[184.7, 0.0, 23.0] SR:46 DR:47 LR:-191.8 LO:191.8);ALT=T[chr1:32689635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35449601	+	chr1	35450813	+	.	33	0	106412_1	87.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=106412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:35449601(+)-1:35450813(-)__1_35427001_35452001D;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:80 GQ:87.2 PL:[87.2, 0.0, 107.0] SR:0 DR:33 LR:-87.26 LO:87.37);ALT=C[chr1:35450813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36102034	+	chr1	36106943	+	.	66	62	108395_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=108395_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36088501_36113501_108C;SPAN=4909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:96 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:62 DR:66 LR:-283.9 LO:283.9);ALT=C[chr1:36106943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36690152	+	chr1	36748129	+	.	34	0	110059_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=110059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36690152(+)-1:36748129(-)__1_36725501_36750501D;SPAN=57977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:32 GQ:9 PL:[99.0, 9.0, 0.0] SR:0 DR:34 LR:-99.02 LO:99.02);ALT=T[chr1:36748129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36859755	+	chr1	36863368	+	.	65	24	110817_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=110817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36848001_36873001_338C;SPAN=3613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:91 GQ:8.6 PL:[209.9, 0.0, 8.6] SR:24 DR:65 LR:-220.4 LO:220.4);ALT=C[chr1:36863368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	37979140	+	chr1	37980257	+	.	36	15	113595_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=113595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_37975001_38000001_17C;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:71 GQ:43.7 PL:[126.2, 0.0, 43.7] SR:15 DR:36 LR:-128.0 LO:128.0);ALT=C[chr1:37980257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39492070	+	chr1	39494394	+	.	117	5	117884_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=117884_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_39494001_39519001_2C;SPAN=2324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:43 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:5 DR:117 LR:-346.6 LO:346.6);ALT=G[chr1:39494394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39492106	+	chr17	27348522	-	.	43	0	117765_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=117765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:39492106(+)-17:27348522(+)__1_39469501_39494501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:34 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=A]chr17:27348522];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	40506524	+	chr1	40525736	+	.	33	0	121105_1	92.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=121105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40506524(+)-1:40525736(-)__1_40523001_40548001D;SPAN=19212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:59 GQ:50 PL:[92.9, 0.0, 50.0] SR:0 DR:33 LR:-93.63 LO:93.63);ALT=G[chr1:40525736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40558228	+	chr1	40562854	+	.	65	0	120961_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=120961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40558228(+)-1:40562854(-)__1_40547501_40572501D;SPAN=4626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:98 GQ:49.4 PL:[188.0, 0.0, 49.4] SR:0 DR:65 LR:-192.5 LO:192.5);ALT=T[chr1:40562854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	42922318	+	chr1	42925264	+	.	38	0	127171_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=127171_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:42922318(+)-1:42925264(-)__1_42899501_42924501D;SPAN=2946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:42 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:38 LR:-122.1 LO:122.1);ALT=G[chr1:42925264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	43124184	+	chr11	111901010	-	CATGCGGCCAACTT	65	6	5004785_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CATGCGGCCAACTT;MAPQ=60;MATEID=5004785_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_11_111891501_111916501_91C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:40 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:6 DR:65 LR:-208.0 LO:208.0);ALT=G]chr11:111901010];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	43831334	+	chr1	43833585	+	.	32	0	129737_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=129737_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:43831334(+)-1:43833585(-)__1_43806001_43831001D;SPAN=2251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:0 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=T[chr1:43833585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45981520	+	chr1	45987349	+	.	174	0	136055_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=136055_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45981520(+)-1:45987349(-)__1_45986501_46011501D;SPAN=5829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:45 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:0 DR:174 LR:-514.9 LO:514.9);ALT=A[chr1:45987349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45984765	+	chr1	45987381	+	.	79	0	136057_1	99.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=136057_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45984765(+)-1:45987381(-)__1_45986501_46011501D;SPAN=2616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:52 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=T[chr1:45987381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46016876	+	chr1	46032232	+	.	33	0	135744_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=135744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46016876(+)-1:46032232(-)__1_46011001_46036001D;SPAN=15356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=T[chr1:46032232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46049805	+	chr1	46067923	+	.	38	0	136446_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=136446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46049805(+)-1:46067923(-)__1_46035501_46060501D;SPAN=18118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:44 GQ:8.4 PL:[122.1, 8.4, 0.0] SR:0 DR:38 LR:-122.5 LO:122.5);ALT=A[chr1:46067923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	45872386	+	chr1	47804186	+	.	60	42	2830453_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TCCCT;MAPQ=60;MATEID=2830453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_45864001_45889001_51C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:29 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:42 DR:60 LR:-211.3 LO:211.3);ALT=]chr6:45872386]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	59096879	+	chr2	32048671	+	.	38	0	168730_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=168730_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:59096879(+)-2:32048671(-)__1_59094001_59119001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:64 GQ:45.5 PL:[108.2, 0.0, 45.5] SR:0 DR:38 LR:-109.4 LO:109.4);ALT=A[chr2:32048671[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	71544391	+	chr1	71546623	+	.	44	9	197185_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=197185_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_1_71540001_71565001_274C;SPAN=2232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:73 GQ:29.9 PL:[145.4, 0.0, 29.9] SR:9 DR:44 LR:-149.4 LO:149.4);ALT=T[chr1:71546623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84517939	+	chr1	84524630	+	.	41	15	224957_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGATTTGTTTTTCT;MAPQ=60;MATEID=224957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84500501_84525501_206C;SPAN=6691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:62 GQ:6.5 PL:[141.8, 0.0, 6.5] SR:15 DR:41 LR:-148.6 LO:148.6);ALT=T[chr1:84524630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	109590094	+	chr1	84971740	+	.	53	0	225534_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=225534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:84971740(-)-23:109590094(+)__1_84966001_84991001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:72 GQ:17 PL:[155.6, 0.0, 17.0] SR:0 DR:53 LR:-161.6 LO:161.6);ALT=]chrX:109590094]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	87170654	+	chr1	87181404	+	.	33	15	231018_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=231018_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_87146501_87171501_143C;SPAN=10750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:29 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:15 DR:33 LR:-112.2 LO:112.2);ALT=G[chr1:87181404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	87369132	+	chr1	87379708	+	.	74	16	231094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=231094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_87367001_87392001_123C;SPAN=10576;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:61 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:16 DR:74 LR:-237.7 LO:237.7);ALT=C[chr1:87379708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	88972810	-	chr17	32063850	+	.	48	19	6371204_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6371204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_32046001_32071001_107C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:41 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:19 DR:48 LR:-158.4 LO:158.4);ALT=[chr17:32063850[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	89570519	+	chr12	57081784	+	.	125	0	5205294_1	99.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=5205294_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:89570519(+)-12:57081784(-)__12_57060501_57085501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:72 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:0 DR:125 LR:-369.7 LO:369.7);ALT=T[chr12:57081784[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	93297682	+	chr1	93299099	+	.	50	0	240745_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=240745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93297682(+)-1:93299099(-)__1_93296001_93321001D;SPAN=1417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:128 GQ:99 PL:[130.4, 0.0, 179.9] SR:0 DR:50 LR:-130.4 LO:130.8);ALT=G[chr1:93299099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93805158	+	chr1	93811280	+	.	59	0	241420_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=241420_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93805158(+)-1:93811280(-)__1_93810501_93835501D;SPAN=6122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:19 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=T[chr1:93811280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	94288375	+	chr1	94291257	+	.	69	27	242166_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CCA;MAPQ=60;MATEID=242166_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_94276001_94301001_16C;SPAN=2882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:22 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:27 DR:69 LR:-254.2 LO:254.2);ALT=A[chr1:94291257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	94343442	+	chr1	94344635	+	.	35	0	242407_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=242407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:94343442(+)-1:94344635(-)__1_94325001_94350001D;SPAN=1193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:57 GQ:37.4 PL:[100.1, 0.0, 37.4] SR:0 DR:35 LR:-101.6 LO:101.6);ALT=G[chr1:94344635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109958043	+	chr1	109968976	+	.	44	0	263428_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=263428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109958043(+)-1:109968976(-)__1_109956001_109981001D;SPAN=10933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:60 GQ:16.7 PL:[128.9, 0.0, 16.7] SR:0 DR:44 LR:-134.0 LO:134.0);ALT=C[chr1:109968976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110230551	+	chr6	111368672	-	.	82	0	2984550_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2984550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110230551(+)-6:111368672(+)__6_111352501_111377501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:47 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=A]chr6:111368672];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	110944251	+	chr1	110950206	+	.	40	0	265035_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=265035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110944251(+)-1:110950206(-)__1_110936001_110961001D;SPAN=5955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:74 GQ:65.9 PL:[112.1, 0.0, 65.9] SR:0 DR:40 LR:-112.6 LO:112.6);ALT=C[chr1:110950206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110946658	+	chr1	110950208	+	AATGAAGAATCCCTCCATTGTTGGAGTCCTGTGCACAGATTCACAAGGACTTAATCTGGGTT	61	52	265041_1	99.0	.	DISC_MAPQ=39;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATGAAGAATCCCTCCATTGTTGGAGTCCTGTGCACAGATTCACAAGGACTTAATCTGGGTT;MAPQ=60;MATEID=265041_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_110936001_110961001_85C;SPAN=3550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:79 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:52 DR:61 LR:-290.5 LO:290.5);ALT=C[chr1:110950208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111415871	+	chr1	111434012	+	.	37	10	265768_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=265768_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_111426001_111451001_77C;SPAN=18141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:23 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:10 DR:37 LR:-112.2 LO:112.2);ALT=G[chr1:111434012[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111415908	+	chr1	111434965	+	.	72	0	265771_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=265771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111415908(+)-1:111434965(-)__1_111426001_111451001D;SPAN=19057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:41 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:0 DR:72 LR:-211.3 LO:211.3);ALT=A[chr1:111434965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111992219	+	chr1	111996831	+	.	83	0	266598_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=266598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111992219(+)-1:111996831(-)__1_111989501_112014501D;SPAN=4612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:71 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:0 DR:83 LR:-244.3 LO:244.3);ALT=C[chr1:111996831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112691792	+	chr1	112704704	+	.	68	26	267593_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=267593_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_1_112675501_112700501_71C;SPAN=12912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:7 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:26 DR:68 LR:-241.0 LO:241.0);ALT=G[chr1:112704704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	44038799	+	chr1	146649791	+	.	36	0	5938554_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5938554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146649791(-)-15:44038799(+)__15_44026501_44051501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:61 GQ:43.1 PL:[102.5, 0.0, 43.1] SR:0 DR:36 LR:-103.5 LO:103.5);ALT=]chr15:44038799]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	146676498	+	chr21	30445877	+	.	74	0	307153_1	99.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=307153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146676498(+)-21:30445877(-)__1_146657001_146682001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:65 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:0 DR:74 LR:-217.9 LO:217.9);ALT=G[chr21:30445877[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	146702258	-	chr1	146818239	+	.	31	0	307686_1	89.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=307686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146702258(-)-1:146818239(-)__1_146804001_146829001D;SPAN=115981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:48 GQ:26.6 PL:[89.3, 0.0, 26.6] SR:0 DR:31 LR:-91.16 LO:91.16);ALT=[chr1:146818239[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	150266371	+	chr1	150280474	+	.	52	0	321972_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=321972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150266371(+)-1:150280474(-)__1_150258501_150283501D;SPAN=14103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:150 GQ:99 PL:[131.0, 0.0, 233.3] SR:0 DR:52 LR:-131.0 LO:132.6);ALT=A[chr1:150280474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150266869	+	chr1	150280478	+	.	35	51	321977_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ACAG;MAPQ=60;MATEID=321977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150258501_150283501_326C;SPAN=13609;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:134 GQ:86 PL:[237.8, 0.0, 86.0] SR:51 DR:35 LR:-241.5 LO:241.5);ALT=G[chr1:150280478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150730506	+	chr1	150738173	+	.	66	0	324108_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=324108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150730506(+)-1:150738173(-)__1_150724001_150749001D;SPAN=7667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:91 GQ:25.1 PL:[193.4, 0.0, 25.1] SR:0 DR:66 LR:-200.4 LO:200.4);ALT=A[chr1:150738173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151028472	+	chr1	151031954	+	.	44	11	325374_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=325374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151018001_151043001_167C;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:106 GQ:99 PL:[133.1, 0.0, 123.2] SR:11 DR:44 LR:-133.0 LO:133.0);ALT=G[chr1:151031954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151227321	+	chr10	95719620	-	.	76	0	4663360_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4663360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151227321(+)-10:95719620(+)__10_95697001_95722001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:31 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:0 DR:76 LR:-224.5 LO:224.5);ALT=G]chr10:95719620];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	151955849	+	chr1	151966225	+	.	91	0	329503_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=329503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151955849(+)-1:151966225(-)__1_151949001_151974001D;SPAN=10376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:91 DP:191 GQ:99 PL:[248.9, 0.0, 212.6] SR:0 DR:91 LR:-248.8 LO:248.8);ALT=T[chr1:151966225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151958729	+	chr1	151966227	+	.	142	17	329512_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=329512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151949001_151974001_205C;SPAN=7498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:151 DP:241 GQ:99 PL:[433.4, 0.0, 149.5] SR:17 DR:142 LR:-440.6 LO:440.6);ALT=T[chr1:151966227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	152005335	+	chr1	152009385	+	.	40	0	329888_1	95.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=329888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:152005335(+)-1:152009385(-)__1_151998001_152023001D;SPAN=4050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:136 GQ:95.3 PL:[95.3, 0.0, 233.9] SR:0 DR:40 LR:-95.2 LO:98.46);ALT=A[chr1:152009385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	152006277	+	chr1	152009388	+	.	120	24	329893_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=329893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151998001_152023001_209C;SPAN=3111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:141 DP:150 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:24 DR:120 LR:-445.6 LO:445.6);ALT=C[chr1:152009388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153330909	+	chr1	153333118	+	.	91	147	333846_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=333846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_153321001_153346001_137C;SPAN=2209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:218 DP:315 GQ:99 PL:[634.4, 0.0, 129.4] SR:147 DR:91 LR:-653.0 LO:653.0);ALT=G[chr1:153333118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153516400	+	chr1	153518229	+	CCCAAGAAGCTGGGCAGCTCCCGGGTCAGCAGCTCCTTTAGTTCTGACTTGTTGAGCTTGAACTTGTCACCCTCTTTGCCCGAGTACTTGTGGAAGGTGGACACCATCACATCCAGGGCCTTCTCCAGAGGGCACGCCATGACAGCAGTCAGGAT	50	99	334414_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCCAAGAAGCTGGGCAGCTCCCGGGTCAGCAGCTCCTTTAGTTCTGACTTGTTGAGCTTGAACTTGTCACCCTCTTTGCCCGAGTACTTGTGGAAGGTGGACACCATCACATCCAGGGCCTTCTCCAGAGGGCACGCCATGACAGCAGTCAGGAT;MAPQ=60;MATEID=334414_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_153492501_153517501_92C;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:123 DP:340 GQ:99 PL:[313.9, 0.0, 512.0] SR:99 DR:50 LR:-313.9 LO:316.5);ALT=C[chr1:153518229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153641105	+	chr1	153643392	+	.	58	0	334932_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=334932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153641105(+)-1:153643392(-)__1_153639501_153664501D;SPAN=2287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:111 GQ:99 PL:[161.6, 0.0, 105.5] SR:0 DR:58 LR:-161.9 LO:161.9);ALT=C[chr1:153643392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56374762	+	chr1	153958676	+	.	32	0	5202764_1	92.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5202764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153958676(-)-12:56374762(+)__12_56374501_56399501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:47 GQ:20.3 PL:[92.9, 0.0, 20.3] SR:0 DR:32 LR:-95.43 LO:95.43);ALT=]chr12:56374762]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	154148745	+	chr1	154155474	+	.	94	0	337633_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=337633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154148745(+)-1:154155474(-)__1_154154001_154179001D;SPAN=6729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:97 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:0 DR:94 LR:-287.2 LO:287.2);ALT=G[chr1:154155474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155145951	+	chr1	155151248	+	.	49	13	341400_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=341400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155134001_155159001_20C;SPAN=5297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:82 GQ:47.3 PL:[149.6, 0.0, 47.3] SR:13 DR:49 LR:-152.2 LO:152.2);ALT=C[chr1:155151248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155658973	+	chr1	155686794	+	.	35	0	343834_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=343834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155658973(+)-1:155686794(-)__1_155648501_155673501D;SPAN=27821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:54 GQ:28.4 PL:[101.0, 0.0, 28.4] SR:0 DR:35 LR:-103.0 LO:103.0);ALT=A[chr1:155686794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155984907	+	chr1	155990678	+	.	33	0	345740_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=345740_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155984907(+)-1:155990678(-)__1_155967001_155992001D;SPAN=5771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:149 GQ:68.6 PL:[68.6, 0.0, 293.0] SR:0 DR:33 LR:-68.57 LO:76.45);ALT=G[chr1:155990678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155988214	+	chr1	155990676	+	.	93	0	345760_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=345760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155988214(+)-1:155990676(-)__1_155967001_155992001D;SPAN=2462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:93 DP:145 GQ:83 PL:[267.8, 0.0, 83.0] SR:0 DR:93 LR:-273.0 LO:273.0);ALT=C[chr1:155990676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156304760	+	chr1	156307943	+	.	57	0	346887_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=346887_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156304760(+)-1:156307943(-)__1_156285501_156310501D;SPAN=3183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:134 GQ:99 PL:[152.0, 0.0, 171.8] SR:0 DR:57 LR:-151.9 LO:151.9);ALT=G[chr1:156307943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156526723	+	chr1	156528936	+	.	110	73	347636_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAATTGAGTAGCTCAGC;MAPQ=60;MATEID=347636_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_1_156506001_156531001_299C;SPAN=2213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:48 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:73 DR:110 LR:-432.4 LO:432.4);ALT=C[chr1:156528936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156708559	+	chr1	156710804	+	.	73	2	348902_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=348902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156702001_156727001_150C;SPAN=2245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:122 GQ:86 PL:[208.1, 0.0, 86.0] SR:2 DR:73 LR:-210.6 LO:210.6);ALT=G[chr1:156710804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	157348495	+	chr1	157457782	-	.	31	0	350898_1	89.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=350898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:157348495(+)-1:157457782(+)__1_157437001_157462001D;SPAN=109287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:27 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=T]chr1:157457782];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	158961355	+	chr1	158966212	+	CATGGT	129	74	355055_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=CATGGT;MAPQ=60;MATEID=355055_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_158956001_158981001_36C;SPAN=4857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:166 DP:55 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:74 DR:129 LR:-491.8 LO:491.8);ALT=G[chr1:158966212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159889673	+	chr1	159895237	+	.	92	0	358330_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=358330_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159889673(+)-1:159895237(-)__1_159887001_159912001D;SPAN=5564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:304 GQ:99 PL:[221.5, 0.0, 515.3] SR:0 DR:92 LR:-221.3 LO:227.8);ALT=C[chr1:159895237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159890358	+	chr1	159895237	+	.	112	0	358338_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=358338_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159890358(+)-1:159895237(-)__1_159887001_159912001D;SPAN=4879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:295 GQ:99 PL:[289.9, 0.0, 425.3] SR:0 DR:112 LR:-289.8 LO:291.2);ALT=C[chr1:159895237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	21958921	+	chr1	160864770	+	.	36	0	361704_1	99.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=361704_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:160864770(-)-23:21958921(+)__1_160842501_160867501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:70 GQ:70.1 PL:[99.8, 0.0, 70.1] SR:0 DR:36 LR:-100.2 LO:100.2);ALT=]chrX:21958921]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	161072167	+	chr1	161087738	+	.	142	20	362607_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCACCT;MAPQ=60;MATEID=362607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161063001_161088001_274C;SPAN=15571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:113 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:20 DR:142 LR:-448.9 LO:448.9);ALT=T[chr1:161087738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161123910	+	chr1	161126739	+	.	46	60	362922_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=362922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161112001_161137001_325C;SPAN=2829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:84 DP:132 GQ:76.7 PL:[241.7, 0.0, 76.7] SR:60 DR:46 LR:-246.1 LO:246.1);ALT=G[chr1:161126739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161123929	+	chr1	161127042	+	.	40	0	362924_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=362924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161123929(+)-1:161127042(-)__1_161112001_161137001D;SPAN=3113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:137 GQ:95 PL:[95.0, 0.0, 236.9] SR:0 DR:40 LR:-94.92 LO:98.31);ALT=G[chr1:161127042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161172305	+	chr1	161176195	+	.	35	0	362703_1	86.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=362703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161172305(+)-1:161176195(-)__1_161161001_161186001D;SPAN=3890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:109 GQ:86 PL:[86.0, 0.0, 178.4] SR:0 DR:35 LR:-86.01 LO:87.78);ALT=C[chr1:161176195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161185160	+	chr1	161187773	+	.	38	2	362759_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=362759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161161001_161186001_355C;SPAN=2613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:2 DR:38 LR:-120.9 LO:120.9);ALT=G[chr1:161187773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600530	+	chr1	165619075	+	.	52	14	379424_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=379424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165595501_165620501_23C;SPAN=18545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:161 GQ:99 PL:[138.2, 0.0, 250.4] SR:14 DR:52 LR:-137.9 LO:139.8);ALT=G[chr1:165619075[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600578	+	chr1	165621212	+	.	41	0	379508_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=379508_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:165600578(+)-1:165621212(-)__1_165620001_165645001D;SPAN=20634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:61 GQ:26.6 PL:[119.0, 0.0, 26.6] SR:0 DR:41 LR:-121.8 LO:121.8);ALT=G[chr1:165621212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600581	+	chr1	165620247	+	.	90	0	379509_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=379509_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:165600581(+)-1:165620247(-)__1_165620001_165645001D;SPAN=19666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:88 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:0 DR:90 LR:-267.4 LO:267.4);ALT=C[chr1:165620247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167599667	+	chr1	167653135	+	.	31	24	386823_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=386823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167580001_167605001_296C;SPAN=53468;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:74 GQ:52.7 PL:[125.3, 0.0, 52.7] SR:24 DR:31 LR:-126.7 LO:126.7);ALT=G[chr1:167653135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168024574	+	chr1	168025733	+	.	106	53	387728_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGGCTTAAGTTTTT;MAPQ=60;MATEID=387728_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_168021001_168046001_352C;SPAN=1159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:82 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:53 DR:106 LR:-379.6 LO:379.6);ALT=T[chr1:168025733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168186489	+	chr3	53175885	+	TT	83	83	388883_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TT;MAPQ=60;MATEID=388883_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_168168001_168193001_141C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:62 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:83 DR:83 LR:-366.4 LO:366.4);ALT=T[chr3:53175885[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	169677993	+	chr1	169680636	+	.	40	0	393052_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=393052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169677993(+)-1:169680636(-)__1_169662501_169687501D;SPAN=2643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:112 GQ:99 PL:[101.9, 0.0, 167.9] SR:0 DR:40 LR:-101.7 LO:102.6);ALT=A[chr1:169680636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	173446631	+	chr1	173450465	+	.	100	60	404769_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=404769_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_173435501_173460501_334C;SPAN=3834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:118 GQ:36 PL:[396.0, 36.0, 0.0] SR:60 DR:100 LR:-396.1 LO:396.1);ALT=C[chr1:173450465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	174969358	+	chr1	174973747	+	.	52	0	410248_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=410248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:174969358(+)-1:174973747(-)__1_174954501_174979501D;SPAN=4389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:110 GQ:99 PL:[141.8, 0.0, 125.3] SR:0 DR:52 LR:-141.9 LO:141.9);ALT=A[chr1:174973747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	175200569	+	chr1	175201937	-	.	50	55	411167_1	99.0	.	DISC_MAPQ=28;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=411167_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_175199501_175224501_362C;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:64 GQ:24 PL:[264.0, 24.0, 0.0] SR:55 DR:50 LR:-264.1 LO:264.1);ALT=A]chr1:175201937];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	182274475	+	chr17	74319261	+	AAAAAAAAAAAA	38	25	435733_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=AAAAAAAAAAAA;MAPQ=60;MATEID=435733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_182255501_182280501_315C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:52 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:25 DR:38 LR:-155.1 LO:155.1);ALT=A[chr17:74319261[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	182357889	+	chr1	182360814	+	.	84	13	435488_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=435488_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_182353501_182378501_373C;SPAN=2925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:122 GQ:23.3 PL:[270.8, 0.0, 23.3] SR:13 DR:84 LR:-282.5 LO:282.5);ALT=G[chr1:182360814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183602343	+	chr1	183604752	+	.	62	0	439783_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=439783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:183602343(+)-1:183604752(-)__1_183603001_183628001D;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:89 GQ:35.3 PL:[180.5, 0.0, 35.3] SR:0 DR:62 LR:-186.1 LO:186.1);ALT=A[chr1:183604752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201181092	+	chr1	201179775	+	.	31	0	492236_1	69.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=492236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201179775(-)-1:201181092(+)__1_201169501_201194501D;SPAN=1317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:122 GQ:69.5 PL:[69.5, 0.0, 224.6] SR:0 DR:31 LR:-69.28 LO:73.96);ALT=]chr1:201181092]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	201459515	+	chr1	201476196	+	.	33	0	493183_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=493183_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201459515(+)-1:201476196(-)__1_201463501_201488501D;SPAN=16681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:43 GQ:5 PL:[97.4, 0.0, 5.0] SR:0 DR:33 LR:-101.9 LO:101.9);ALT=G[chr1:201476196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202920292	+	chr1	202927313	+	.	56	8	498953_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=498953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_202909001_202934001_304C;SPAN=7021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:109 GQ:99 PL:[165.2, 0.0, 99.2] SR:8 DR:56 LR:-166.1 LO:166.1);ALT=A[chr1:202927313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	203830843	+	chr19	5576940	-	.	86	0	6708348_1	99.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=6708348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:203830843(+)-19:5576940(+)__19_5561501_5586501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:47 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:0 DR:86 LR:-254.2 LO:254.2);ALT=T]chr19:5576940];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	203830843	+	chr9	6748969	-	.	35	0	4132425_1	99.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4132425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:203830843(+)-9:6748969(+)__9_6737501_6762501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:27 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:35 LR:-102.3 LO:102.3);ALT=T]chr9:6748969];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	221913157	+	chr1	221915340	+	.	32	0	561828_1	78.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=561828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:221913157(+)-1:221915340(-)__1_221896501_221921501D;SPAN=2183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:101 GQ:78.5 PL:[78.5, 0.0, 164.3] SR:0 DR:32 LR:-78.27 LO:80.03);ALT=A[chr1:221915340[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	225133672	+	chr1	225248642	+	.	49	0	574239_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=574239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:225133672(+)-1:225248642(-)__1_225228501_225253501D;SPAN=114970;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:20 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:49 LR:-145.2 LO:145.2);ALT=C[chr1:225248642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228270547	+	chr1	228284776	+	.	140	0	585393_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=585393_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228270547(+)-1:228284776(-)__1_228266501_228291501D;SPAN=14229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:78 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:0 DR:140 LR:-415.9 LO:415.9);ALT=T[chr1:228284776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228295620	+	chr1	228296902	+	.	35	0	585862_1	93.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=585862_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228295620(+)-1:228296902(-)__1_228291001_228316001D;SPAN=1282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:80 GQ:93.8 PL:[93.8, 0.0, 100.4] SR:0 DR:35 LR:-93.86 LO:93.87);ALT=T[chr1:228296902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228328065	+	chr1	228333211	+	.	50	15	585707_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=585707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_228315501_228340501_25C;SPAN=5146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:148 GQ:99 PL:[144.8, 0.0, 214.1] SR:15 DR:50 LR:-144.8 LO:145.5);ALT=G[chr1:228333211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228328100	+	chr1	228334539	+	.	56	0	585709_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=585709_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228328100(+)-1:228334539(-)__1_228315501_228340501D;SPAN=6439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:118 GQ:99 PL:[152.9, 0.0, 133.1] SR:0 DR:56 LR:-153.0 LO:153.0);ALT=G[chr1:228334539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	229812537	+	chr1	229820837	+	.	100	80	591106_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTGT;MAPQ=60;MATEID=591106_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_1_229810001_229835001_227C;SPAN=8300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:38 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:80 DR:100 LR:-435.7 LO:435.7);ALT=T[chr1:229820837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235291967	-	chrX	72443018	+	.	34	0	611479_1	77.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=611479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235291967(-)-23:72443018(-)__1_235273501_235298501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:130 GQ:77 PL:[77.0, 0.0, 238.7] SR:0 DR:34 LR:-77.01 LO:81.62);ALT=[chrX:72443018[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	235993764	+	chr1	236030139	+	.	58	0	614263_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=614263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235993764(+)-1:236030139(-)__1_235984001_236009001D;SPAN=36375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:45 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=C[chr1:236030139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	236549103	+	chr1	236551330	+	.	69	56	616486_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TAATAATTTGAAAGTTA;MAPQ=60;MATEID=616486_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_236547501_236572501_394C;SPAN=2227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:37 GQ:27 PL:[297.0, 27.0, 0.0] SR:56 DR:69 LR:-297.1 LO:297.1);ALT=A[chr1:236551330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246091389	+	chr1	246350042	+	.	37	0	649825_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=649825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:246091389(+)-1:246350042(-)__1_246347501_246372501D;SPAN=258653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:76 GQ:81.8 PL:[101.6, 0.0, 81.8] SR:0 DR:37 LR:-101.6 LO:101.6);ALT=A[chr1:246350042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246729965	+	chr1	246754812	+	.	99	23	651890_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=651890_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_246715001_246740001_455C;SPAN=24847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:73 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:23 DR:99 LR:-359.8 LO:359.8);ALT=G[chr1:246754812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	247850475	+	chr1	247856516	+	.	100	60	655719_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=GAAAAGAAAGATC;MAPQ=60;MATEID=655719_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_247842001_247867001_25C;SPAN=6041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:49 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:60 DR:100 LR:-389.5 LO:389.5);ALT=C[chr1:247856516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	248051492	+	chr1	248057639	+	.	111	60	656454_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCATGTATTTATTT;MAPQ=60;MATEID=656454_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_1_248038001_248063001_31C;SPAN=6147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:42 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:60 DR:111 LR:-406.0 LO:406.0);ALT=T[chr1:248057639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	265011	+	chr2	271865	+	.	79	11	660263_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTAA;MAPQ=60;MATEID=660263_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_245001_270001_312C;SPAN=6854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:55 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:11 DR:79 LR:-237.7 LO:237.7);ALT=A[chr2:271865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	4781310	+	chr2	4787357	+	.	79	37	671921_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAGATACTGCA;MAPQ=60;MATEID=671921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_4777501_4802501_273C;SPAN=6047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:106 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:37 DR:79 LR:-312.5 LO:312.5);ALT=A[chr2:4787357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26459896	+	chr2	26467411	+	.	64	0	725439_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=725439_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:26459896(+)-2:26467411(-)__2_26460001_26485001D;SPAN=7515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:54 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=G[chr2:26467411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27593578	+	chr2	27595487	+	.	35	0	728801_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27593578(+)-2:27595487(-)__2_27587001_27612001D;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:0 DR:35 LR:-91.97 LO:92.16);ALT=T[chr2:27595487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27651632	+	chr2	27656113	+	.	39	0	729136_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=729136_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27651632(+)-2:27656113(-)__2_27636001_27661001D;SPAN=4481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:76 GQ:75.2 PL:[108.2, 0.0, 75.2] SR:0 DR:39 LR:-108.4 LO:108.4);ALT=A[chr2:27656113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27995252	+	chr2	28002300	+	TTGCCAAGAGCAAGTCAAA	148	7	730465_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTGCCAAGAGCAAGTCAAA;MAPQ=60;MATEID=730465_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_27979001_28004001_56C;SPAN=7048;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:133 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:7 DR:148 LR:-448.9 LO:448.9);ALT=G[chr2:28002300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28113759	+	chr2	28117396	+	.	33	0	730591_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=730591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:28113759(+)-2:28117396(-)__2_28101501_28126501D;SPAN=3637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:86 GQ:85.7 PL:[85.7, 0.0, 122.0] SR:0 DR:33 LR:-85.63 LO:86.0);ALT=G[chr2:28117396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	30369956	+	chr2	30378726	+	.	82	0	736719_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=736719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:30369956(+)-2:30378726(-)__2_30355501_30380501D;SPAN=8770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:69 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=G[chr2:30378726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41238369	+	chr2	41250294	+	.	50	32	764464_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGA;MAPQ=60;MATEID=764464_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41233501_41258501_84C;SPAN=11925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:40 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:32 DR:50 LR:-204.7 LO:204.7);ALT=A[chr2:41250294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41775966	+	chr2	41781284	+	G	57	55	765669_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=765669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41772501_41797501_165C;SPAN=5318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:25 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:55 DR:57 LR:-267.4 LO:267.4);ALT=T[chr2:41781284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41973156	+	chr2	41975866	+	.	79	54	766256_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAACCTCACATGC;MAPQ=60;MATEID=766256_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41968501_41993501_127C;SPAN=2710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:46 GQ:27 PL:[297.0, 27.0, 0.0] SR:54 DR:79 LR:-297.1 LO:297.1);ALT=C[chr2:41975866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42052666	+	chr4	66413930	+	.	42	0	766432_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=766432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:42052666(+)-4:66413930(-)__2_42042001_42067001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:39 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=A[chr4:66413930[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	42346259	+	chr2	42347319	+	TGTA	32	20	767122_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTA;MAPQ=60;MATEID=767122_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_42336001_42361001_22C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:59 GQ:36.8 PL:[106.1, 0.0, 36.8] SR:20 DR:32 LR:-108.0 LO:108.0);ALT=C[chr2:42347319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42578554	+	chr2	42588232	+	.	62	0	767923_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=767923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:42578554(+)-2:42588232(-)__2_42581001_42606001D;SPAN=9678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:61 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:0 DR:62 LR:-181.5 LO:181.5);ALT=T[chr2:42588232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42580486	+	chr2	42588229	+	.	165	41	767924_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=767924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_42581001_42606001_294C;SPAN=7743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:59 GQ:46 PL:[505.0, 46.0, 0.0] SR:41 DR:165 LR:-505.0 LO:505.0);ALT=G[chr2:42588229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47389830	+	chr2	47403577	+	.	106	0	781617_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=781617_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:47389830(+)-2:47403577(-)__2_47383001_47408001D;SPAN=13747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:81 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=T[chr2:47403577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47403577	-	chr10	71923415	+	.	54	0	781682_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=781682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:47403577(-)-10:71923415(-)__2_47383001_47408001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:45 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=[chr10:71923415[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	48541953	+	chr2	48573339	+	.	40	7	784914_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=784914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48559001_48584001_122C;SPAN=31386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:65 GQ:32 PL:[124.4, 0.0, 32.0] SR:7 DR:40 LR:-127.2 LO:127.2);ALT=G[chr2:48573339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	48781852	+	chr2	48784868	+	.	60	37	785747_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAAGTGCAAAATTTTTT;MAPQ=60;MATEID=785747_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48779501_48804501_359C;SPAN=3016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:60 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:37 DR:60 LR:-217.9 LO:217.9);ALT=T[chr2:48784868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	48851192	+	chr2	48857953	+	.	49	45	785640_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=785640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48853001_48878001_52C;SPAN=6761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:22 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:45 DR:49 LR:-221.2 LO:221.2);ALT=A[chr2:48857953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	63816227	+	chr2	63821669	+	.	59	0	821676_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=821676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63816227(+)-2:63821669(-)__2_63822501_63847501D;SPAN=5442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:0 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=T[chr2:63821669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	68592526	+	chr2	68607458	+	.	96	19	834109_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=834109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_68600001_68625001_162C;SPAN=14932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:48 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:19 DR:96 LR:-300.4 LO:300.4);ALT=G[chr2:68607458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	69969349	+	chr2	70031662	+	.	34	0	837624_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=837624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:69969349(+)-2:70031662(-)__2_70021001_70046001D;SPAN=62313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:47 GQ:13.7 PL:[99.5, 0.0, 13.7] SR:0 DR:34 LR:-103.1 LO:103.1);ALT=C[chr2:70031662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70662448	+	chr2	70661187	+	.	50	0	840263_1	99.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=840263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70661187(-)-2:70662448(+)__2_70658001_70683001D;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:78 GQ:44.9 PL:[143.9, 0.0, 44.9] SR:0 DR:50 LR:-146.7 LO:146.7);ALT=]chr2:70662448]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	73461512	+	chr2	73466770	+	.	50	8	846958_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=846958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_73451001_73476001_311C;SPAN=5258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:108 GQ:99 PL:[145.7, 0.0, 116.0] SR:8 DR:50 LR:-145.9 LO:145.9);ALT=G[chr2:73466770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73461550	+	chr2	73467562	+	.	31	0	846961_1	77.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=846961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:73461550(+)-2:73467562(-)__2_73451001_73476001D;SPAN=6012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:93 GQ:77.3 PL:[77.3, 0.0, 146.6] SR:0 DR:31 LR:-77.14 LO:78.38);ALT=C[chr2:73467562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74154180	+	chr2	74173845	+	.	57	39	849414_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=849414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74137001_74162001_15C;SPAN=19665;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:63 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:39 DR:57 LR:-221.2 LO:221.2);ALT=G[chr2:74173845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	76526512	+	chr2	76528894	+	.	48	40	855560_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTTTTCCATGTTTT;MAPQ=60;MATEID=855560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_76513501_76538501_253C;SPAN=2382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:34 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:40 DR:48 LR:-221.2 LO:221.2);ALT=T[chr2:76528894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84670575	+	chr2	84686302	+	.	71	0	873023_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=873023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:84670575(+)-2:84686302(-)__2_84672001_84697001D;SPAN=15727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:40 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=A[chr2:84686302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84676876	+	chr2	84686297	+	.	35	10	873035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=873035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_84672001_84697001_74C;SPAN=9421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:67 GQ:61.1 PL:[100.7, 0.0, 61.1] SR:10 DR:35 LR:-101.2 LO:101.2);ALT=A[chr2:84686297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85629118	+	chr2	85637404	+	.	147	0	875683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=875683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85629118(+)-2:85637404(-)__2_85627501_85652501D;SPAN=8286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:85 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:0 DR:147 LR:-435.7 LO:435.7);ALT=A[chr2:85637404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85629142	+	chr2	85641105	+	.	42	0	875684_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=875684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85629142(+)-2:85641105(-)__2_85627501_85652501D;SPAN=11963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:97 GQ:99 PL:[112.4, 0.0, 122.3] SR:0 DR:42 LR:-112.4 LO:112.4);ALT=A[chr2:85641105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85804773	+	chr2	85806131	+	.	106	5	876458_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=876458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85799001_85824001_256C;SPAN=1358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:143 DP:268 GQ:99 PL:[399.5, 0.0, 250.9] SR:5 DR:106 LR:-401.2 LO:401.2);ALT=G[chr2:85806131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85804826	+	chr2	85808698	+	.	94	0	876460_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=876460_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85804826(+)-2:85808698(-)__2_85799001_85824001D;SPAN=3872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:161 GQ:99 PL:[266.9, 0.0, 121.7] SR:0 DR:94 LR:-269.5 LO:269.5);ALT=C[chr2:85808698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86756521	+	chr2	86790425	+	CCTTATTTGCCTGTCAACAACTCTCATTTCCTTTCTTATCTTCAATGACCACTCATTG	32	20	879231_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=CCTTATTTGCCTGTCAACAACTCTCATTTCCTTTCTTATCTTCAATGACCACTCATTG;MAPQ=60;MATEID=879231_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_86754501_86779501_183C;SPAN=33904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:20 DR:32 LR:-118.8 LO:118.8);ALT=C[chr2:86790425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	89029246	+	chr2	89032283	+	.	82	30	887260_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATATTAAAACTAAG;MAPQ=60;MATEID=887260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_89008501_89033501_104C;SPAN=3037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:99 DP:164 GQ:99 PL:[282.5, 0.0, 114.2] SR:30 DR:82 LR:-286.2 LO:286.2);ALT=G[chr2:89032283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	89850662	+	chr2	89853637	+	.	44	25	893566_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATTTGAGTCCATTCCATCCCACTCCATT;MAPQ=60;MATEID=893566_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_89841501_89866501_311C;SPAN=2975;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:138 GQ:99 PL:[177.2, 0.0, 157.4] SR:25 DR:44 LR:-177.2 LO:177.2);ALT=T[chr2:89853637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99343031	+	chr2	99347510	+	.	32	3	910762_1	97.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=910762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_99323001_99348001_166C;SPAN=4479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:55 GQ:34.7 PL:[97.4, 0.0, 34.7] SR:3 DR:32 LR:-98.87 LO:98.87);ALT=C[chr2:99347510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	118572439	+	chr2	118575019	+	.	36	34	962222_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=962222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_118555501_118580501_305C;SPAN=2580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:89 GQ:18.8 PL:[197.0, 0.0, 18.8] SR:34 DR:36 LR:-205.7 LO:205.7);ALT=G[chr2:118575019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	119653329	+	chr2	119659369	+	.	63	48	964901_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CGGCACTGGCTT;MAPQ=60;MATEID=964901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_119633501_119658501_153C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:28 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:48 DR:63 LR:-274.0 LO:274.0);ALT=T[chr2:119659369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120124668	+	chr2	120125759	+	.	63	0	965746_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=965746_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:120124668(+)-2:120125759(-)__2_120123501_120148501D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:97 GQ:53 PL:[181.7, 0.0, 53.0] SR:0 DR:63 LR:-185.5 LO:185.5);ALT=T[chr2:120125759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120418488	+	chr2	120417080	+	GGC	37	72	966609_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GGC;MAPQ=60;MATEID=966609_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_120417501_120442501_334C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:25 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:72 DR:37 LR:-260.8 LO:260.8);ALT=]chr2:120418488]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	126443251	+	chr2	126451832	+	.	95	53	981173_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAAC;MAPQ=60;MATEID=981173_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_126444501_126469501_206C;SPAN=8581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:13 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:53 DR:95 LR:-373.0 LO:373.0);ALT=C[chr2:126451832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	127674758	+	chr2	127677273	+	.	85	53	983779_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=983779_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_127669501_127694501_17C;SPAN=2515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:27 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:53 DR:85 LR:-343.3 LO:343.3);ALT=C[chr2:127677273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	128528625	+	chr2	128568654	+	.	33	0	986631_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=986631_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:128528625(+)-2:128568654(-)__2_128527001_128552001D;SPAN=40029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:33 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:0 DR:33 LR:-95.72 LO:95.72);ALT=C[chr2:128568654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	139046347	+	chr17	1303411	+	.	35	0	6282323_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6282323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:139046347(+)-17:1303411(-)__17_1298501_1323501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:56 GQ:34.4 PL:[100.4, 0.0, 34.4] SR:0 DR:35 LR:-102.1 LO:102.1);ALT=T[chr17:1303411[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	153572641	+	chr2	153573870	+	.	34	6	1047485_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1047485_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_153566001_153591001_334C;SPAN=1229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:75 GQ:72.2 PL:[108.5, 0.0, 72.2] SR:6 DR:34 LR:-108.8 LO:108.8);ALT=C[chr2:153573870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	155007024	+	chr2	167545932	-	.	36	0	1079414_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=1079414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:155007024(+)-2:167545932(+)__2_167531001_167556001D;SPAN=12538908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:10 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=T]chr2:167545932];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	167545960	+	chr2	167547086	+	.	31	0	1079442_1	89.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=1079442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:167545960(+)-2:167547086(-)__2_167531001_167556001D;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:16 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=T[chr2:167547086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170105133	+	chr2	170111163	+	.	51	21	1085145_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAACAGCAATGTTGA;MAPQ=60;MATEID=1085145_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_170103501_170128501_12C;SPAN=6030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:55 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:21 DR:51 LR:-171.6 LO:171.6);ALT=A[chr2:170111163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170641518	+	chr2	170643952	+	.	70	41	1086336_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=TCATTATTTTC;MAPQ=60;MATEID=1086336_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_170618001_170643001_86C;SPAN=2434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:31 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:41 DR:70 LR:-280.6 LO:280.6);ALT=C[chr2:170643952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170655507	+	chr2	170661981	+	.	36	0	1086235_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1086235_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170655507(+)-2:170661981(-)__2_170642501_170667501D;SPAN=6474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:79 GQ:94.1 PL:[97.4, 0.0, 94.1] SR:0 DR:36 LR:-97.44 LO:97.44);ALT=A[chr2:170661981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	173004263	+	chr2	173007481	+	.	85	36	1092750_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GTAGAGATGGGGTTT;MAPQ=60;MATEID=1092750_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172994501_173019501_230C;SPAN=3218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:25 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:36 DR:85 LR:-290.5 LO:290.5);ALT=T[chr2:173007481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	175094189	+	chr2	175113178	+	.	58	0	1098190_1	99.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=1098190_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:175094189(+)-2:175113178(-)__2_175101501_175126501D;SPAN=18989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:31 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=A[chr2:175113178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42504992	+	chr2	175113176	+	.	61	0	7311591_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7311591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:175113176(-)-22:42504992(+)__22_42483001_42508001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:66 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:0 DR:61 LR:-194.7 LO:194.7);ALT=]chr22:42504992]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	176044031	+	chr2	176046382	+	.	87	0	1100781_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1100781_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:176044031(+)-2:176046382(-)__2_176032501_176057501D;SPAN=2351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:210 GQ:99 PL:[230.3, 0.0, 279.8] SR:0 DR:87 LR:-230.3 LO:230.6);ALT=T[chr2:176046382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176044956	+	chr2	176046382	+	.	97	0	1100786_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1100786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:176044956(+)-2:176046382(-)__2_176032501_176057501D;SPAN=1426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:201 GQ:99 PL:[266.0, 0.0, 219.8] SR:0 DR:97 LR:-265.9 LO:265.9);ALT=T[chr2:176046382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	177265645	+	chr2	177272041	+	.	97	76	1103493_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATT;MAPQ=60;MATEID=1103493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_177257501_177282501_173C;SPAN=6396;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:39 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:76 DR:97 LR:-412.6 LO:412.6);ALT=T[chr2:177272041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187351185	+	chr2	187359960	+	.	59	72	1126341_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1126341_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_187327001_187352001_151C;SPAN=8775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:57 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:72 DR:59 LR:-283.9 LO:283.9);ALT=G[chr2:187359960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	194545044	+	chr14	65447291	+	TTTTTTTTTTATTTTTATTTTTTTTTTTTTTTT	43	47	5775820_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TTTTA;INSERTION=TTTTTTTTTTATTTTTATTTTTTTTTTTTTTTT;MAPQ=60;MATEID=5775820_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_65439501_65464501_193C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:36 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:47 DR:43 LR:-224.5 LO:224.5);ALT=A[chr14:65447291[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	194689502	+	chr2	194698766	+	.	60	50	1142905_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1142905_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_194677001_194702001_27C;SPAN=9264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:25 GQ:24 PL:[264.0, 24.0, 0.0] SR:50 DR:60 LR:-264.1 LO:264.1);ALT=G[chr2:194698766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198288700	+	chr2	198299696	+	.	37	12	1151306_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1151306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198278501_198303501_370C;SPAN=10996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:102 GQ:99 PL:[127.7, 0.0, 117.8] SR:12 DR:37 LR:-127.5 LO:127.5);ALT=T[chr2:198299696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198362139	+	chr2	198364504	+	.	39	0	1151938_1	88.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=1151938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198362139(+)-2:198364504(-)__2_198352001_198377001D;SPAN=2365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:149 GQ:88.4 PL:[88.4, 0.0, 273.2] SR:0 DR:39 LR:-88.37 LO:93.64);ALT=G[chr2:198364504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201676743	+	chr2	201680061	+	.	55	0	1159312_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1159312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201676743(+)-2:201680061(-)__2_201659501_201684501D;SPAN=3318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:77 GQ:25.4 PL:[160.7, 0.0, 25.4] SR:0 DR:55 LR:-166.2 LO:166.2);ALT=C[chr2:201680061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	202146658	+	chr2	202149441	+	.	79	50	1160930_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCAAATTCTT;MAPQ=60;MATEID=1160930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_202149501_202174501_306C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:7 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:50 DR:79 LR:-333.4 LO:333.4);ALT=T[chr2:202149441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135347363	+	chr2	203104274	+	.	66	0	3621391_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=3621391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:203104274(-)-7:135347363(+)__7_135338001_135363001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:98 GQ:46.1 PL:[191.3, 0.0, 46.1] SR:0 DR:66 LR:-196.2 LO:196.2);ALT=]chr7:135347363]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	203638956	+	chr4	89444837	+	.	33	0	2080293_1	89.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=2080293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:203638956(+)-4:89444837(-)__4_89425001_89450001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:71 GQ:80 PL:[89.9, 0.0, 80.0] SR:0 DR:33 LR:-89.71 LO:89.71);ALT=T[chr4:89444837[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	208474495	+	chr2	208476785	+	.	77	33	1177710_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGAAAACCTATTC;MAPQ=60;MATEID=1177710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_208470501_208495501_63C;SPAN=2290;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:35 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:33 DR:77 LR:-287.2 LO:287.2);ALT=C[chr2:208476785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209033773	+	chr17	19995679	-	.	39	0	6342394_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6342394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:209033773(+)-17:19995679(+)__17_19992001_20017001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:32 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:39 LR:-115.5 LO:115.5);ALT=T]chr17:19995679];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	209131139	+	chr2	209136232	+	.	34	20	1179659_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1179659_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_209132001_209157001_38C;SPAN=5093;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:52 GQ:2.6 PL:[121.4, 0.0, 2.6] SR:20 DR:34 LR:-127.7 LO:127.7);ALT=G[chr2:209136232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216974181	+	chr2	216977737	+	.	35	9	1198042_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=1198042_2;MATENM=0;NM=0;NUMPARTS=7;REPSEQ=GG;SCTG=c_2_216972001_216997001_267C;SPAN=3556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:103 GQ:99 PL:[110.9, 0.0, 137.3] SR:9 DR:35 LR:-110.7 LO:110.9);ALT=G[chr2:216977737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216974226	+	chr2	216981379	+	.	36	0	1198045_1	91.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1198045_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:216974226(+)-2:216981379(-)__2_216972001_216997001D;SPAN=7153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:102 GQ:91.4 PL:[91.4, 0.0, 154.1] SR:0 DR:36 LR:-91.2 LO:92.14);ALT=C[chr2:216981379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217089943	+	chr2	217092499	+	.	79	45	1198277_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GCCATGTGTTCTT;MAPQ=60;MATEID=1198277_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_2_217070001_217095001_328C;SPAN=2556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:322 GQ:99 PL:[249.7, 0.0, 530.3] SR:45 DR:79 LR:-249.5 LO:255.1);ALT=T[chr2:217092499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217955896	+	chr2	217957267	+	.	41	33	1200419_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTGG;MAPQ=60;MATEID=1200419_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_217952001_217977001_18C;SPAN=1371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:45 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:33 DR:41 LR:-184.8 LO:184.8);ALT=G[chr2:217957267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219082086	+	chr2	219093456	+	.	104	0	1203182_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1203182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219082086(+)-2:219093456(-)__2_219079001_219104001D;SPAN=11370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:104 DP:160 GQ:88.7 PL:[299.9, 0.0, 88.7] SR:0 DR:104 LR:-306.3 LO:306.3);ALT=C[chr2:219093456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	228258379	+	chr2	228241100	+	.	51	23	1227072_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CACTTT;MAPQ=60;MATEID=1227072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_228242001_228267001_31C;SPAN=17279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:40 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:23 DR:51 LR:-191.4 LO:191.4);ALT=]chr2:228258379]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	230877120	+	chr2	230879677	+	.	69	49	1233472_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCTG;MAPQ=60;MATEID=1233472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_230863501_230888501_111C;SPAN=2557;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:62 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:49 DR:69 LR:-270.7 LO:270.7);ALT=G[chr2:230879677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231729788	+	chr2	231738130	+	.	53	0	1235889_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1235889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231729788(+)-2:231738130(-)__2_231721001_231746001D;SPAN=8342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:92 GQ:71 PL:[150.2, 0.0, 71.0] SR:0 DR:53 LR:-151.5 LO:151.5);ALT=C[chr2:231738130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232326730	+	chr2	232329046	+	CTTCTCCACTGCTATCATCTTCTTCATCTTCTGACATTTCCTCATCTTCACTATCTTCTTCTACCTCCTTTGGAGGAGGAGCCATTTTCTTGGGGTCACCTTGATTTTTACCTG	49	162	1237734_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTTCTCCACTGCTATCATCTTCTTCATCTTCTGACATTTCCTCATCTTCACTATCTTCTTCTACCTCCTTTGGAGGAGGAGCCATTTTCTTGGGGTCACCTTGATTTTTACCTG;MAPQ=60;MATEID=1237734_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_232309001_232334001_332C;SPAN=2316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:181 DP:130 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:162 DR:49 LR:-534.7 LO:534.7);ALT=T[chr2:232329046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232328079	+	chr2	232329114	+	.	106	0	1237741_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1237741_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232328079(+)-2:232329114(-)__2_232309001_232334001D;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:99 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=A[chr2:232329114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	238875775	+	chr2	238881731	+	.	53	13	1255559_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=1255559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_238875001_238900001_298C;SPAN=5956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:54 GQ:15 PL:[165.0, 15.0, 0.0] SR:13 DR:53 LR:-165.0 LO:165.0);ALT=G[chr2:238881731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9834882	+	chr3	9841864	+	.	57	0	1281018_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1281018_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:9834882(+)-3:9841864(-)__3_9824501_9849501D;SPAN=6982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:90 GQ:54.8 PL:[163.7, 0.0, 54.8] SR:0 DR:57 LR:-166.8 LO:166.8);ALT=G[chr3:9841864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9839462	+	chr3	9841865	+	.	31	68	1281026_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TCAGG;MAPQ=60;MATEID=1281026_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_3_9824501_9849501_273C;SPAN=2403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:112 GQ:6.2 PL:[263.6, 0.0, 6.2] SR:68 DR:31 LR:-278.0 LO:278.0);ALT=G[chr3:9841865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10157503	+	chr3	10167309	+	.	72	83	1281931_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1281931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_10143001_10168001_182C;SPAN=9806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:109 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:83 DR:72 LR:-379.6 LO:379.6);ALT=G[chr3:10167309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10157541	+	chr3	10167951	+	.	71	0	1281932_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1281932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10157541(+)-3:10167951(-)__3_10143001_10168001D;SPAN=10410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:90 GQ:8.6 PL:[209.9, 0.0, 8.6] SR:0 DR:71 LR:-221.2 LO:221.2);ALT=G[chr3:10167951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10354465	+	chr3	10362729	+	.	32	0	1282488_1	87.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1282488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10354465(+)-3:10362729(-)__3_10339001_10364001D;SPAN=8264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:66 GQ:71.3 PL:[87.8, 0.0, 71.3] SR:0 DR:32 LR:-87.83 LO:87.83);ALT=T[chr3:10362729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10357149	+	chr3	10362730	+	.	34	0	1282492_1	97.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1282492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10357149(+)-3:10362730(-)__3_10339001_10364001D;SPAN=5581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:54 GQ:31.7 PL:[97.7, 0.0, 31.7] SR:0 DR:34 LR:-99.33 LO:99.33);ALT=T[chr3:10362730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	17914057	+	chr10	71993020	+	.	53	14	1294793_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TGAGGAAGACTCGGTACTCCAGGGAGAAGGG;MAPQ=42;MATEID=1294793_2;MATENM=0;NM=9;NUMPARTS=2;SCTG=c_3_17909501_17934501_217C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:32 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:14 DR:53 LR:-188.1 LO:188.1);ALT=G[chr10:71993020[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	23847580	+	chr3	23848726	+	.	41	4	1302368_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1302368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_23838501_23863501_262C;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:41 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:4 DR:41 LR:-125.4 LO:125.4);ALT=G[chr3:23848726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32433559	+	chr3	32483331	+	.	31	38	1338760_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1338760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32462501_32487501_398C;SPAN=49772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:67 GQ:8.3 PL:[153.5, 0.0, 8.3] SR:38 DR:31 LR:-161.2 LO:161.2);ALT=T[chr3:32483331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32806763	+	chr3	32808062	+	.	50	18	1340216_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=TTGCAGTGAGCCAAGAT;MAPQ=60;MATEID=1340216_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_32805501_32830501_315C;SPAN=1299;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:78 GQ:15.2 PL:[173.6, 0.0, 15.2] SR:18 DR:50 LR:-181.4 LO:181.4);ALT=T[chr3:32808062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	37449928	+	chr3	39676077	-	.	36	42	1356067_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGTGAGCCAAGATCATGCCACTACACTCCAGCCTG;MAPQ=60;MATEID=1356067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37436001_37461001_212C;SPAN=2226149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:44 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:42 DR:36 LR:-221.2 LO:221.2);ALT=G]chr3:39676077];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	37450057	-	chr3	39675868	+	.	46	0	1356068_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1356068_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:37450057(-)-3:39675868(-)__3_37436001_37461001D;SPAN=2225811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:60 GQ:10.1 PL:[135.5, 0.0, 10.1] SR:0 DR:46 LR:-142.0 LO:142.0);ALT=[chr3:39675868[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	40498968	+	chr12	63359104	+	.	92	9	5220782_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5220782_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_63357001_63382001_5C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:101 DP:1279 GQ:12.8 PL:[0.0, 12.8, 3132.0] SR:9 DR:92 LR:13.11 LO:185.0);ALT=G[chr12:63359104[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	41818076	+	chr3	41821494	+	.	43	24	1370814_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAGGTACAAAATG;MAPQ=60;MATEID=1370814_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_41821501_41846501_79C;SPAN=3418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:27 GQ:15 PL:[165.0, 15.0, 0.0] SR:24 DR:43 LR:-165.0 LO:165.0);ALT=G[chr3:41821494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42633146	+	chr3	42635913	+	.	40	0	1374140_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1374140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:42633146(+)-3:42635913(-)__3_42630001_42655001D;SPAN=2767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:110 GQ:99 PL:[102.2, 0.0, 164.9] SR:0 DR:40 LR:-102.2 LO:103.0);ALT=G[chr3:42635913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42838373	+	chr3	42840811	+	.	107	53	1374684_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGAATCTTATAACTTCC;MAPQ=60;MATEID=1374684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_42826001_42851001_299C;SPAN=2438;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:40 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:53 DR:107 LR:-452.2 LO:452.2);ALT=C[chr3:42840811[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	44740991	-	chr3	44742263	+	.	78	81	1381228_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCACTTTGGGA;MAPQ=60;MATEID=1381228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_251C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:101 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:81 DR:78 LR:-429.1 LO:429.1);ALT=[chr3:44742263[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	44741013	+	chr3	44742285	-	.	61	63	1381229_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TCCCAAAGTGCTGGGATTACAGG;MAPQ=60;MATEID=1381229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_127C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:105 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:63 DR:61 LR:-326.8 LO:326.8);ALT=A]chr3:44742285];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	47490669	+	chr3	47493441	+	.	78	40	1391327_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=1391327_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47481001_47506001_157C;SPAN=2772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:73 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:40 DR:78 LR:-283.9 LO:283.9);ALT=C[chr3:47493441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48511243	+	chr3	48514417	+	.	53	10	1396355_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=28;MATEID=1396355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48510001_48535001_18C;SPAN=3174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:130 GQ:99 PL:[162.8, 0.0, 152.9] SR:10 DR:53 LR:-162.9 LO:162.9);ALT=C[chr3:48514417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48643336	+	chr3	48647003	+	.	63	0	1396662_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1396662_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48643336(+)-3:48647003(-)__3_48632501_48657501D;SPAN=3667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:107 GQ:80 PL:[179.0, 0.0, 80.0] SR:0 DR:63 LR:-181.0 LO:181.0);ALT=G[chr3:48647003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49397817	+	chr3	49399928	+	.	33	46	1400882_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1400882_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_49392001_49417001_2C;SPAN=2111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:120 GQ:89.6 PL:[201.8, 0.0, 89.6] SR:46 DR:33 LR:-204.2 LO:204.2);ALT=T[chr3:49399928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49413026	+	chr3	49449253	+	.	134	51	1400982_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1400982_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49392001_49417001_476C;SPAN=36227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:142 DP:181 GQ:17.2 PL:[419.9, 0.0, 17.2] SR:51 DR:134 LR:-441.6 LO:441.6);ALT=T[chr3:49449253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52005866	+	chr3	52007978	+	.	97	0	1410901_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1410901_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52005866(+)-3:52007978(-)__3_51989001_52014001D;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:118 GQ:2.1 PL:[290.4, 2.1, 0.0] SR:0 DR:97 LR:-306.6 LO:306.6);ALT=G[chr3:52007978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52009220	+	chr3	52011886	+	.	42	12	1410917_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1410917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51989001_52014001_151C;SPAN=2666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:112 GQ:99 PL:[118.4, 0.0, 151.4] SR:12 DR:42 LR:-118.2 LO:118.5);ALT=G[chr3:52011886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52266194	+	chr3	52273015	+	.	105	0	1411874_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1411874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52266194(+)-3:52273015(-)__3_52258501_52283501D;SPAN=6821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:103 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:0 DR:105 LR:-310.3 LO:310.3);ALT=G[chr3:52273015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52269123	+	chr3	52273008	+	.	51	35	1411885_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1411885_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_52258501_52283501_34C;SPAN=3885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:94 GQ:67.1 PL:[159.5, 0.0, 67.1] SR:35 DR:51 LR:-161.3 LO:161.3);ALT=C[chr3:52273008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53275312	+	chr3	53289851	+	.	76	0	1416153_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1416153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53275312(+)-3:53289851(-)__3_53287501_53312501D;SPAN=14539;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:87 GQ:16.8 PL:[244.2, 16.8, 0.0] SR:0 DR:76 LR:-246.4 LO:246.4);ALT=T[chr3:53289851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53312247	+	chr3	53315559	+	.	41	37	1416276_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AAGTGATC;MAPQ=27;MATEID=1416276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53287501_53312501_18C;SPAN=3312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:29 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:37 DR:41 LR:-188.1 LO:188.1);ALT=C[chr3:53315559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57505598	+	chr3	141457288	-	.	56	0	1691813_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=1691813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:57505598(+)-3:141457288(+)__3_141438501_141463501D;SPAN=83951690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:76 GQ:19.1 PL:[164.3, 0.0, 19.1] SR:0 DR:56 LR:-170.8 LO:170.8);ALT=C]chr3:141457288];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	67493708	+	chr3	67496800	+	.	47	25	1463988_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAATTAGATCTC;MAPQ=60;MATEID=1463988_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_67473001_67498001_289C;SPAN=3092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:58 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:25 DR:47 LR:-178.2 LO:178.2);ALT=C[chr3:67496800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69134376	+	chr3	69150989	+	.	68	91	1469160_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=1469160_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_69114501_69139501_192C;SPAN=16613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:87 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:91 DR:68 LR:-406.0 LO:406.0);ALT=T[chr3:69150989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	95465768	+	chr3	95470764	+	.	53	45	1540653_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CAAG;MAPQ=60;MATEID=1540653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_95C;SPAN=4996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:104 GQ:8.1 PL:[267.3, 8.1, 0.0] SR:45 DR:53 LR:-276.8 LO:276.8);ALT=G[chr3:95470764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	95471000	+	chr3	95468117	+	TGCATAGGG	43	35	1540655_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGCATAGGG;MAPQ=60;MATEID=1540655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_267C;SPAN=2883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:97 GQ:72.8 PL:[161.9, 0.0, 72.8] SR:35 DR:43 LR:-163.7 LO:163.7);ALT=]chr3:95471000]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	98899063	+	chr3	98902390	+	.	43	29	1550958_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=1550958_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_98882001_98907001_475C;SPAN=3327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:57 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:29 DR:43 LR:-168.3 LO:168.3);ALT=T[chr3:98902390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	100053691	+	chr3	100058657	+	.	42	0	1554362_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1554362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:100053691(+)-3:100058657(-)__3_100058001_100083001D;SPAN=4966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:58 GQ:17.3 PL:[122.9, 0.0, 17.3] SR:0 DR:42 LR:-127.4 LO:127.4);ALT=G[chr3:100058657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	101293131	+	chr3	101298430	+	.	59	0	1558296_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1558296_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101293131(+)-3:101298430(-)__3_101283001_101308001D;SPAN=5299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:105 GQ:87.2 PL:[166.4, 0.0, 87.2] SR:0 DR:59 LR:-167.6 LO:167.6);ALT=C[chr3:101298430[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	101293152	+	chr13	48902558	-	.	41	0	5490003_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5490003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101293152(+)-13:48902558(+)__13_48877501_48902501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:18 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=C]chr13:48902558];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	42924510	+	chr3	101405405	+	.	38	0	2819974_1	67.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2819974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101405405(-)-6:42924510(+)__6_42899501_42924501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:213 GQ:67.9 PL:[67.9, 0.0, 447.5] SR:0 DR:38 LR:-67.73 LO:84.01);ALT=]chr6:42924510]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	120315385	+	chr3	120319956	+	.	36	0	1618392_1	86.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1618392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:120315385(+)-3:120319956(-)__3_120295001_120320001D;SPAN=4571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:121 GQ:86.3 PL:[86.3, 0.0, 205.1] SR:0 DR:36 LR:-86.05 LO:88.83);ALT=T[chr3:120319956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121366339	+	chr3	121379674	+	.	36	0	1621519_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1621519_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121366339(+)-3:121379674(-)__3_121373001_121398001D;SPAN=13335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:62 GQ:46.1 PL:[102.2, 0.0, 46.1] SR:0 DR:36 LR:-103.1 LO:103.1);ALT=T[chr3:121379674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121376246	+	chr3	121379670	+	.	63	0	1621541_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1621541_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121376246(+)-3:121379670(-)__3_121373001_121398001D;SPAN=3424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:115 GQ:99 PL:[176.9, 0.0, 101.0] SR:0 DR:63 LR:-177.9 LO:177.9);ALT=A[chr3:121379670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121377196	+	chr3	121379667	+	.	34	13	1621548_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1621548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121373001_121398001_176C;SPAN=2471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:127 GQ:84.5 PL:[84.5, 0.0, 223.1] SR:13 DR:34 LR:-84.43 LO:87.92);ALT=T[chr3:121379667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121554238	+	chr3	121563300	+	.	39	39	1622097_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=1622097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121544501_121569501_65C;SPAN=9062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:110 GQ:99 PL:[148.4, 0.0, 118.7] SR:39 DR:39 LR:-148.6 LO:148.6);ALT=T[chr3:121563300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122044207	+	chr3	122056392	+	.	33	30	1623628_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1623628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122034501_122059501_147C;SPAN=12185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:113 GQ:99 PL:[134.6, 0.0, 137.9] SR:30 DR:33 LR:-134.4 LO:134.4);ALT=T[chr3:122056392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122044235	+	chr3	122060281	+	.	71	0	1623683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1623683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:122044235(+)-3:122060281(-)__3_122059001_122084001D;SPAN=16046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:55 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=G[chr3:122060281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122103147	+	chr3	122121605	+	.	53	10	1623847_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1623847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122108001_122133001_270C;SPAN=18458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:56 GQ:15 PL:[165.0, 15.0, 0.0] SR:10 DR:53 LR:-165.0 LO:165.0);ALT=G[chr3:122121605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122103185	+	chr3	122123104	+	.	32	0	1623849_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1623849_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:122103185(+)-3:122123104(-)__3_122108001_122133001D;SPAN=19919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:51 GQ:29.3 PL:[92.0, 0.0, 29.3] SR:0 DR:32 LR:-93.4 LO:93.4);ALT=G[chr3:122123104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127540682	+	chr3	127541926	+	.	43	21	1643512_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1643512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127522501_127547501_87C;SPAN=1244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:113 GQ:99 PL:[131.3, 0.0, 141.2] SR:21 DR:43 LR:-131.1 LO:131.2);ALT=C[chr3:127541926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128445118	+	chr3	128514201	+	.	49	0	1646917_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1646917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:128445118(+)-3:128514201(-)__3_128502501_128527501D;SPAN=69083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:66 GQ:15.2 PL:[143.9, 0.0, 15.2] SR:0 DR:49 LR:-149.8 LO:149.8);ALT=C[chr3:128514201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128890617	+	chr3	128902619	+	.	255	26	1648624_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=1648624_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128870001_128895001_315C;SPAN=12002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:258 DP:72 GQ:69.7 PL:[765.7, 69.7, 0.0] SR:26 DR:255 LR:-765.8 LO:765.8);ALT=T[chr3:128902619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	129763382	+	chr3	129806746	+	.	64	34	1652305_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=1652305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_129801001_129826001_158C;SPAN=43364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:39 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:34 DR:64 LR:-237.7 LO:237.7);ALT=C[chr3:129806746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	143219592	+	chr3	143221217	+	.	40	35	1698113_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATGTTA;MAPQ=60;MATEID=1698113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_143202501_143227501_296C;SPAN=1625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:56 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:35 DR:40 LR:-181.5 LO:181.5);ALT=A[chr3:143221217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	148709434	+	chr3	148711927	+	.	32	12	1714640_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1714640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148690501_148715501_306C;SPAN=2493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:112 GQ:92 PL:[92.0, 0.0, 177.8] SR:12 DR:32 LR:-91.79 LO:93.37);ALT=G[chr3:148711927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150264665	+	chr3	150280328	+	.	45	0	1720105_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1720105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150264665(+)-3:150280328(-)__3_150258501_150283501D;SPAN=15663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:93 GQ:99 PL:[123.5, 0.0, 100.4] SR:0 DR:45 LR:-123.5 LO:123.5);ALT=T[chr3:150280328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	151962215	+	chr3	152017192	+	TAAAGCATAG	54	7	1726448_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TAAAGCATAG;MAPQ=60;MATEID=1726448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_151998001_152023001_33C;SPAN=54977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:80 GQ:24.5 PL:[169.7, 0.0, 24.5] SR:7 DR:54 LR:-176.0 LO:176.0);ALT=T[chr3:152017192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	152311738	+	chr3	152313156	+	.	75	42	1727140_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAGGTCACTGTTT;MAPQ=60;MATEID=1727140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_152292001_152317001_39C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:96 DP:235 GQ:99 PL:[253.4, 0.0, 316.1] SR:42 DR:75 LR:-253.2 LO:253.6);ALT=T[chr3:152313156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	158350740	+	chr3	158351912	+	.	60	35	1746939_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1746939_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_158343501_158368501_258C;SPAN=1172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:68 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:35 DR:60 LR:-217.9 LO:217.9);ALT=C[chr3:158351912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	163919285	+	chr10	36760446	+	.	50	39	4574086_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=4574086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_36750001_36775001_210C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:38 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:50 LR:-201.3 LO:201.3);ALT=A[chr10:36760446[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	169684685	+	chr3	169694728	+	.	35	0	1781870_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1781870_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:169684685(+)-3:169694728(-)__3_169687001_169712001D;SPAN=10043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:57 GQ:37.4 PL:[100.1, 0.0, 37.4] SR:0 DR:35 LR:-101.6 LO:101.6);ALT=C[chr3:169694728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	170586204	+	chr3	170587947	+	.	54	0	1784532_1	99.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1784532_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:170586204(+)-3:170587947(-)__3_170569001_170594001D;SPAN=1743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:149 GQ:99 PL:[137.9, 0.0, 223.7] SR:0 DR:54 LR:-137.9 LO:139.0);ALT=T[chr3:170587947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179320586	+	chr3	179322313	+	.	39	9	1813245_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1813245_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179315501_179340501_263C;SPAN=1727;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:109 GQ:99 PL:[102.5, 0.0, 161.9] SR:9 DR:39 LR:-102.5 LO:103.2);ALT=C[chr3:179322313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179322727	+	chr3	179332758	+	.	58	44	1813256_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1813256_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GTCGTC;SCTG=c_3_179315501_179340501_325C;SPAN=10031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:103 DP:136 GQ:12.8 PL:[231.3, 0.0, 12.8] SR:44 DR:58 LR:-244.7 LO:244.7);ALT=G[chr3:179332758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	180707414	-	chr14	45759196	+	.	36	0	5726304_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5726304_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:180707414(-)-14:45759196(-)__14_45741501_45766501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:51 GQ:16.1 PL:[105.2, 0.0, 16.1] SR:0 DR:36 LR:-108.4 LO:108.4);ALT=[chr14:45759196[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	183585850	+	chr3	183602508	+	.	52	27	1828389_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=1828389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183578501_183603501_240C;SPAN=16658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:130 GQ:99 PL:[176.0, 0.0, 139.7] SR:27 DR:52 LR:-176.3 LO:176.3);ALT=T[chr3:183602508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183892749	+	chr3	183894737	+	.	60	13	1828920_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1828920_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183872501_183897501_12C;SPAN=1988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:136 GQ:99 PL:[177.8, 0.0, 151.4] SR:13 DR:60 LR:-177.8 LO:177.8);ALT=T[chr3:183894737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183892781	+	chr3	183896641	+	.	60	0	1828921_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1828921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:183892781(+)-3:183896641(-)__3_183872501_183897501D;SPAN=3860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:128 GQ:99 PL:[163.4, 0.0, 146.9] SR:0 DR:60 LR:-163.4 LO:163.4);ALT=A[chr3:183896641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184081353	+	chr3	184082752	+	.	43	20	1829901_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1829901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_184068501_184093501_123C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:118 GQ:99 PL:[133.1, 0.0, 152.9] SR:20 DR:43 LR:-133.1 LO:133.2);ALT=G[chr3:184082752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186501450	+	chrX	52862812	-	.	41	0	7424856_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7424856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186501450(+)-23:52862812(+)__23_52846501_52871501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:28 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=G]chrX:52862812];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	186581033	+	chr3	186585285	+	.	75	42	1839808_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GAAAAATATTGCAAATAG;MAPQ=60;MATEID=1839808_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_186567501_186592501_262C;SPAN=4252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:85 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:42 DR:75 LR:-293.8 LO:293.8);ALT=G[chr3:186585285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	192875332	+	chr3	192885406	+	.	46	38	1860239_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TCT;MAPQ=60;MATEID=1860239_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_192864001_192889001_30C;SPAN=10074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:70 GQ:15.6 PL:[201.3, 15.6, 0.0] SR:38 DR:46 LR:-202.4 LO:202.4);ALT=T[chr3:192885406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	194546431	+	chr3	194543310	+	.	78	92	1866318_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1866318_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_194530001_194555001_83C;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:99 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:92 DR:78 LR:-429.1 LO:429.1);ALT=]chr3:194546431]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	196366747	+	chr3	196381398	+	.	45	13	1875112_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1875112_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_196343001_196368001_446C;SPAN=14651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:48 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:13 DR:45 LR:-145.2 LO:145.2);ALT=G[chr3:196381398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196467029	+	chr3	196509496	+	.	50	58	1875735_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1875735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196465501_196490501_162C;SPAN=42467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:70 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:58 DR:50 LR:-250.9 LO:250.9);ALT=G[chr3:196509496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196934573	+	chr3	196939256	+	CAGACT	56	38	1877108_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CAGACT;MAPQ=60;MATEID=1877108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196931001_196956001_77C;SPAN=4683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:70 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:38 DR:56 LR:-217.9 LO:217.9);ALT=A[chr3:196939256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197843929	+	chr3	197850167	+	.	92	79	1881562_1	99.0	.	DISC_MAPQ=25;EVDNC=ASDIS;HOMSEQ=GGC;MAPQ=60;MATEID=1881562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_197837501_197862501_505C;SPAN=6238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:36 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:79 DR:92 LR:-425.8 LO:425.8);ALT=C[chr3:197850167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	666358	+	chr4	667998	+	.	48	0	1883237_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1883237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:666358(+)-4:667998(-)__4_661501_686501D;SPAN=1640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:164 GQ:99 PL:[114.2, 0.0, 282.5] SR:0 DR:48 LR:-114.0 LO:118.0);ALT=T[chr4:667998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1267490	+	chr4	1266053	+	.	37	0	1885387_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=1885387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1266053(-)-4:1267490(+)__4_1249501_1274501D;SPAN=1437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:71 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.2 LO:103.2);ALT=]chr4:1267490]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	6651593	+	chr4	6652911	+	.	63	47	1895414_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CAGA;MAPQ=60;MATEID=1895414_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_6639501_6664501_271C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:24 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:47 DR:63 LR:-270.7 LO:270.7);ALT=A[chr4:6652911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	7995809	+	chr4	7996894	+	.	63	32	1898035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGGAAGCATTCTT;MAPQ=60;MATEID=1898035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_7987001_8012001_254C;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:104 GQ:8.3 PL:[242.6, 0.0, 8.3] SR:32 DR:63 LR:-255.4 LO:255.4);ALT=T[chr4:7996894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	10105658	+	chr4	10118307	+	.	32	0	1902634_1	94.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1902634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:10105658(+)-4:10118307(-)__4_10094001_10119001D;SPAN=12649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:42 GQ:5.3 PL:[94.4, 0.0, 5.3] SR:0 DR:32 LR:-98.59 LO:98.59);ALT=A[chr4:10118307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	10211267	+	chr4	10234568	+	.	65	49	1902852_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTTTCAA;MAPQ=60;MATEID=1902852_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_10192001_10217001_168C;SPAN=23301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:12 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:49 DR:65 LR:-267.4 LO:267.4);ALT=A[chr4:10234568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	17579208	+	chr6	36641580	+	.	43	0	1913378_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1913378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:17579208(+)-6:36641580(-)__4_17566501_17591501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:23 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=G[chr6:36641580[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	18420151	+	chr12	131712545	-	.	33	0	5397687_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5397687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:18420151(+)-12:131712545(+)__12_131712001_131737001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:33 LR:-102.3 LO:102.3);ALT=G]chr12:131712545];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	71523073	+	chr4	71532143	+	.	71	0	2022425_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=2022425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:71523073(+)-4:71532143(-)__4_71515501_71540501D;SPAN=9070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:98 GQ:29.6 PL:[207.8, 0.0, 29.6] SR:0 DR:71 LR:-215.5 LO:215.5);ALT=G[chr4:71532143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71527935	+	chr4	71532144	+	.	94	21	2022439_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=2022439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_71515501_71540501_247C;SPAN=4209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:112 GQ:30 PL:[330.0, 30.0, 0.0] SR:21 DR:94 LR:-330.1 LO:330.1);ALT=T[chr4:71532144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	75023999	+	chr4	75025770	+	.	34	25	2033312_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2033312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_75019001_75044001_219C;SPAN=1771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:135 GQ:99 PL:[115.4, 0.0, 211.1] SR:25 DR:34 LR:-115.3 LO:116.8);ALT=G[chr4:75025770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	79269134	+	chr4	79275196	+	.	56	15	2047479_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAGCTTCAAGATA;MAPQ=60;MATEID=2047479_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_79257501_79282501_431C;SPAN=6062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:199 GQ:99 PL:[154.1, 0.0, 329.0] SR:15 DR:56 LR:-154.1 LO:157.5);ALT=A[chr4:79275196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83196114	-	chr12	51717804	+	.	54	4	2059126_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=ACCTTCTCCTGGGCCCTGCT;MAPQ=43;MATEID=2059126_2;MATENM=0;NM=7;NUMPARTS=2;SCTG=c_4_83177501_83202501_264C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:57 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:4 DR:54 LR:-171.6 LO:171.6);ALT=[chr12:51717804[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	83616163	+	chr5	134263298	+	AAC	33	18	2060658_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AAC;MAPQ=60;MATEID=2060658_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_83594001_83619001_229C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:58 GQ:0.8 PL:[139.4, 0.0, 0.8] SR:18 DR:33 LR:-147.8 LO:147.8);ALT=C[chr5:134263298[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	84026199	+	chr4	84035817	+	.	50	0	2062620_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=2062620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84026199(+)-4:84035817(-)__4_84035001_84060001D;SPAN=9618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:50 LR:-161.7 LO:161.7);ALT=T[chr4:84035817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84029103	+	chr4	84035819	+	.	84	10	2062621_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;MAPQ=60;MATEID=2062621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_84035001_84060001_125C;SPAN=6716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:61 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:10 DR:84 LR:-250.9 LO:250.9);ALT=A[chr4:84035819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	132611296	+	chr4	84035816	+	.	65	0	5400324_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5400324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84035816(-)-12:132611296(+)__12_132594001_132619001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:36 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=]chr12:132611296]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	88303516	+	chr4	88312013	+	.	35	67	2076300_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2076300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_88298001_88323001_247C;SPAN=8497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:127 GQ:87.8 PL:[219.8, 0.0, 87.8] SR:67 DR:35 LR:-222.8 LO:222.8);ALT=T[chr4:88312013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88483900	+	chr4	88486313	+	.	88	56	2077334_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAGTTACAAACAAC;MAPQ=60;MATEID=2077334_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_88469501_88494501_334C;SPAN=2413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:51 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:56 DR:88 LR:-340.0 LO:340.0);ALT=C[chr4:88486313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88847164	-	chr4	88858700	+	A	115	69	2078496_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=2078496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_88837001_88862001_254C;SPAN=11536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:68 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:69 DR:115 LR:-458.8 LO:458.8);ALT=[chr4:88858700[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	94559454	+	chr4	94565491	+	.	107	64	2094967_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAAAACTTGCATCTT;MAPQ=60;MATEID=2094967_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_94545501_94570501_233C;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:46 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:64 DR:107 LR:-399.4 LO:399.4);ALT=T[chr4:94565491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	95518746	+	chr7	46904659	+	.	95	84	3290388_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAGCC;MAPQ=60;MATEID=3290388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_46893001_46918001_396C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:45 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:84 DR:95 LR:-432.4 LO:432.4);ALT=C[chr7:46904659[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	5273545	+	chr4	103748338	+	.	57	0	2122682_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2122682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:103748338(-)-20:5273545(+)__4_103733001_103758001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:93 GQ:60.8 PL:[163.1, 0.0, 60.8] SR:0 DR:57 LR:-165.4 LO:165.4);ALT=]chr20:5273545]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	107056578	+	chr4	107063363	+	CA	32	33	2132529_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CA;MAPQ=60;MATEID=2132529_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_107040501_107065501_326C;SPAN=6785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:51 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:33 DR:32 LR:-148.5 LO:148.5);ALT=C[chr4:107063363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107237794	+	chr4	107248607	+	.	42	0	2133059_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2133059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107237794(+)-4:107248607(-)__4_107236501_107261501D;SPAN=10813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:105 GQ:99 PL:[110.3, 0.0, 143.3] SR:0 DR:42 LR:-110.2 LO:110.5);ALT=T[chr4:107248607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108127828	+	chr4	108131715	+	.	93	61	2135501_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAACATTAGGATTCTCTTT;MAPQ=60;MATEID=2135501_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108118501_108143501_113C;SPAN=3887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:127 DP:34 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:61 DR:93 LR:-376.3 LO:376.3);ALT=T[chr4:108131715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108276701	+	chr4	108279505	+	.	61	66	2135779_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAC;MAPQ=60;MATEID=2135779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108265501_108290501_170C;SPAN=2804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:41 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:66 DR:61 LR:-310.3 LO:310.3);ALT=C[chr4:108279505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115507821	+	chr4	115513865	+	TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT	33	61	2158821_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT;MAPQ=60;MATEID=2158821_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_115493001_115518001_217C;SPAN=6044;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:66 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:61 DR:33 LR:-241.0 LO:241.0);ALT=G[chr4:115513865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115928723	+	chr4	115931874	+	.	48	36	2160360_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTGA;MAPQ=60;MATEID=2160360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_115909501_115934501_351C;SPAN=3151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:61 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:36 DR:48 LR:-201.3 LO:201.3);ALT=A[chr4:115931874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	130961892	+	chr4	131004550	+	CCT	60	55	2206992_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCT;MAPQ=60;MATEID=2206992_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_131001501_131026501_192C;SPAN=42658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:48 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:55 DR:60 LR:-274.0 LO:274.0);ALT=C[chr4:131004550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	138966211	+	chr4	138967219	+	T	49	30	2231112_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=2231112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_138964001_138989001_336C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:63 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:30 DR:49 LR:-184.8 LO:184.8);ALT=G[chr4:138967219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140587233	+	chr4	140599697	+	.	35	49	2236749_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=2236749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_140581001_140606001_221C;SPAN=12464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:131 GQ:99 PL:[189.2, 0.0, 126.5] SR:49 DR:35 LR:-189.6 LO:189.6);ALT=T[chr4:140599697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	142230783	+	chr4	142233063	+	.	112	70	2241959_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGCC;MAPQ=60;MATEID=2241959_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_142222501_142247501_77C;SPAN=2280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:38 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:70 DR:112 LR:-445.6 LO:445.6);ALT=C[chr4:142233063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	146919581	+	chr4	146927741	+	.	46	28	2256404_1	99.0	.	DISC_MAPQ=14;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=0;MATEID=2256404_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_4_146926501_146951501_360C;SECONDARY;SPAN=8160;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:36 GQ:18 PL:[198.0, 18.0, 0.0] SR:28 DR:46 LR:-198.0 LO:198.0);ALT=T[chr4:146927741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147208406	+	chr4	147206794	+	.	91	0	2257297_1	99.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=2257297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:147206794(-)-4:147208406(+)__4_147196001_147221001D;SPAN=1612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:101 GQ:27 PL:[297.0, 27.0, 0.0] SR:0 DR:91 LR:-297.1 LO:297.1);ALT=]chr4:147208406]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1043012	+	chr5	1041007	+	.	50	0	2400174_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2400174_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:1041007(-)-5:1043012(+)__5_1029001_1054001D;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:42 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=]chr5:1043012]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1178294	+	chr5	1180733	+	.	51	30	2400027_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=2400027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_1176001_1201001_111C;SPAN=2439;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:15 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:30 DR:51 LR:-211.3 LO:211.3);ALT=T[chr5:1180733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	1801690	+	chr5	1814450	+	.	84	0	2401318_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2401318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:1801690(+)-5:1814450(-)__5_1813001_1838001D;SPAN=12760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:67 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=C[chr5:1814450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32585763	+	chr5	32591666	+	.	79	0	2446915_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2446915_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:32585763(+)-5:32591666(-)__5_32585001_32610001D;SPAN=5903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:70 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=T[chr5:32591666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76145980	+	chr5	76166020	+	.	63	6	2507680_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2507680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_76146001_76171001_250C;SPAN=20040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:60 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:6 DR:63 LR:-194.7 LO:194.7);ALT=G[chr5:76166020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76146022	+	chr5	76171125	+	.	50	0	2507682_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2507682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:76146022(+)-5:76171125(-)__5_76146001_76171001D;SPAN=25103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:20 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=A[chr5:76171125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	81572339	+	chr5	81574137	+	.	60	0	2516215_1	0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2516215_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:81572339(+)-5:81574137(-)__5_81560501_81585501D;SPAN=1798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:60 DP:1079 GQ:94 PL:[0.0, 94.0, 2809.0] SR:0 DR:60 LR:94.27 LO:100.5);ALT=T[chr5:81574137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108230344	+	chr6	31774531	+	.	85	0	2775157_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=2775157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:108230344(+)-6:31774531(-)__6_31752001_31777001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:77 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:0 DR:85 LR:-250.9 LO:250.9);ALT=T[chr6:31774531[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	108595089	+	chr5	108601122	+	.	63	36	2550904_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAAATAAGAATGG;MAPQ=60;MATEID=2550904_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_108584001_108609001_141C;SPAN=6033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:40 GQ:21 PL:[231.0, 21.0, 0.0] SR:36 DR:63 LR:-231.1 LO:231.1);ALT=G[chr5:108601122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	112197123	+	chr18	56835763	+	.	40	0	6640949_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6640949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:112197123(+)-18:56835763(-)__18_56815501_56840501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:40 LR:-130.9 LO:130.9);ALT=T[chr18:56835763[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	131746735	+	chr5	131755513	+	.	34	11	2582387_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2582387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_131736501_131761501_94C;SPAN=8778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:70 GQ:63.5 PL:[106.4, 0.0, 63.5] SR:11 DR:34 LR:-107.1 LO:107.1);ALT=T[chr5:131755513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131825177	+	chr5	131826237	+	.	39	48	2582587_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2582587_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TGCTGC;SCTG=c_5_131810001_131835001_214C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:69 GQ:18.5 PL:[161.2, 18.5, 0.0] SR:48 DR:39 LR:-161.3 LO:161.3);ALT=T[chr5:131826237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133134710	+	chr5	133136486	+	.	51	0	2584716_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2584716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133134710(+)-5:133136486(-)__5_133133001_133158001D;SPAN=1776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:10 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:51 LR:-148.5 LO:148.5);ALT=A[chr5:133136486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49397979	+	chr5	133340188	+	.	98	0	7419751_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7419751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133340188(-)-23:49397979(+)__23_49392001_49417001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:36 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:0 DR:98 LR:-290.5 LO:290.5);ALT=]chrX:49397979]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	133496836	+	chr5	133512576	+	.	39	0	2585645_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2585645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133496836(+)-5:133512576(-)__5_133500501_133525501D;SPAN=15740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:98 GQ:99 PL:[102.2, 0.0, 135.2] SR:0 DR:39 LR:-102.2 LO:102.4);ALT=G[chr5:133512576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133509713	+	chr5	133512546	+	.	61	43	2585664_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;MAPQ=20;MATEID=2585664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133500501_133525501_277C;SPAN=2833;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:63 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:43 DR:61 LR:-270.7 LO:270.7);ALT=T[chr5:133512546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134094645	+	chr5	134099593	+	.	79	53	2586727_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2586727_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_134088501_134113501_116C;SPAN=4948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:86 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:53 DR:79 LR:-307.0 LO:307.0);ALT=G[chr5:134099593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134724816	+	chr5	134734752	+	.	135	30	2587827_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=2587827_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134725501_134750501_2C;SPAN=9936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:165 DP:47 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:30 DR:135 LR:-488.5 LO:488.5);ALT=A[chr5:134734752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	136854719	+	chr5	136856379	+	.	58	0	2590927_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2590927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:136854719(+)-5:136856379(-)__5_136857001_136882001D;SPAN=1660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:0 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=T[chr5:136856379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138677671	+	chr5	138699447	+	.	99	31	2594459_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2594459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138694501_138719501_118C;SPAN=21776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:42 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:31 DR:99 LR:-343.3 LO:343.3);ALT=T[chr5:138699447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140025311	+	chr5	140026841	+	.	40	3	2596901_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2596901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_140017501_140042501_157C;SPAN=1530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:85 GQ:89.3 PL:[115.7, 0.0, 89.3] SR:3 DR:40 LR:-115.8 LO:115.8);ALT=C[chr5:140026841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140080115	+	chr5	140081588	+	.	53	0	2596835_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2596835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140080115(+)-5:140081588(-)__5_140066501_140091501D;SPAN=1473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:65 GQ:0.9 PL:[158.4, 0.9, 0.0] SR:0 DR:53 LR:-167.0 LO:167.0);ALT=A[chr5:140081588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176258026	+	chr5	176259412	+	AAGTTC	59	57	2652125_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=AAGTTC;MAPQ=60;MATEID=2652125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176253001_176278001_254C;SPAN=1386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:31 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:57 DR:59 LR:-280.6 LO:280.6);ALT=A[chr5:176259412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176387587	+	chr5	176390181	+	.	44	27	2652209_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAAA;MAPQ=60;MATEID=2652209_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176375501_176400501_273C;SPAN=2594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:51 DP:725 GQ:27.7 PL:[0.0, 27.7, 1815.0] SR:27 DR:44 LR:28.07 LO:90.75);ALT=A[chr5:176390181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176785072	+	chr5	176793176	+	TCTGGCTGTGTCAGATGG	37	20	2653323_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCTGGCTGTGTCAGATGG;MAPQ=60;MATEID=2653323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176767501_176792501_208C;SPAN=8104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:38 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:20 DR:37 LR:-118.8 LO:118.8);ALT=T[chr5:176793176[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177580808	-	chr10	93976191	+	.	41	0	2654873_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2654873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:177580808(-)-10:93976191(-)__5_177576001_177601001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:74 GQ:62.6 PL:[115.4, 0.0, 62.6] SR:0 DR:41 LR:-116.1 LO:116.1);ALT=[chr10:93976191[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	179126103	+	chr5	179132678	+	.	68	14	2657864_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2657864_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_179119501_179144501_79C;SPAN=6575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:56 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:14 DR:68 LR:-208.0 LO:208.0);ALT=G[chr5:179132678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179221139	+	chr5	179222583	+	.	56	16	2658165_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2658165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179217501_179242501_156C;SPAN=1444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:50 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:16 DR:56 LR:-168.3 LO:168.3);ALT=G[chr5:179222583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179467649	+	chr5	179498456	+	.	38	52	2658587_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2658587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179487001_179512001_255C;SPAN=30807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:25 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:52 DR:38 LR:-217.9 LO:217.9);ALT=T[chr5:179498456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180668687	+	chr5	180670762	+	.	56	0	2660767_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2660767_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:180668687(+)-5:180670762(-)__5_180663001_180688001D;SPAN=2075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:492 GQ:51.8 PL:[51.8, 0.0, 1141.0] SR:0 DR:56 LR:-51.56 LO:111.9);ALT=T[chr5:180670762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180669347	+	chr5	180670692	+	.	127	131	2660770_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2660770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_180663001_180688001_277C;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:195 DP:604 GQ:99 PL:[480.3, 0.0, 985.3] SR:131 DR:127 LR:-480.1 LO:489.6);ALT=T[chr5:180670692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2834248	+	chr6	2836090	+	.	67	39	2670598_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2670598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2817501_2842501_366C;SPAN=1842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:130 GQ:67.1 PL:[248.6, 0.0, 67.1] SR:39 DR:67 LR:-254.5 LO:254.5);ALT=T[chr6:2836090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2838979	+	chr6	2842045	+	.	120	0	2670628_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2670628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2838979(+)-6:2842045(-)__6_2817501_2842501D;SPAN=3066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:120 DP:362 GQ:99 PL:[298.3, 0.0, 578.9] SR:0 DR:120 LR:-298.0 LO:303.0);ALT=C[chr6:2842045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2840854	+	chr6	2842043	+	.	136	0	2670639_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2670639_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2840854(+)-6:2842043(-)__6_2817501_2842501D;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:136 DP:333 GQ:99 PL:[358.9, 0.0, 448.0] SR:0 DR:136 LR:-358.7 LO:359.3);ALT=G[chr6:2842043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2959576	+	chr6	2971765	+	.	37	13	2671034_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=2671034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2964501_2989501_302C;SPAN=12189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:52 GQ:0.6 PL:[125.4, 0.6, 0.0] SR:13 DR:37 LR:-131.9 LO:131.9);ALT=C[chr6:2971765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6589103	+	chr6	6625158	+	.	72	60	2683742_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2683742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_6566001_6591001_182C;SPAN=36055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:74 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:60 DR:72 LR:-307.0 LO:307.0);ALT=G[chr6:6625158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6589120	+	chr6	6626525	+	.	46	0	2683744_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2683744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6589120(+)-6:6626525(-)__6_6566001_6591001D;SPAN=37405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:54 GQ:7.8 PL:[145.2, 7.8, 0.0] SR:0 DR:46 LR:-147.4 LO:147.4);ALT=C[chr6:6626525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7310308	+	chr6	7313328	+	.	43	0	2686608_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2686608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:7310308(+)-6:7313328(-)__6_7301001_7326001D;SPAN=3020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:99 GQ:99 PL:[115.1, 0.0, 125.0] SR:0 DR:43 LR:-115.1 LO:115.1);ALT=A[chr6:7313328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	8097702	+	chr6	8102668	+	.	38	8	2689588_1	58.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2689588_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCGCTCGC;SCTG=c_6_8085001_8110001_71C;SPAN=4966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:96 GQ:58.3 PL:[58.3, 0.0, 62.2] SR:8 DR:38 LR:-57.99 LO:58.02);ALT=T[chr6:8102668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723474	+	chr6	10724788	+	.	36	17	2698243_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2698243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_394C;SPAN=1314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:155 GQ:99 PL:[113.3, 0.0, 261.8] SR:17 DR:36 LR:-113.2 LO:116.4);ALT=G[chr6:10724788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723474	+	chr6	10725193	+	.	46	3	2698244_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2698244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_153C;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:180 GQ:99 PL:[113.0, 0.0, 324.2] SR:3 DR:46 LR:-113.0 LO:118.6);ALT=G[chr6:10725193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723511	+	chr6	10726136	+	.	32	0	2698248_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2698248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10723511(+)-6:10726136(-)__6_10706501_10731501D;SPAN=2625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:106 GQ:77 PL:[77.0, 0.0, 179.3] SR:0 DR:32 LR:-76.91 LO:79.21);ALT=C[chr6:10726136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10748157	+	chr10	70304647	-	.	111	0	4621447_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4621447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10748157(+)-10:70304647(+)__10_70290501_70315501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:37 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:111 LR:-326.8 LO:326.8);ALT=A]chr10:70304647];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	13191492	+	chr17	64637274	+	.	37	0	6472096_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6472096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:13191492(+)-17:64637274(-)__17_64631001_64656001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:47 GQ:3.8 PL:[109.4, 0.0, 3.8] SR:0 DR:37 LR:-115.2 LO:115.2);ALT=T[chr17:64637274[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	19765125	+	chr6	19771185	+	.	115	29	2731437_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGAAAAAAAAACTAACTGG;MAPQ=60;MATEID=2731437_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_19747001_19772001_100C;SECONDARY;SPAN=6060;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:131 DP:4255 GQ:99 PL:[0.0, 719.4, 11770.0] SR:29 DR:115 LR:720.4 LO:185.3);ALT=G[chr6:19771185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	27748738	+	chr15	55489062	+	.	61	0	5956060_1	99.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=5956060_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:27748738(+)-15:55489062(-)__15_55468001_55493001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:49 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:61 LR:-178.2 LO:178.2);ALT=C[chr15:55489062[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	29685488	+	chr6	29688081	+	.	105	24	2766515_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAGAAAGACCCAAGCCT;MAPQ=60;MATEID=2766515_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_29669501_29694501_51C;SPAN=2593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:112 DP:2059 GQ:99 PL:[0.0, 187.7, 5377.0] SR:24 DR:105 LR:188.1 LO:186.4);ALT=T[chr6:29688081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29814750	+	chr12	133088578	-	.	36	0	5401718_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5401718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29814750(+)-12:133088578(+)__12_133084001_133109001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:22 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=G]chr12:133088578];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	29899782	+	chr6	29901527	+	.	109	86	2767610_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=AAGAATTGAGGAGC;MAPQ=60;MATEID=2767610_2;MATENM=7;NM=1;NUMPARTS=2;SCTG=c_6_29890001_29915001_228C;SPAN=1745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:172 DP:37 GQ:46.3 PL:[508.3, 46.3, 0.0] SR:86 DR:109 LR:-508.3 LO:508.3);ALT=C[chr6:29901527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30585720	+	chr6	30587483	+	.	31	0	2769820_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2769820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30585720(+)-6:30587483(-)__6_30576001_30601001D;SPAN=1763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:108 GQ:73.1 PL:[73.1, 0.0, 188.6] SR:0 DR:31 LR:-73.07 LO:75.91);ALT=G[chr6:30587483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31211630	+	chr6	31213117	+	.	118	39	2772820_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AATACCCACCACCC;MAPQ=60;MATEID=2772820_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_31188501_31213501_461C;SPAN=1487;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:219 GQ:99 PL:[402.8, 0.0, 128.8] SR:39 DR:118 LR:-410.6 LO:410.6);ALT=C[chr6:31213117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31337861	+	chr6	31341967	+	.	34	34	2773094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCCA;MAPQ=60;MATEID=2773094_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_31335501_31360501_28C;SPAN=4106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:56 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:34 DR:34 LR:-178.2 LO:178.2);ALT=A[chr6:31341967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31555096	+	chr6	31556294	+	.	127	31	2773950_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2773950_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31531501_31556501_153C;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:148 DP:232 GQ:99 PL:[425.9, 0.0, 135.4] SR:31 DR:127 LR:-433.8 LO:433.8);ALT=G[chr6:31556294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31633994	+	chr6	31635642	+	.	86	0	2774553_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2774553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31633994(+)-6:31635642(-)__6_31629501_31654501D;SPAN=1648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:103 GQ:7.8 PL:[264.0, 7.8, 0.0] SR:0 DR:86 LR:-273.4 LO:273.4);ALT=G[chr6:31635642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31702042	+	chr6	31704038	+	.	166	17	2774836_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2774836_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31678501_31703501_77C;SPAN=1996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:74 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:17 DR:166 LR:-514.9 LO:514.9);ALT=T[chr6:31704038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31765887	+	chr6	31774529	+	.	32	0	2775239_1	74.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2775239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31765887(+)-6:31774529(-)__6_31752001_31777001D;SPAN=8642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:115 GQ:74.6 PL:[74.6, 0.0, 203.3] SR:0 DR:32 LR:-74.48 LO:77.84);ALT=T[chr6:31774529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31924828	+	chr6	31926667	+	.	59	0	2776166_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2776166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31924828(+)-6:31926667(-)__6_31923501_31948501D;SPAN=1839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:102 GQ:78.2 PL:[167.3, 0.0, 78.2] SR:0 DR:59 LR:-168.8 LO:168.8);ALT=G[chr6:31926667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32407809	+	chr6	32410223	+	.	162	94	2778079_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2778079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32389001_32414001_126C;SPAN=2414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:223 DP:621 GQ:99 PL:[568.2, 0.0, 937.9] SR:94 DR:162 LR:-567.9 LO:572.9);ALT=G[chr6:32410223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32487430	+	chr6	32489682	+	.	51	30	2779870_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2779870_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32487001_32512001_788C;SPAN=2252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:101 GQ:29 PL:[213.8, 0.0, 29.0] SR:30 DR:51 LR:-221.4 LO:221.4);ALT=T[chr6:32489682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32489951	+	chr6	32497902	+	.	147	77	2779892_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=2779892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32487001_32512001_80C;SPAN=7951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:175 DP:376 GQ:99 PL:[475.9, 0.0, 436.3] SR:77 DR:147 LR:-475.9 LO:475.9);ALT=G[chr6:32497902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32552155	+	chr6	32557420	+	.	162	48	2781961_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2781961_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32536001_32561001_813C;SPAN=5265;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:194 DP:324 GQ:99 PL:[552.8, 0.0, 232.6] SR:48 DR:162 LR:-559.7 LO:559.7);ALT=G[chr6:32557420[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32561965	+	chr6	32564609	+	.	88	68	2778886_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATTATTTTTC;MAPQ=60;MATEID=2778886_2;MATENM=0;NM=12;NUMPARTS=2;SCTG=c_6_32560501_32585501_315C;SPAN=2644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:39 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:68 DR:88 LR:-359.8 LO:359.8);ALT=C[chr6:32564609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32605317	+	chr6	32609086	+	.	119	57	2781019_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2781019_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32585001_32610001_973C;SPAN=3769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:183 GQ:13 PL:[468.7, 13.0, 0.0] SR:57 DR:119 LR:-486.7 LO:486.7);ALT=G[chr6:32609086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32719382	+	chr6	32620142	+	.	36	0	2779320_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2779320_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32620142(-)-6:32719382(+)__6_32609501_32634501D;SPAN=99240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:7 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=]chr6:32719382]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32623587	+	chr6	32624623	+	.	31	0	2779362_1	89.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2779362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32623587(+)-6:32624623(-)__6_32609501_32634501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:5 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=C[chr6:32624623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32632845	+	chr6	32634276	+	.	122	15	2778436_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=43;MATEID=2778436_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32634001_32659001_128C;SPAN=1431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:107 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:15 DR:122 LR:-402.7 LO:402.7);ALT=C[chr6:32634276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32778699	+	chr6	32779819	+	.	87	0	2780350_1	99.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2780350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32778699(+)-6:32779819(-)__6_32756501_32781501D;SPAN=1120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:28 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:0 DR:87 LR:-257.5 LO:257.5);ALT=C[chr6:32779819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32822066	+	chr6	32825039	+	ACCACCATCATGGCAGTGGAGTTTGACGGGGGCGTTGTGATGGGTTCTGATTCCCGAGTGTCTGCAG	90	93	2780593_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACCACCATCATGGCAGTGGAGTTTGACGGGGGCGTTGTGATGGGTTCTGATTCCCGAGTGTCTGCAG;MAPQ=60;MATEID=2780593_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32805501_32830501_416C;SPAN=2973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:124 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:93 DR:90 LR:-435.7 LO:435.7);ALT=G[chr6:32825039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32918582	+	chr6	32920726	+	.	151	38	2781158_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2781158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32903501_32928501_173C;SPAN=2144;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:164 DP:166 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:38 DR:151 LR:-491.8 LO:491.8);ALT=T[chr6:32920726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33037664	+	chr6	33041248	+	.	183	104	2782450_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2782450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_199C;SPAN=3584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:238 DP:410 GQ:99 PL:[674.5, 0.0, 321.4] SR:104 DR:183 LR:-681.4 LO:681.4);ALT=C[chr6:33041248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33043918	+	chr6	33048455	+	AGAATG	175	163	2782470_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AGAATG;MAPQ=60;MATEID=2782470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_206C;SPAN=4537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:302 DP:539 GQ:99 PL:[850.9, 0.0, 458.1] SR:163 DR:175 LR:-857.2 LO:857.2);ALT=G[chr6:33048455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34205094	+	chr6	34208513	+	.	119	104	2787700_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2787700_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GCGC;SCTG=c_6_34202001_34227001_392C;SPAN=3419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:188 DP:119 GQ:50.8 PL:[557.8, 50.8, 0.0] SR:104 DR:119 LR:-557.8 LO:557.8);ALT=G[chr6:34208513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35265732	+	chr6	35277445	+	.	50	10	2791568_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=2791568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35255501_35280501_285C;SPAN=11713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:101 GQ:91.7 PL:[151.1, 0.0, 91.7] SR:10 DR:50 LR:-151.6 LO:151.6);ALT=G[chr6:35277445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35626434	+	chr6	35629745	+	.	83	77	2793238_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2793238_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35623001_35648001_95C;SPAN=3311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:38 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:77 DR:83 LR:-406.0 LO:406.0);ALT=G[chr6:35629745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35766788	+	chr6	35754561	+	.	96	58	2794250_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAC;MAPQ=60;MATEID=2794250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35745501_35770501_86C;SPAN=12227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:130 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:58 DR:96 LR:-386.2 LO:386.2);ALT=]chr6:35766788]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	36562258	+	chr6	36564537	+	.	131	25	2797146_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2797146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36554001_36579001_207C;SPAN=2279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:135 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:25 DR:131 LR:-448.9 LO:448.9);ALT=G[chr6:36564537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37451113	+	chr6	37467595	+	.	31	0	2800705_1	83.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2800705_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:37451113(+)-6:37467595(-)__6_37460501_37485501D;SPAN=16482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:68 GQ:80.6 PL:[83.9, 0.0, 80.6] SR:0 DR:31 LR:-83.91 LO:83.91);ALT=T[chr6:37467595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37452972	+	chr6	37467598	+	.	48	8	2800707_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2800707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_37460501_37485501_440C;SPAN=14626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:72 GQ:33.5 PL:[139.1, 0.0, 33.5] SR:8 DR:48 LR:-142.3 LO:142.3);ALT=T[chr6:37467598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41755564	+	chr6	41756968	+	.	52	112	2814998_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2814998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_41748001_41773001_83C;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:119 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:112 DR:52 LR:-422.5 LO:422.5);ALT=G[chr6:41756968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41755578	+	chr12	125541044	-	.	37	0	2814999_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2814999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:41755578(+)-12:125541044(+)__6_41748001_41773001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:28 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:0 DR:37 LR:-108.9 LO:108.9);ALT=G]chr12:125541044];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	43025973	+	chr6	43027024	+	.	39	12	2820592_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2820592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_43022001_43047001_309C;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:108 GQ:99 PL:[119.3, 0.0, 142.4] SR:12 DR:39 LR:-119.3 LO:119.4);ALT=T[chr6:43027024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44081993	+	chr6	44095079	+	.	37	0	2824769_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2824769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44081993(+)-6:44095079(-)__6_44075501_44100501D;SPAN=13086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:136 GQ:85.4 PL:[85.4, 0.0, 243.8] SR:0 DR:37 LR:-85.29 LO:89.57);ALT=C[chr6:44095079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44214926	+	chr6	44217111	+	.	34	0	2825377_1	76.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2825377_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44214926(+)-6:44217111(-)__6_44198001_44223001D;SPAN=2185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:134 GQ:76.1 PL:[76.1, 0.0, 247.7] SR:0 DR:34 LR:-75.93 LO:81.1);ALT=T[chr6:44217111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44214931	+	chr6	44216351	+	.	72	0	2825378_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2825378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44214931(+)-6:44216351(-)__6_44198001_44223001D;SPAN=1420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:115 GQ:71.3 PL:[206.6, 0.0, 71.3] SR:0 DR:72 LR:-210.0 LO:210.0);ALT=A[chr6:44216351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	102283809	+	chr8	107556938	+	.	34	0	4012507_1	98.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4012507_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:102283809(+)-8:107556938(-)__8_107555001_107580001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:52 GQ:25.7 PL:[98.3, 0.0, 25.7] SR:0 DR:34 LR:-100.3 LO:100.3);ALT=T[chr8:107556938[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	107307807	+	chr8	105231728	+	CCATGATCAGTGGCCATG	32	57	2973824_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;INSERTION=CCATGATCAGTGGCCATG;MAPQ=60;MATEID=2973824_2;MATENM=1;NM=1;NUMPARTS=3;SCTG=c_6_107285501_107310501_193C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:42 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:57 DR:32 LR:-201.3 LO:201.3);ALT=C[chr8:105231728[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	105231899	+	chr6	107307808	+	CCATGATCAGTGGCCATG	32	38	4006369_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AC;INSERTION=CCATGATCAGTGGCCATG;MAPQ=60;MATEID=4006369_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_8_105227501_105252501_237C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:53 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:38 DR:32 LR:-178.2 LO:178.2);ALT=]chr8:105231899]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	108544251	+	chr6	108581964	+	.	72	99	2977550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2977550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_108559501_108584501_115C;SPAN=37713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:62 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:99 DR:72 LR:-406.0 LO:406.0);ALT=T[chr6:108581964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	111280048	+	chrX	106374932	+	.	52	0	7492079_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7492079_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:111280048(+)-23:106374932(-)__23_106354501_106379501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:26 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=A[chrX:106374932[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	139350013	+	chr6	139355290	+	.	31	40	3047348_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3047348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_139331501_139356501_335C;SPAN=5277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:96 GQ:76.4 PL:[155.6, 0.0, 76.4] SR:40 DR:31 LR:-157.0 LO:157.0);ALT=G[chr6:139355290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	149433833	+	chr20	16710782	-	.	33	0	6938925_1	92.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=6938925_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:149433833(+)-20:16710782(+)__20_16709001_16734001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:62 GQ:56 PL:[92.3, 0.0, 56.0] SR:0 DR:33 LR:-92.54 LO:92.54);ALT=A]chr20:16710782];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	154620006	+	chr6	154621505	+	.	123	77	3082933_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GGAAGCTGAGGCAGGAG;MAPQ=60;MATEID=3082933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_154595001_154620001_361C;SPAN=1499;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:19 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:77 DR:123 LR:-452.2 LO:452.2);ALT=G[chr6:154621505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	157699920	+	chr6	157703237	+	.	47	18	3090020_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCTCCCAGGTTCAAGCGATTCTCCTGCCTCAGCCTCCTGAGTAGCTGGGA;MAPQ=60;MATEID=3090020_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_6_157682001_157707001_3C;SPAN=3317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:38 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:18 DR:47 LR:-171.6 LO:171.6);ALT=A[chr6:157703237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	158589482	+	chr6	158613006	+	.	45	0	3092858_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3092858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:158589482(+)-6:158613006(-)__6_158613001_158638001D;SPAN=23524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:36 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=G[chr6:158613006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159968217	+	chr6	159970838	+	.	57	26	3096791_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGTACCACATTTTTTA;MAPQ=60;MATEID=3096791_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_159960501_159985501_195C;SPAN=2621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:59 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:26 DR:57 LR:-217.9 LO:217.9);ALT=A[chr6:159970838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	151134	+	chr7	160558	+	TGGCG	70	49	3125958_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TGGCG;MAPQ=60;MATEID=3125958_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_147001_172001_320C;SPAN=9424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:77 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:49 DR:70 LR:-293.8 LO:293.8);ALT=A[chr7:160558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1185078	+	chr7	1187655	+	.	57	20	3129900_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CACTCTTAAGTTTT;MAPQ=60;MATEID=3129900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1176001_1201001_348C;SPAN=2577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:67 DP:1556 GQ:99 PL:[0.0, 199.9, 4179.0] SR:20 DR:57 LR:200.4 LO:104.6);ALT=T[chr7:1187655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2284362	+	chr7	2289490	+	.	67	97	3133587_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3133587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_2278501_2303501_64C;SPAN=5128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:156 GQ:28.9 PL:[435.7, 28.9, 0.0] SR:97 DR:67 LR:-440.4 LO:440.4);ALT=G[chr7:2289490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	4081265	+	chr7	4082297	+	.	60	47	3140500_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3140500_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_7_4067001_4092001_137C;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:65 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:47 DR:60 LR:-241.0 LO:241.0);ALT=C[chr7:4082297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	8463551	+	chr7	8465542	+	.	61	26	3159575_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=3159575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_8452501_8477501_231C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:67 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:26 DR:61 LR:-214.6 LO:214.6);ALT=A[chr7:8465542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	9634650	+	chr7	9635978	+	.	123	69	3163237_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGAAAAGAGACTACTG;MAPQ=60;MATEID=3163237_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_9628501_9653501_19C;SPAN=1328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:44 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:69 DR:123 LR:-448.9 LO:448.9);ALT=G[chr7:9635978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	10491065	-	chr11	122932781	+	.	91	0	5033453_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5033453_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:10491065(-)-11:122932781(-)__11_122916501_122941501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:91 DP:165 GQ:99 PL:[255.8, 0.0, 143.6] SR:0 DR:91 LR:-257.3 LO:257.3);ALT=[chr11:122932781[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	26233316	+	chr7	26236021	+	CCAGGTCCTCCTCCATACCCATTATAGCCATCCCCAAATCCACGTCCACTGCCATATCCAT	43	75	3217639_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCAGGTCCTCCTCCATACCCATTATAGCCATCCCCAAATCCACGTCCACTGCCATATCCAT;MAPQ=60;MATEID=3217639_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26215001_26240001_244C;SPAN=2705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:131 GQ:8.7 PL:[333.3, 8.7, 0.0] SR:75 DR:43 LR:-346.1 LO:346.1);ALT=T[chr7:26236021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26237488	+	chr7	26240192	+	.	82	19	3217816_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3217816_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26239501_26264501_355C;SPAN=2704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:101 DP:135 GQ:29.6 PL:[296.9, 0.0, 29.6] SR:19 DR:82 LR:-309.4 LO:309.4);ALT=T[chr7:26240192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26241446	+	chr7	26245987	+	AATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA	33	97	3217824_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=GGCTCTGCCTCTTCAACTTTTTTACTCTTTCCATTCTGTTTTTTTCCCATTTTTTGCAATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA;INSERTION=AATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA;MAPQ=60;MATEID=3217824_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26239501_26264501_0C;SECONDARY;SPAN=4541;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:101 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:97 DR:33 LR:-366.4 LO:366.4);ALT=A[chr7:26245987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27779888	+	chr7	27788136	+	.	48	11	3224296_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3224296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27783001_27808001_516C;SPAN=8248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:11 DR:48 LR:-163.7 LO:163.7);ALT=G[chr7:27788136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	31315559	+	chr7	31318954	+	.	90	41	3235743_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GGTGGCTCACGCCTGTAATCCCAGCACTTTGG;MAPQ=60;MATEID=3235743_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_7_31311001_31336001_78C;SPAN=3395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:93 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:41 DR:90 LR:-349.9 LO:349.9);ALT=G[chr7:31318954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32390165	+	chr7	32393113	+	.	78	40	3239179_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTGACTAATATAT;MAPQ=60;MATEID=3239179_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_32389001_32414001_54C;SPAN=2948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:38 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:40 DR:78 LR:-290.5 LO:290.5);ALT=T[chr7:32393113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32526950	+	chr7	32529930	+	.	36	0	3239537_1	80.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3239537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:32526950(+)-7:32529930(-)__7_32511501_32536501D;SPAN=2980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:142 GQ:80.6 PL:[80.6, 0.0, 262.1] SR:0 DR:36 LR:-80.37 LO:85.85);ALT=G[chr7:32529930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32527411	+	chr7	32529930	+	.	53	0	3239539_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3239539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:32527411(+)-7:32529930(-)__7_32511501_32536501D;SPAN=2519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:144 GQ:99 PL:[136.1, 0.0, 212.0] SR:0 DR:53 LR:-135.9 LO:136.9);ALT=A[chr7:32529930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38218024	+	chr7	38247045	+	.	70	13	3259293_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGGT;MAPQ=60;MATEID=3259293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38195501_38220501_359C;SPAN=29021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:64 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:13 DR:70 LR:-211.3 LO:211.3);ALT=T[chr7:38247045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38289174	+	chr7	38295938	+	.	41	6	3259379_1	99.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3259379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38269001_38294001_169C;SPAN=6764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:63 GQ:16.1 PL:[134.9, 0.0, 16.1] SR:6 DR:41 LR:-139.9 LO:139.9);ALT=C[chr7:38295938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42964437	+	chr7	42971715	+	.	55	0	3275343_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3275343_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:42964437(+)-7:42971715(-)__7_42948501_42973501D;SPAN=7278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:159 GQ:99 PL:[138.5, 0.0, 247.4] SR:0 DR:55 LR:-138.5 LO:140.2);ALT=T[chr7:42971715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42966297	+	chr7	42971716	+	.	133	0	3275350_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3275350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:42966297(+)-7:42971716(-)__7_42948501_42973501D;SPAN=5419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:152 GQ:31 PL:[429.1, 31.0, 0.0] SR:0 DR:133 LR:-431.5 LO:431.5);ALT=T[chr7:42971716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	43906631	+	chr7	43908906	+	.	78	0	3278797_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3278797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:43906631(+)-7:43908906(-)__7_43904001_43929001D;SPAN=2275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:119 GQ:63.5 PL:[225.2, 0.0, 63.5] SR:0 DR:78 LR:-230.3 LO:230.3);ALT=C[chr7:43908906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44084420	+	chr7	44091428	+	GCTCTCTTTACCTATGAAGGCAACAGCAATGACATCCGCGTGGCTGGCACAGGG	65	56	3280111_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GCTCTCTTTACCTATGAAGGCAACAGCAATGACATCCGCGTGGCTGGCACAGGG;MAPQ=60;MATEID=3280111_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_7_44075501_44100501_437C;SPAN=7008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:134 GQ:56.3 PL:[267.5, 0.0, 56.3] SR:56 DR:65 LR:-275.0 LO:275.0);ALT=G[chr7:44091428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44880622	+	chr7	44887566	+	.	52	0	3283069_1	99.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3283069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44880622(+)-7:44887566(-)__7_44859501_44884501D;SPAN=6944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:58 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:52 LR:-171.1 LO:171.1);ALT=G[chr7:44887566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93277465	+	chr7	44887593	+	.	73	0	6038799_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6038799_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44887593(-)-15:93277465(+)__15_93271501_93296501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:92 GQ:5 PL:[216.2, 0.0, 5.0] SR:0 DR:73 LR:-227.9 LO:227.9);ALT=]chr15:93277465]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	45016673	+	chr7	45018464	+	.	45	21	3283667_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=3283667_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_45006501_45031501_206C;SPAN=1791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:119 GQ:99 PL:[139.4, 0.0, 149.3] SR:21 DR:45 LR:-139.4 LO:139.4);ALT=G[chr7:45018464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	45024073	+	chr7	45026145	+	.	35	0	3283706_1	83.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3283706_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:45024073(+)-7:45026145(-)__7_45006501_45031501D;SPAN=2072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:119 GQ:83.3 PL:[83.3, 0.0, 205.4] SR:0 DR:35 LR:-83.3 LO:86.15);ALT=C[chr7:45026145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	61848994	+	chr7	61857679	+	CAAATAT	53	48	3333354_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;INSERTION=CAAATAT;MAPQ=47;MATEID=3333354_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_7_61838001_61863001_89C;SPAN=8685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:144 GQ:93.2 PL:[254.9, 0.0, 93.2] SR:48 DR:53 LR:-258.8 LO:258.8);ALT=C[chr7:61857679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	62002310	+	chr7	62004852	+	.	89	35	3333854_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTTCTTTTGATAGAACAGTTTTGAAACACTCTTT;MAPQ=60;MATEID=3333854_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_61985001_62010001_172C;SPAN=2542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:26 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:35 DR:89 LR:-326.8 LO:326.8);ALT=T[chr7:62004852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64315824	+	chr7	64318059	+	.	84	38	3344483_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAATTTTATTTTATC;MAPQ=60;MATEID=3344483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_64312501_64337501_113C;SPAN=2235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:30 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:38 DR:84 LR:-300.4 LO:300.4);ALT=C[chr7:64318059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	65589705	+	chr7	65591966	+	.	42	42	3351273_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=3351273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65586501_65611501_276C;SPAN=2261;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:74 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:42 DR:42 LR:-217.9 LO:217.9);ALT=C[chr7:65591966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66030576	+	chr7	66258667	-	ACCTGCT	39	29	3353859_1	99.0	.	DISC_MAPQ=32;EVDNC=TSI_L;INSERTION=ACCTGCT;MAPQ=60;MATEID=3353859_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_7_66027501_66052501_45C;SPAN=228091;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:77 GQ:5.6 PL:[180.5, 0.0, 5.6] SR:29 DR:39 LR:-190.3 LO:190.3);ALT=C]chr7:66258667];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	66697505	+	chr7	66699292	+	.	45	18	3356890_1	99.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTGGG;MAPQ=60;MATEID=3356890_2;MATENM=0;NM=2;NUMPARTS=2;REPSEQ=GGG;SCTG=c_7_66689001_66714001_393C;SECONDARY;SPAN=1787;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:80 GQ:21.2 PL:[173.0, 0.0, 21.2] SR:18 DR:45 LR:-180.0 LO:180.0);ALT=G[chr7:66699292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	70426185	-	chr7	70438880	+	.	41	43	3372272_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=3372272_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_70437501_70462501_158C;SPAN=12695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:48 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:43 DR:41 LR:-224.5 LO:224.5);ALT=[chr7:70438880[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	71211913	+	chr7	71212956	+	.	51	32	3375663_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAAA;MAPQ=60;MATEID=3375663_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_71197001_71222001_193C;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:67 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:32 DR:51 LR:-208.0 LO:208.0);ALT=A[chr7:71212956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73549766	+	chr7	73550967	+	.	34	45	3387402_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTGAGA;MAPQ=60;MATEID=3387402_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_73549001_73574001_217C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:26 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:45 DR:34 LR:-204.7 LO:204.7);ALT=A[chr7:73550967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73624418	+	chr7	73629150	+	.	74	7	3387642_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3387642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_73622501_73647501_218C;SPAN=4732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:109 GQ:39.8 PL:[224.6, 0.0, 39.8] SR:7 DR:74 LR:-232.0 LO:232.0);ALT=G[chr7:73629150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75363121	+	chr7	75368118	+	.	55	21	3398591_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=3398591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75362001_75387001_343C;SPAN=4997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:137 GQ:99 PL:[174.2, 0.0, 157.7] SR:21 DR:55 LR:-174.2 LO:174.2);ALT=G[chr7:75368118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75677544	+	chr7	75684146	+	.	110	54	3400448_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3400448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75656001_75681001_239C;SPAN=6602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:47 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:54 DR:110 LR:-412.6 LO:412.6);ALT=G[chr7:75684146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80268062	+	chr7	80275402	+	.	61	22	3417511_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3417511_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_80262001_80287001_273C;SPAN=7340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:134 GQ:86 PL:[237.8, 0.0, 86.0] SR:22 DR:61 LR:-241.5 LO:241.5);ALT=G[chr7:80275402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	81789164	+	chr10	60902930	-	.	84	47	3422222_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=3422222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_81781001_81806001_162C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:43 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:47 DR:84 LR:-326.8 LO:326.8);ALT=T]chr10:60902930];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	89810409	+	chr7	89812600	+	.	81	81	3446317_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=3446317_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_89792501_89817501_168C;SPAN=2191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:37 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:81 DR:81 LR:-399.4 LO:399.4);ALT=C[chr7:89812600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98972405	+	chr7	98983323	+	.	95	27	3478075_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3478075_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98980001_99005001_174C;SPAN=10918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:72 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:27 DR:95 LR:-280.6 LO:280.6);ALT=G[chr7:98983323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99006156	-	chr12	119632708	+	.	41	0	5361551_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5361551_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99006156(-)-12:119632708(-)__12_119609001_119634001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:41 LR:-132.0 LO:132.0);ALT=[chr12:119632708[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	99006678	+	chr7	99008684	+	.	37	0	3478319_1	95.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3478319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99006678(+)-7:99008684(-)__7_99004501_99029501D;SPAN=2006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:98 GQ:95.6 PL:[95.6, 0.0, 141.8] SR:0 DR:37 LR:-95.59 LO:96.09);ALT=A[chr7:99008684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99041062	+	chr12	56211447	+	.	51	0	5202108_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5202108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99041062(+)-12:56211447(-)__12_56203001_56228001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:68 GQ:14.6 PL:[149.9, 0.0, 14.6] SR:0 DR:51 LR:-156.4 LO:156.4);ALT=A[chr12:56211447[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	99056908	+	chr7	99063733	+	.	31	0	3478463_1	67.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=3478463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99056908(+)-7:99063733(-)__7_99053501_99078501D;SPAN=6825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:128 GQ:67.7 PL:[67.7, 0.0, 242.6] SR:0 DR:31 LR:-67.65 LO:73.21);ALT=A[chr7:99063733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99697418	+	chr7	99698897	+	.	33	0	3480936_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3480936_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99697418(+)-7:99698897(-)__7_99690501_99715501D;SPAN=1479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:87 GQ:85.4 PL:[85.4, 0.0, 125.0] SR:0 DR:33 LR:-85.36 LO:85.79);ALT=A[chr7:99698897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99746760	+	chr7	99751020	+	.	122	0	3481465_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3481465_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99746760(+)-7:99751020(-)__7_99739501_99764501D;SPAN=4260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:149 GQ:0.6 PL:[363.0, 0.6, 0.0] SR:0 DR:122 LR:-385.1 LO:385.1);ALT=G[chr7:99751020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99747240	+	chr7	99751488	+	.	31	0	3481468_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3481468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99747240(+)-7:99751488(-)__7_99739501_99764501D;SPAN=4248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:164 GQ:58.1 PL:[58.1, 0.0, 338.6] SR:0 DR:31 LR:-57.9 LO:69.4);ALT=A[chr7:99751488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99930229	+	chr7	99933460	+	.	35	0	3482947_1	86.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=3482947_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99930229(+)-7:99933460(-)__7_99911001_99936001D;SPAN=3231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:106 GQ:86.9 PL:[86.9, 0.0, 169.4] SR:0 DR:35 LR:-86.82 LO:88.31);ALT=A[chr7:99933460[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100271547	+	chr7	100273797	+	.	91	13	3484111_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3484111_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_100254001_100279001_52C;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:97 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:13 DR:91 LR:-287.2 LO:287.2);ALT=G[chr7:100273797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100533453	+	chr7	100536238	+	.	60	45	3485291_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAGGTTGCAGTGAG;MAPQ=60;MATEID=3485291_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_100523501_100548501_71C;SPAN=2785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:87 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:45 DR:60 LR:-256.6 LO:256.6);ALT=G[chr7:100536238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100861545	+	chr7	100865880	+	.	51	0	3486487_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3486487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100861545(+)-7:100865880(-)__7_100842001_100867001D;SPAN=4335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:109 GQ:99 PL:[138.8, 0.0, 125.6] SR:0 DR:51 LR:-138.9 LO:138.9);ALT=C[chr7:100865880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100861549	+	chr7	100866756	+	.	33	0	3487180_1	91.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3487180_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100861549(+)-7:100866756(-)__7_100866501_100891501D;SPAN=5207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=G[chr7:100866756[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100884188	+	chr7	100888241	+	CTCGAGCAGCACGATGCCTTTACGGATGTCATCATTGTACTTGCTCCGCACCAGGCACCAGGCGTACTCAAACTGCGTGCTCTTGGACACCGAGCCTGCTGCCTTCTCAGACTGAAATTTCTTTTCAAACTT	37	101	3487264_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTCGAGCAGCACGATGCCTTTACGGATGTCATCATTGTACTTGCTCCGCACCAGGCACCAGGCGTACTCAAACTGCGTGCTCTTGGACACCGAGCCTGCTGCCTTCTCAGACTGAAATTTCTTTTCAAACTT;MAPQ=60;MATEID=3487264_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_100866501_100891501_246C;SPAN=4053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:138 GQ:2.3 PL:[332.3, 0.0, 2.3] SR:101 DR:37 LR:-352.4 LO:352.4);ALT=C[chr7:100888241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101001266	+	chr7	101003796	+	.	50	28	3489005_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCAATTTTTGTATTTTT;MAPQ=38;MATEID=3489005_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_7_100989001_101014001_394C;SPAN=2530;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:56 GQ:21 PL:[231.0, 21.0, 0.0] SR:28 DR:50 LR:-231.1 LO:231.1);ALT=T[chr7:101003796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101059188	+	chr7	101060267	+	.	45	36	3488111_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CCCGCCTCAGCCTCCCAAAGTGCTGGGATTA;MAPQ=60;MATEID=3488111_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_7_101038001_101063001_241C;SPAN=1079;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:72 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:36 DR:45 LR:-211.3 LO:211.3);ALT=A[chr7:101060267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101459373	+	chr7	101559392	+	.	36	9	3490506_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=3490506_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_101552501_101577501_190C;SPAN=100019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:9 DR:36 LR:-118.8 LO:118.8);ALT=G[chr7:101559392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104612302	+	chr7	104485067	+	.	57	37	3503166_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3503166_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104590501_104615501_205C;SPAN=127235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:82 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:37 DR:57 LR:-244.3 LO:244.3);ALT=]chr7:104612302]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	105739729	+	chr7	105752586	+	.	76	44	3507980_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3507980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105717501_105742501_365C;SPAN=12857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:68 GQ:24 PL:[264.0, 24.0, 0.0] SR:44 DR:76 LR:-264.1 LO:264.1);ALT=C[chr7:105752586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	125264220	+	chr12	74014367	+	ATTATA	49	58	3568962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTATA;MAPQ=60;MATEID=3568962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_125244001_125269001_225C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:61 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:58 DR:49 LR:-254.2 LO:254.2);ALT=C[chr12:74014367[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	125746123	+	chr7	126166901	+	T	47	38	3570834_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=3570834_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_126150501_126175501_101C;SPAN=420778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:63 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:38 DR:47 LR:-211.3 LO:211.3);ALT=A[chr7:126166901[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	126045889	+	chr7	126051448	+	.	50	53	3570696_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=3570696_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_126028001_126053001_151C;SPAN=5559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:25 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:53 DR:50 LR:-257.5 LO:257.5);ALT=C[chr7:126051448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	126098488	-	chr7	126167441	+	.	39	48	3570835_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAT;MAPQ=60;MATEID=3570835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_126150501_126175501_371C;SPAN=68953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:72 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:48 DR:39 LR:-234.4 LO:234.4);ALT=[chr7:126167441[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	128096078	+	chr7	128097253	+	.	35	12	3580607_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3580607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_128086001_128111001_215C;SPAN=1175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:173 GQ:75.5 PL:[75.5, 0.0, 342.8] SR:12 DR:35 LR:-75.27 LO:85.08);ALT=G[chr7:128097253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128503047	+	chr12	48478956	+	.	40	0	3583351_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3583351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128503047(+)-12:48478956(-)__7_128502501_128527501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:128 GQ:97.4 PL:[97.4, 0.0, 212.9] SR:0 DR:40 LR:-97.36 LO:99.74);ALT=A[chr12:48478956[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	128503128	+	chr7	128505428	+	.	56	0	3583352_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3583352_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128503128(+)-7:128505428(-)__7_128502501_128527501D;SPAN=2300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:173 GQ:99 PL:[138.2, 0.0, 280.1] SR:0 DR:56 LR:-138.0 LO:140.7);ALT=C[chr7:128505428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128578155	+	chr7	128582120	+	.	38	0	3584032_1	86.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3584032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128578155(+)-7:128582120(-)__7_128576001_128601001D;SPAN=3965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:146 GQ:86 PL:[86.0, 0.0, 267.5] SR:0 DR:38 LR:-85.88 LO:91.13);ALT=C[chr7:128582120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	129050411	+	chr9	116037593	+	.	33	0	3586964_1	91.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=3586964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:129050411(+)-9:116037593(-)__7_129041501_129066501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=T[chr9:116037593[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	133785003	+	chr7	133798330	+	.	129	68	3612727_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=60;MATEID=3612727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_133794501_133819501_217C;SPAN=13327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:161 DP:77 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:68 DR:129 LR:-475.3 LO:475.3);ALT=C[chr7:133798330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135347372	+	chr7	135358838	+	.	62	0	3621458_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3621458_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:135347372(+)-7:135358838(-)__7_135338001_135363001D;SPAN=11466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:189 GQ:99 PL:[153.5, 0.0, 305.3] SR:0 DR:62 LR:-153.5 LO:156.2);ALT=G[chr7:135358838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	137613141	+	chr7	137620615	+	.	32	0	3632445_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3632445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:137613141(+)-7:137620615(-)__7_137616501_137641501D;SPAN=7474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:61 GQ:56.3 PL:[89.3, 0.0, 56.3] SR:0 DR:32 LR:-89.43 LO:89.43);ALT=G[chr7:137620615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139026270	+	chr7	139030246	+	.	46	32	3641275_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=3641275_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139013001_139038001_355C;SPAN=3976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:177 GQ:99 PL:[160.1, 0.0, 269.0] SR:32 DR:46 LR:-160.0 LO:161.5);ALT=T[chr7:139030246[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139218974	-	chr14	69864948	+	.	85	8	3642952_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CATCGCGCCAAACTCT;MAPQ=32;MATEID=3642952_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_7_139209001_139234001_457C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:83 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:8 DR:85 LR:-267.4 LO:267.4);ALT=[chr14:69864948[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	140397086	+	chr7	140402665	+	.	69	0	3650450_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3650450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:140397086(+)-7:140402665(-)__7_140385001_140410001D;SPAN=5579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:209 GQ:99 PL:[171.2, 0.0, 336.2] SR:0 DR:69 LR:-171.1 LO:174.1);ALT=T[chr7:140402665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140710474	+	chr7	140714709	+	.	33	0	3651988_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3651988_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:140710474(+)-7:140714709(-)__7_140703501_140728501D;SPAN=4235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:188 GQ:58 PL:[58.0, 0.0, 398.0] SR:0 DR:33 LR:-58.0 LO:72.7);ALT=G[chr7:140714709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142824847	+	chr7	142893908	+	.	109	47	3661916_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTAAA;MAPQ=60;MATEID=3661916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_142884001_142909001_275C;SPAN=69061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:54 GQ:36 PL:[396.0, 36.0, 0.0] SR:47 DR:109 LR:-396.1 LO:396.1);ALT=A[chr7:142893908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150746657	+	chr15	84810725	+	.	44	33	3692179_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3692179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_150724001_150749001_17C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:31 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:33 DR:44 LR:-191.4 LO:191.4);ALT=C[chr15:84810725[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	152281703	+	chr7	152284306	+	.	43	38	3695637_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=CACATGTTTTA;MAPQ=60;MATEID=3695637_2;MATENM=2;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_7_152267501_152292501_263C;SPAN=2603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:37 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:38 DR:43 LR:-194.7 LO:194.7);ALT=A[chr7:152284306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11245561	+	chr8	11247208	+	.	48	45	3743746_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAG;MAPQ=60;MATEID=3743746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11245501_11270501_317C;SPAN=1647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:66 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:45 DR:48 LR:-208.0 LO:208.0);ALT=G[chr8:11247208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11660441	+	chr8	11666300	+	.	50	23	3745060_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3745060_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_11662001_11687001_301C;SPAN=5859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:60 GQ:9.6 PL:[165.0, 9.6, 0.0] SR:23 DR:50 LR:-167.9 LO:167.9);ALT=G[chr8:11666300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11710989	+	chr8	11725507	+	.	40	6	3745233_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=3745233_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11686501_11711501_378C;SPAN=14518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:51 GQ:2.9 PL:[118.4, 0.0, 2.9] SR:6 DR:40 LR:-124.4 LO:124.4);ALT=C[chr8:11725507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	12427810	+	chr8	12432836	+	GGAATTTTGTG	36	29	3752489_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;INSERTION=GGAATTTTGTG;MAPQ=60;MATEID=3752489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_12421501_12446501_1306C;SPAN=5026;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:256 GQ:99 PL:[118.9, 0.0, 501.8] SR:29 DR:36 LR:-118.8 LO:132.2);ALT=G[chr8:12432836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	15289364	+	chr13	74314062	-	.	57	70	3757473_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TATGTT;MAPQ=60;MATEID=3757473_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_15288001_15313001_184C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:31 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:70 DR:57 LR:-326.8 LO:326.8);ALT=T]chr13:74314062];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	15289367	-	chr13	74313858	+	.	72	80	3757475_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGGC;MAPQ=60;MATEID=3757475_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_15288001_15313001_68C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:31 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:80 DR:72 LR:-369.7 LO:369.7);ALT=[chr13:74313858[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	29927576	+	chr8	29940363	+	.	33	29	3801846_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3801846_2;MATENM=0;NM=2;NUMPARTS=3;REPSEQ=GGG;SCTG=c_8_29939001_29964001_338C;SPAN=12787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:139 GQ:99 PL:[120.8, 0.0, 216.5] SR:29 DR:33 LR:-120.8 LO:122.3);ALT=C[chr8:29940363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29931572	+	chr8	29940363	+	.	84	90	3801848_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3801848_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_29939001_29964001_156C;SPAN=8791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:139 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:90 DR:84 LR:-412.6 LO:412.6);ALT=C[chr8:29940363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29953095	+	chr8	29961815	+	.	72	0	3801898_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3801898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:29953095(+)-8:29961815(-)__8_29939001_29964001D;SPAN=8720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:95 GQ:17.3 PL:[212.0, 0.0, 17.3] SR:0 DR:72 LR:-221.5 LO:221.5);ALT=G[chr8:29961815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7167959	+	chr8	30145402	+	.	35	43	6301911_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=T;MAPQ=60;MATEID=6301911_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_17_7154001_7179001_15C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:50 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:43 DR:35 LR:-201.3 LO:201.3);ALT=]chr17:7167959]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	37888239	+	chr8	37914597	+	.	69	72	3824402_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGGTA;MAPQ=60;MATEID=3824402_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_37901501_37926501_31C;SPAN=26358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:53 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:72 DR:69 LR:-356.5 LO:356.5);ALT=A[chr8:37914597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	39232074	+	chr8	39387229	+	T	46	32	3829053_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=3829053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_39371501_39396501_56C;SPAN=155155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:21 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:32 DR:46 LR:-188.1 LO:188.1);ALT=G[chr8:39387229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	40289707	+	chr8	40296198	+	.	76	59	3832045_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAAAATACACAGGA;MAPQ=60;MATEID=3832045_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_8_40278001_40303001_55C;SPAN=6491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:33 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:59 DR:76 LR:-303.7 LO:303.7);ALT=A[chr8:40296198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42190485	+	chr8	42194353	+	.	95	0	3837614_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCTACTCGGGAGGCTGAGGCAGGAGAATCGCTTGAACCCGGGAGGCAGAGGTTGCAGTGAGCCGAGATCGTGCCATTGCACTCC;MAPQ=60;MATEID=3837614_2;MATENM=2;NM=4;NUMPARTS=2;SCTG=c_8_42189001_42214001_113C;SPAN=3868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:5 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:0 DR:95 LR:-280.6 LO:280.6);ALT=C[chr8:42194353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	71583571	+	chr8	71584644	+	.	84	72	3909790_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATGATCTCATTTTTTT;MAPQ=60;MATEID=3909790_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_71564501_71589501_137C;SPAN=1073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:52 GQ:33 PL:[363.0, 33.0, 0.0] SR:72 DR:84 LR:-363.1 LO:363.1);ALT=T[chr8:71584644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	72214752	+	chr8	72217809	+	.	45	33	3911452_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGCTGA;MAPQ=60;MATEID=3911452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_72201501_72226501_151C;SPAN=3057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:33 DR:45 LR:-205.9 LO:205.9);ALT=A[chr8:72217809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	73787775	+	chr8	73793824	+	.	62	57	3915763_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGCAAATCTT;MAPQ=60;MATEID=3915763_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_73769501_73794501_251C;SPAN=6049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:127 GQ:5.3 PL:[302.3, 0.0, 5.3] SR:57 DR:62 LR:-319.7 LO:319.7);ALT=T[chr8:73793824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	75362871	+	chr8	75367000	+	CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA	34	56	3920406_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA;MAPQ=60;MATEID=3920406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_75337501_75362501_106C;SPAN=4129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:0 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:56 DR:34 LR:-208.0 LO:208.0);ALT=A[chr8:75367000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	82045018	+	chr8	82046625	+	TTACGT	70	36	3937783_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;INSERTION=TTACGT;MAPQ=60;MATEID=3937783_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_8_82026001_82051001_324C;SPAN=1607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:59 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:36 DR:70 LR:-267.4 LO:267.4);ALT=G[chr8:82046625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	82192863	+	chr11	59549161	-	.	58	0	4874864_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=4874864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:82192863(+)-11:59549161(+)__11_59535001_59560001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:43 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=G]chr11:59549161];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	83269755	+	chr8	83295603	+	.	41	27	3941214_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTATCT;MAPQ=60;MATEID=3941214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_83251001_83276001_12C;SPAN=25848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:29 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:27 DR:41 LR:-151.8 LO:151.8);ALT=T[chr8:83295603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	99055064	+	chr8	99057733	+	.	34	0	3987718_1	0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=3987718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:99055064(+)-8:99057733(-)__8_99053501_99078501D;SPAN=2669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:34 DP:814 GQ:99 PL:[0.0, 107.9, 2192.0] SR:0 DR:34 LR:108.3 LO:52.63);ALT=G[chr8:99057733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	100899897	+	chr8	100905864	+	.	45	0	3992816_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3992816_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:100899897(+)-8:100905864(-)__8_100891001_100916001D;SPAN=5967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:148 GQ:99 PL:[108.5, 0.0, 250.4] SR:0 DR:45 LR:-108.4 LO:111.6);ALT=G[chr8:100905864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	100904324	+	chr8	100905793	+	.	61	0	3992830_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3992830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:100904324(+)-8:100905793(-)__8_100891001_100916001D;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:79 GQ:11.6 PL:[179.9, 0.0, 11.6] SR:0 DR:61 LR:-188.7 LO:188.7);ALT=A[chr8:100905793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101162981	+	chr8	101164049	+	.	46	0	3993692_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3993692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101162981(+)-8:101164049(-)__8_101160501_101185501D;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:104 GQ:99 PL:[123.8, 0.0, 127.1] SR:0 DR:46 LR:-123.7 LO:123.7);ALT=C[chr8:101164049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101162989	+	chr8	101165521	+	.	47	0	3993693_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3993693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101162989(+)-8:101165521(-)__8_101160501_101185501D;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:100 GQ:99 PL:[128.0, 0.0, 114.8] SR:0 DR:47 LR:-128.1 LO:128.1);ALT=G[chr8:101165521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101961128	+	chr8	101964156	+	.	106	0	3996479_1	99.0	.	DISC_MAPQ=5;EVDNC=DSCRD;IMPRECISE;MAPQ=5;MATEID=3996479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101961128(+)-8:101964156(-)__8_101944501_101969501D;SPAN=3028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:96 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=T[chr8:101964156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101964157	-	chr10	23425817	+	.	31	15	4543359_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCGCCACCACCCACTCCGGACACAG;MAPQ=60;MATEID=4543359_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_23422001_23447001_75C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:54 GQ:18.5 PL:[110.9, 0.0, 18.5] SR:15 DR:31 LR:-114.4 LO:114.4);ALT=[chr10:23425817[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	109252371	+	chr8	109260871	+	.	110	0	4017307_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=4017307_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:109252371(+)-8:109260871(-)__8_109245501_109270501D;SPAN=8500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:90 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:110 LR:-326.8 LO:326.8);ALT=A[chr8:109260871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109254166	+	chr8	109260881	+	.	143	0	4017313_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=4017313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:109254166(+)-8:109260881(-)__8_109245501_109270501D;SPAN=6715;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:163 GQ:34 PL:[462.1, 34.0, 0.0] SR:0 DR:143 LR:-464.5 LO:464.5);ALT=A[chr8:109260881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110346705	+	chr8	110348356	+	.	31	33	4020045_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4020045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110323501_110348501_3C;SPAN=1651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:128 GQ:99 PL:[130.4, 0.0, 179.9] SR:33 DR:31 LR:-130.4 LO:130.8);ALT=T[chr8:110348356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110346718	+	chr8	110351547	+	.	31	0	4020047_1	84.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4020047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:110346718(+)-8:110351547(-)__8_110323501_110348501D;SPAN=4829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:66 GQ:74.6 PL:[84.5, 0.0, 74.6] SR:0 DR:31 LR:-84.47 LO:84.47);ALT=T[chr8:110351547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	112294052	+	chr8	112297140	+	.	108	86	4024740_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4024740_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_112283501_112308501_73C;SPAN=3088;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:41 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:86 DR:108 LR:-458.8 LO:458.8);ALT=G[chr8:112297140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	125551262	-	chr10	64981924	+	.	45	0	4060953_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4060953_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:125551262(-)-10:64981924(-)__8_125538001_125563001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:0 DR:45 LR:-141.9 LO:141.9);ALT=[chr10:64981924[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	125551528	+	chr8	125555326	+	.	121	37	4060956_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4060956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_125538001_125563001_3C;SPAN=3798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:119 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:37 DR:121 LR:-422.5 LO:422.5);ALT=G[chr8:125555326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	126595129	+	chr8	126601135	+	.	104	46	4064665_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACTCACA;MAPQ=60;MATEID=4064665_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_126591501_126616501_153C;SPAN=6006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:156 GQ:19 PL:[415.9, 19.0, 0.0] SR:46 DR:104 LR:-426.4 LO:426.4);ALT=A[chr8:126601135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	127192205	+	chr8	127194572	+	T	47	42	4065851_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=4065851_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_127179501_127204501_144C;SPAN=2367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:60 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:42 DR:47 LR:-224.5 LO:224.5);ALT=C[chr8:127194572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	134972222	-	chr18	57070970	+	.	45	0	6641939_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6641939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:134972222(-)-18:57070970(-)__18_57060501_57085501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:33 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=[chr18:57070970[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	144100003	+	chr8	144102299	+	.	57	18	4114262_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4114262_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_144084501_144109501_279C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:70 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:18 DR:57 LR:-208.0 LO:208.0);ALT=G[chr8:144102299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145651208	+	chr8	145653869	+	.	52	0	4119069_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4119069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145651208(+)-8:145653869(-)__8_145628001_145653001D;SPAN=2661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:29 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=C[chr8:145653869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34618018	+	chr9	34620362	+	.	42	0	4179209_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4179209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:34618018(+)-9:34620362(-)__9_34594001_34619001D;SPAN=2344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:47 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:42 LR:-137.9 LO:137.9);ALT=C[chr9:34620362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34618759	+	chr9	34620363	+	.	51	25	4179028_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=4179028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_34618501_34643501_268C;SPAN=1604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:115 GQ:99 PL:[163.7, 0.0, 114.2] SR:25 DR:51 LR:-164.0 LO:164.0);ALT=T[chr9:34620363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35725727	+	chr9	35732069	+	.	51	5	4183288_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCTG;MAPQ=60;MATEID=4183288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35721001_35746001_51C;SPAN=6342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:97 GQ:79.4 PL:[155.3, 0.0, 79.4] SR:5 DR:51 LR:-156.6 LO:156.6);ALT=G[chr9:35732069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35813784	+	chr9	35814894	+	.	58	20	4183550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=4183550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35794501_35819501_373C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:133 GQ:99 PL:[191.9, 0.0, 129.2] SR:20 DR:58 LR:-192.3 LO:192.3);ALT=G[chr9:35814894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136870	+	chr9	36147778	+	.	31	0	4184927_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4184927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136870(+)-9:36147778(-)__9_36113001_36138001D;SPAN=10908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:36 GQ:6.3 PL:[99.0, 6.3, 0.0] SR:0 DR:31 LR:-99.82 LO:99.82);ALT=G[chr9:36147778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136870	+	chr9	36148542	+	.	47	0	4184928_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4184928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136870(+)-9:36148542(-)__9_36113001_36138001D;SPAN=11672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:36 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=G[chr9:36148542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36362896	+	chr9	36364080	+	.	134	101	4185954_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GCCTCCCAAAGTGCT;MAPQ=0;MATEID=4185954_2;MATENM=1;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_9_36358001_36383001_217C;SECONDARY;SPAN=1184;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:222 DP:39 GQ:59.8 PL:[656.8, 59.8, 0.0] SR:101 DR:134 LR:-656.9 LO:656.9);ALT=T[chr9:36364080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37422830	+	chr9	37424842	+	.	86	43	4189930_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4189930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37411501_37436501_296C;SPAN=2012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:109 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:43 DR:86 LR:-326.8 LO:326.8);ALT=A[chr9:37424842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37588930	+	chr9	37592307	+	.	58	4	4190789_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4190789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37583001_37608001_124C;SPAN=3377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:106 GQ:83.6 PL:[172.7, 0.0, 83.6] SR:4 DR:58 LR:-174.3 LO:174.3);ALT=C[chr9:37592307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37637304	+	chr11	66036196	-	.	49	0	4894603_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4894603_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:37637304(+)-11:66036196(+)__11_66027501_66052501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:44 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:49 LR:-145.2 LO:145.2);ALT=G]chr11:66036196];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	38243898	+	chr15	63770026	+	.	31	0	5969671_1	89.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5969671_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:38243898(+)-15:63770026(-)__15_63749001_63774001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:20 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=A[chr15:63770026[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	93564288	+	chr9	93606135	+	.	48	0	4329568_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4329568_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:93564288(+)-9:93606135(-)__9_93590001_93615001D;SPAN=41847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:55 GQ:11.4 PL:[155.1, 11.4, 0.0] SR:0 DR:48 LR:-155.5 LO:155.5);ALT=G[chr9:93606135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	94395817	+	chr9	94403299	+	.	51	46	4332069_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=4332069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_94374001_94399001_58C;SPAN=7482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:45 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:46 DR:51 LR:-227.8 LO:227.8);ALT=A[chr9:94403299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95858634	+	chr9	95869954	+	.	63	21	4337099_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4337099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_95868501_95893501_16C;SPAN=11320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:58 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:21 DR:63 LR:-201.3 LO:201.3);ALT=G[chr9:95869954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95888921	+	chr9	95896425	+	.	44	9	4337300_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4337300_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_95893001_95918001_203C;SPAN=7504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:35 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:9 DR:44 LR:-145.2 LO:145.2);ALT=C[chr9:95896425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	101984648	+	chr9	101990179	+	CTGCCGGACAGTGGATCCCGCCGCCCGGGCGGCCACTGCTTTGCTGGGAGAGCGCCCTGAGGATCCCACGTTAGTGCCACTGGGGGTCGGACCAGG	62	146	4358926_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTGCCGGACAGTGGATCCCGCCGCCCGGGCGGCCACTGCTTTGCTGGGAGAGCGCCCTGAGGATCCCACGTTAGTGCCACTGGGGGTCGGACCAGG;MAPQ=60;MATEID=4358926_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_101969001_101994001_136C;SPAN=5531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:185 DP:150 GQ:49.9 PL:[547.9, 49.9, 0.0] SR:146 DR:62 LR:-547.9 LO:547.9);ALT=G[chr9:101990179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	105967270	+	chr17	74553940	-	.	99	0	6501910_1	99.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=6501910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:105967270(+)-17:74553940(+)__17_74529001_74554001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:39 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:0 DR:99 LR:-293.8 LO:293.8);ALT=C]chr17:74553940];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	106568322	+	chr9	106569729	+	.	45	0	4371896_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4371896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:106568322(+)-9:106569729(-)__9_106550501_106575501D;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=A[chr9:106569729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	107510133	+	chr9	107513233	+	.	46	18	4374800_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=4374800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_107506001_107531001_333C;SPAN=3100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:112 GQ:99 PL:[151.4, 0.0, 118.4] SR:18 DR:46 LR:-151.4 LO:151.4);ALT=G[chr9:107513233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110033454	+	chr9	110035446	+	.	62	22	4382962_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATTATTATTATT;MAPQ=60;MATEID=4382962_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_110029501_110054501_364C;SPAN=1992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:66 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:22 DR:62 LR:-227.8 LO:227.8);ALT=T[chr9:110035446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110537535	+	chr9	110540596	+	.	78	34	4384765_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TAAAAATATTTTGTA;MAPQ=60;MATEID=4384765_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_110519501_110544501_1C;SPAN=3061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:53 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:34 DR:78 LR:-283.9 LO:283.9);ALT=A[chr9:110540596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	117350201	+	chr9	117354832	+	.	87	52	4408633_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4408633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_117330501_117355501_306C;SPAN=4631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:119 DP:185 GQ:99 PL:[342.8, 0.0, 105.2] SR:52 DR:87 LR:-349.6 LO:349.6);ALT=G[chr9:117354832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124030552	+	chr9	124064234	+	.	84	0	4429176_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4429176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:124030552(+)-9:124064234(-)__9_124043501_124068501D;SPAN=33682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:67 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=G[chr9:124064234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124043840	+	chr9	124064239	+	.	33	47	4429179_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4429179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_124043501_124068501_195C;SPAN=20399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:132 GQ:99 PL:[202.1, 0.0, 116.3] SR:47 DR:33 LR:-203.1 LO:203.1);ALT=G[chr9:124064239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127176335	+	chr9	127177645	+	.	55	0	4439715_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4439715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127176335(+)-9:127177645(-)__9_127155001_127180001D;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:112 GQ:99 PL:[151.4, 0.0, 118.4] SR:0 DR:55 LR:-151.4 LO:151.4);ALT=A[chr9:127177645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127933461	+	chr9	127951923	+	.	33	22	4442688_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4442688_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127939001_127964001_116C;SPAN=18462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:59 GQ:23.6 PL:[119.3, 0.0, 23.6] SR:22 DR:33 LR:-123.0 LO:123.0);ALT=T[chr9:127951923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130922765	+	chr9	130925719	+	.	137	104	4453309_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4453309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_130903501_130928501_315C;SPAN=2954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:198 DP:184 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:104 DR:137 LR:-587.5 LO:587.5);ALT=G[chr9:130925719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131085215	+	chr9	131087419	+	.	32	0	4453969_1	71.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4453969_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131085215(+)-9:131087419(-)__9_131075001_131100001D;SPAN=2204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:128 GQ:71 PL:[71.0, 0.0, 239.3] SR:0 DR:32 LR:-70.95 LO:76.08);ALT=G[chr9:131087419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131403219	+	chr9	131418829	+	GTCTCCCC	32	6	4455770_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTCTCCCC;MAPQ=60;MATEID=4455770_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_131418001_131443001_242C;SPAN=15610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:6 DR:32 LR:-110.1 LO:110.1);ALT=C[chr9:131418829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131412068	+	chr9	131413977	+	.	77	92	4455535_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AGGTCAGGAGTT;MAPQ=60;MATEID=4455535_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_131393501_131418501_219C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:26 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:92 DR:77 LR:-435.7 LO:435.7);ALT=T[chr9:131413977[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132026700	+	chr9	132028070	+	.	112	66	4458261_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCTGGGATTACAGGT;MAPQ=60;MATEID=4458261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132006001_132031001_79C;SPAN=1370;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:148 DP:42 GQ:40 PL:[439.0, 40.0, 0.0] SR:66 DR:112 LR:-439.0 LO:439.0);ALT=T[chr9:132028070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	133383116	+	chr9	133387421	+	GTGATCC	41	51	4463328_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=GTGATCC;MAPQ=60;MATEID=4463328_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_133378001_133403001_411C;SPAN=4305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:71 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:51 DR:41 LR:-254.2 LO:254.2);ALT=C[chr9:133387421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136221872	+	chr9	136223144	+	.	53	0	4473912_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4473912_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136221872(+)-9:136223144(-)__9_136220001_136245001D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:81 GQ:41 PL:[153.2, 0.0, 41.0] SR:0 DR:53 LR:-156.4 LO:156.4);ALT=G[chr9:136223144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	138479103	+	chr9	138480200	+	.	78	48	4481204_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGC;MAPQ=60;MATEID=4481204_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_138474001_138499001_134C;SPAN=1097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:26 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:48 DR:78 LR:-300.4 LO:300.4);ALT=C[chr9:138480200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139757955	+	chr9	139760649	+	.	136	0	4485715_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4485715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139757955(+)-9:139760649(-)__9_139748001_139773001D;SPAN=2694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:122 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:0 DR:136 LR:-402.7 LO:402.7);ALT=A[chr9:139760649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139758325	+	chr9	139760632	+	.	53	46	4485717_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=4485717_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_139748001_139773001_145C;SPAN=2307;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:122 GQ:99 PL:[155.3, 0.0, 138.8] SR:46 DR:53 LR:-155.1 LO:155.1);ALT=T[chr9:139760632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140500287	+	chr9	140507346	+	.	57	33	4488057_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4488057_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140507501_140532501_419C;SPAN=7059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:0 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:33 DR:57 LR:-201.3 LO:201.3);ALT=G[chr9:140507346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140783384	+	chr9	140785281	+	.	66	31	4489230_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4489230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140777001_140802001_444C;SPAN=1897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:173 GQ:99 PL:[240.5, 0.0, 177.8] SR:31 DR:66 LR:-240.8 LO:240.8);ALT=G[chr9:140785281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3109901	+	chr10	3124578	+	.	40	24	4495829_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4495829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3111501_3136501_3C;SPAN=14677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:44 GQ:12 PL:[132.0, 12.0, 0.0] SR:24 DR:40 LR:-132.0 LO:132.0);ALT=T[chr10:3124578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3357536	+	chr10	3356324	+	.	42	0	4496231_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4496231_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:3356324(-)-10:3357536(+)__10_3356501_3381501D;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:20 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=]chr10:3357536]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	3822424	+	chr10	3823832	+	.	33	6	4497208_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4497208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3797501_3822501_18C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:6 DR:33 LR:-115.5 LO:115.5);ALT=G[chr10:3823832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3824410	+	chr10	3827105	+	.	126	139	4496862_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTGT;MAPQ=60;MATEID=4496862_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3822001_3847001_130C;SPAN=2695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:192 DP:254 GQ:50.2 PL:[565.1, 0.0, 50.2] SR:139 DR:126 LR:-590.1 LO:590.1);ALT=T[chr10:3827105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	4290063	+	chr10	4291683	+	.	74	51	4497691_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4497691_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_10_4287501_4312501_0C;SPAN=1620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:26 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:51 DR:74 LR:-293.8 LO:293.8);ALT=C[chr10:4291683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	4376586	+	chr10	4374452	+	.	39	0	4497876_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4497876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:4374452(-)-10:4376586(+)__10_4361001_4386001D;SPAN=2134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:39 LR:-125.4 LO:125.4);ALT=]chr10:4376586]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	4708518	+	chr10	4710523	+	ATAG	50	42	4498208_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATAG;MAPQ=60;MATEID=4498208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_4704001_4729001_49C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:22 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:42 DR:50 LR:-208.0 LO:208.0);ALT=T[chr10:4710523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5889586	+	chr10	5892818	+	.	41	34	4500385_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTCTGCCTCCCAGGTTCAAGCAATTCT;MAPQ=45;MATEID=4500385_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5880001_5905001_252C;SPAN=3232;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:21 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:34 DR:41 LR:-188.1 LO:188.1);ALT=T[chr10:5892818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	6131119	+	chr10	6139007	+	.	39	0	4500777_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4500777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:6131119(+)-10:6139007(-)__10_6125001_6150001D;SPAN=7888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:50 GQ:6.2 PL:[115.1, 0.0, 6.2] SR:0 DR:39 LR:-121.1 LO:121.1);ALT=C[chr10:6139007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	6411580	+	chr10	6417630	+	.	40	24	4501537_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGCAAATCATTTTCCT;MAPQ=60;MATEID=4501537_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_6394501_6419501_193C;SPAN=6050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:139 GQ:99 PL:[147.2, 0.0, 190.1] SR:24 DR:40 LR:-147.2 LO:147.5);ALT=T[chr10:6417630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7077040	+	chr10	7078302	+	A	105	72	4502524_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4502524_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_7056001_7081001_305C;SPAN=1262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:37 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:72 DR:105 LR:-432.4 LO:432.4);ALT=T[chr10:7078302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7132876	+	chr19	17397640	+	.	31	28	6752156_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGAA;MAPQ=60;MATEID=6752156_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_17395001_17420001_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:31 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:28 DR:31 LR:-148.5 LO:148.5);ALT=A[chr19:17397640[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	7830227	+	chr10	7839010	+	ATTCAAGTTCGAAATATGGCAACTTTGAAAGATA	116	42	4503874_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GACTAAAGTCCATCAAAAACATCCAGAAAATTACCAAGTCTATGAAAATGGTAGCGGCAGCAAAATATGCCCGAGCTGAGAGAGAGCTGAAACCAGCTCGAATATATGGATTGGGATCTTTAG;INSERTION=ATTCAAGTTCGAAATATGGCAACTTTGAAAGATA;MAPQ=60;MATEID=4503874_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_7815501_7840501_181C;SECONDARY;SPAN=8783;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:97 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:42 DR:116 LR:-415.9 LO:415.9);ALT=G[chr10:7839010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7830256	+	chr10	7840947	+	.	36	0	4503875_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4503875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:7830256(+)-10:7840947(-)__10_7815501_7840501D;SPAN=10691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:36 LR:-115.5 LO:115.5);ALT=A[chr10:7840947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12077479	+	chr10	12084753	+	.	42	0	4514265_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12077479(+)-10:12084753(-)__10_12054001_12079001D;SPAN=7274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:42 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=G[chr10:12084753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12226998	+	chr10	12237766	+	.	33	0	4514964_1	87.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=4514964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12226998(+)-10:12237766(-)__10_12225501_12250501D;SPAN=10768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:80 GQ:87.2 PL:[87.2, 0.0, 107.0] SR:0 DR:33 LR:-87.26 LO:87.37);ALT=A[chr10:12237766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12228331	+	chr10	12237768	+	.	40	12	4514965_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4514965_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_12225501_12250501_423C;SPAN=9437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:89 GQ:94.7 PL:[121.1, 0.0, 94.7] SR:12 DR:40 LR:-121.3 LO:121.3);ALT=C[chr10:12237768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12238316	+	chr10	12251963	+	.	31	0	4514990_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514990_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12238316(+)-10:12251963(-)__10_12225501_12250501D;SPAN=13647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=G[chr10:12251963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12560473	+	chr10	12562974	+	.	79	58	4516315_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTTATTCATTCTT;MAPQ=60;MATEID=4516315_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_10_12544001_12569001_147C;SPAN=2501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:35 GQ:27 PL:[297.0, 27.0, 0.0] SR:58 DR:79 LR:-297.1 LO:297.1);ALT=T[chr10:12562974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	22605485	+	chr10	22606809	+	.	35	27	4541158_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTAG;MAPQ=60;MATEID=4541158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_22589001_22614001_239C;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:68 GQ:17.9 PL:[146.6, 0.0, 17.9] SR:27 DR:35 LR:-152.4 LO:152.4);ALT=G[chr10:22606809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26999048	+	chr10	27002154	+	.	89	35	4551675_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=GAGGTTGCAGTGAGCCGAGATCACGCCATTGCA;MAPQ=0;MATEID=4551675_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_26999001_27024001_99C;SECONDARY;SPAN=3106;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:35 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:35 DR:89 LR:-320.2 LO:320.2);ALT=A[chr10:27002154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27112237	+	chr10	27149675	+	.	32	26	4552106_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4552106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_27146001_27171001_69C;SPAN=37438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:26 DR:32 LR:-128.7 LO:128.7);ALT=G[chr10:27149675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27224203	+	chr10	27228086	+	.	107	79	4552299_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=4552299_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_10_27219501_27244501_51C;SPAN=3883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:51 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:79 DR:107 LR:-445.6 LO:445.6);ALT=A[chr10:27228086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	30723677	+	chr10	30727844	+	.	38	3	4561932_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4561932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_30723001_30748001_156C;SPAN=4167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:98 GQ:99 PL:[108.8, 0.0, 128.6] SR:3 DR:38 LR:-108.8 LO:108.9);ALT=G[chr10:30727844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	31443368	+	chr10	31444865	+	.	77	42	4564183_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=TTGGGAGGCTGAGGCAGG;MAPQ=60;MATEID=4564183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_31433501_31458501_235C;SPAN=1497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:51 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:42 DR:77 LR:-277.3 LO:277.3);ALT=G[chr10:31444865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	35248436	+	chr10	35255023	+	.	90	52	4571671_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4571671_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_10_35255501_35280501_292C;SPAN=6587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:0 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:52 DR:90 LR:-326.8 LO:326.8);ALT=G[chr10:35255023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	42809246	+	chr10	42805768	+	.	40	0	4580853_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4580853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42805768(-)-10:42809246(+)__10_42801501_42826501D;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:70 GQ:56.9 PL:[113.0, 0.0, 56.9] SR:0 DR:40 LR:-114.1 LO:114.1);ALT=]chr10:42809246]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	43892044	+	chr10	43903163	+	.	31	0	4582649_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4582649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43892044(+)-10:43903163(-)__10_43879501_43904501D;SPAN=11119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:48 GQ:26.6 PL:[89.3, 0.0, 26.6] SR:0 DR:31 LR:-91.16 LO:91.16);ALT=A[chr10:43903163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	60477422	+	chr12	72667074	-	G	34	69	5244021_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=5244021_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_72642501_72667501_147C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:57 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:69 DR:34 LR:-280.6 LO:280.6);ALT=G]chr12:72667074];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	61361964	+	chr10	61365009	+	.	47	29	4608151_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AATCA;MAPQ=60;MATEID=4608151_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_61348001_61373001_127C;SPAN=3045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:16 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:29 DR:47 LR:-184.8 LO:184.8);ALT=A[chr10:61365009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70091992	+	chr10	70096955	+	.	55	14	4620900_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4620900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70070001_70095001_81C;SPAN=4963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:29 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:14 DR:55 LR:-184.8 LO:184.8);ALT=G[chr10:70096955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70716068	+	chr10	70719560	+	.	56	32	4622304_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4622304_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70707001_70732001_245C;SPAN=3492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:73 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:32 DR:56 LR:-214.6 LO:214.6);ALT=G[chr10:70719560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70847994	+	chr10	70856838	+	.	128	42	4622876_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4622876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70854001_70879001_121C;SPAN=8844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:142 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:42 DR:128 LR:-419.2 LO:419.2);ALT=T[chr10:70856838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72645038	+	chr10	72648286	+	.	43	0	4625960_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4625960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:72645038(+)-10:72648286(-)__10_72642501_72667501D;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:73 GQ:53 PL:[122.3, 0.0, 53.0] SR:0 DR:43 LR:-123.5 LO:123.5);ALT=T[chr10:72648286[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72645687	+	chr10	72648287	+	.	55	8	4625962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4625962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_72642501_72667501_263C;SPAN=2600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:83 GQ:23.9 PL:[175.7, 0.0, 23.9] SR:8 DR:55 LR:-182.0 LO:182.0);ALT=C[chr10:72648287[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73521785	+	chr10	73533113	+	.	137	78	4627482_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4627482_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73500001_73525001_60C;SPAN=11328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:173 DP:45 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:78 DR:137 LR:-511.6 LO:511.6);ALT=T[chr10:73533113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73594317	+	chr10	73610945	+	.	60	0	4627819_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4627819_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73594317(+)-10:73610945(-)__10_73598001_73623001D;SPAN=16628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:44 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=C[chr10:73610945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975946	+	chr10	73983639	+	.	71	0	4628454_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4628454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73975946(+)-10:73983639(-)__10_73965501_73990501D;SPAN=7693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:58 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=T[chr10:73983639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975992	+	chr10	73992757	+	.	33	0	4628455_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4628455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73975992(+)-10:73992757(-)__10_73965501_73990501D;SPAN=16765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:39 GQ:3.9 PL:[102.3, 3.9, 0.0] SR:0 DR:33 LR:-105.5 LO:105.5);ALT=T[chr10:73992757[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	32673414	+	chr10	74767593	+	AAACATAACACCTAGATACATCC	42	83	6372196_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=AAACATAACACCTAGATACATCC;MAPQ=60;MATEID=6372196_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_17_32658501_32683501_14C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:25 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:83 DR:42 LR:-340.0 LO:340.0);ALT=]chr17:32673414]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	74767593	-	chr17	32673409	+	ATACATCC	44	67	6372195_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;INSERTION=ATACATCC;MAPQ=57;MATEID=6372195_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_32658501_32683501_57C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:23 GQ:27 PL:[297.0, 27.0, 0.0] SR:67 DR:44 LR:-297.1 LO:297.1);ALT=[chr17:32673409[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	75158173	+	chr10	75173768	+	.	76	0	4630725_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4630725_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:75158173(+)-10:75173768(-)__10_75166001_75191001D;SPAN=15595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:55 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:0 DR:76 LR:-224.5 LO:224.5);ALT=T[chr10:75173768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78255578	+	chr10	78261020	+	.	42	36	4635628_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCAGT;MAPQ=60;MATEID=4635628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_78253001_78278001_187C;SPAN=5442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:18 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:36 DR:42 LR:-178.2 LO:178.2);ALT=T[chr10:78261020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78346604	+	chr10	78351578	+	.	53	25	4636083_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAATACTTAATTT;MAPQ=60;MATEID=4636083_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_78351001_78376001_169C;SPAN=4974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:10 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:25 DR:53 LR:-184.8 LO:184.8);ALT=T[chr10:78351578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	79184909	+	chr22	44376043	-	.	31	33	7319557_1	99.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=ATGGATGGATGGATGGATGGATGGATG;MAPQ=25;MATEID=7319557_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_44369501_44394501_144C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:86 GQ:52.7 PL:[155.0, 0.0, 52.7] SR:33 DR:31 LR:-157.6 LO:157.6);ALT=G]chr22:44376043];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	79793707	+	chr10	79795266	+	.	113	0	4638092_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4638092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:79793707(+)-10:79795266(-)__10_79772001_79797001D;SPAN=1559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:113 DP:146 GQ:20 PL:[333.5, 0.0, 20.0] SR:0 DR:113 LR:-349.9 LO:349.9);ALT=C[chr10:79795266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	84127819	+	chr10	84130365	+	.	32	33	4645094_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTC;MAPQ=60;MATEID=4645094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_84108501_84133501_213C;SPAN=2546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:17 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:33 DR:32 LR:-161.7 LO:161.7);ALT=C[chr10:84130365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104184552	+	chr10	104192283	+	AGGTCGGCCTCCGGGAGGTGTGTCTGGACAAAGGCAAGGAGGGCTGCACTGACGATCCTCTCCAGCTCCATGCTCTCTCTT	66	32	4677795_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=AGGTCGGCCTCCGGGAGGTGTGTCTGGACAAAGGCAAGGAGGGCTGCACTGACGATCCTCTCCAGCTCCATGCTCTCTCTT;MAPQ=60;MATEID=4677795_2;MATENM=0;NM=88;NUMPARTS=3;SCTG=c_10_104174001_104199001_158C;SPAN=7731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:71 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:32 DR:66 LR:-227.8 LO:227.8);ALT=G[chr10:104192283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105152063	+	chr10	105156165	+	.	55	0	4679884_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=4679884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:105152063(+)-10:105156165(-)__10_105154001_105179001D;SPAN=4102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:85 GQ:46.4 PL:[158.6, 0.0, 46.4] SR:0 DR:55 LR:-161.8 LO:161.8);ALT=A[chr10:105156165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105156166	-	chrX	73393696	+	.	119	6	7450102_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGAATTTGCGGCTTTGGCAG;MAPQ=60;MATEID=7450102_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_23_73377501_73402501_55C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:41 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:6 DR:119 LR:-359.8 LO:359.8);ALT=[chrX:73393696[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	106015030	+	chr10	106019330	+	.	83	58	4681482_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=TCAGG;MAPQ=60;MATEID=4681482_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_10_106011501_106036501_111C;SPAN=4300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:82 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:58 DR:83 LR:-356.5 LO:356.5);ALT=G[chr10:106019330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	126150556	+	chr10	126172705	+	.	31	11	4712009_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4712009_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_126126001_126151001_159C;SPAN=22149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:21 GQ:9 PL:[99.0, 9.0, 0.0] SR:11 DR:31 LR:-99.02 LO:99.02);ALT=G[chr10:126172705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127191657	+	chr10	127197235	+	.	81	55	4713856_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=4713856_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_169C;SPAN=5578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:47 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:55 DR:81 LR:-323.5 LO:323.5);ALT=C[chr10:127197235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	129060203	+	chr10	129058857	+	.	34	0	4716743_1	93.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=4716743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:129058857(-)-10:129060203(+)__10_129041501_129066501D;SPAN=1346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:69 GQ:73.7 PL:[93.5, 0.0, 73.7] SR:0 DR:34 LR:-93.66 LO:93.66);ALT=]chr10:129060203]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	131265562	+	chr10	131334504	+	.	63	9	4720138_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=4720138_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_131320001_131345001_266C;SPAN=68942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:31 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:9 DR:63 LR:-201.3 LO:201.3);ALT=T[chr10:131334504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131265613	+	chr10	131506157	+	.	60	0	4719939_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4719939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:131265613(+)-10:131506157(-)__10_131246501_131271501D;SPAN=240544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:25 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=A[chr10:131506157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	132909062	+	chr10	132912780	+	.	48	33	4722583_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCA;MAPQ=60;MATEID=4722583_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_132912501_132937501_31C;SPAN=3718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:11 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:33 DR:48 LR:-204.7 LO:204.7);ALT=A[chr10:132912780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	13023198	+	chr18	53590863	-	.	40	48	4764331_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CATTAGATTCTCATAAGGAGCATGCAGCCTAG;MAPQ=60;MATEID=4764331_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_11_13009501_13034501_28C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:24 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:48 DR:40 LR:-241.0 LO:241.0);ALT=G]chr18:53590863];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	14539330	+	chr11	14541841	+	.	82	0	4768435_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4768435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:14539330(+)-11:14541841(-)__11_14528501_14553501D;SPAN=2511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:116 GQ:41.3 PL:[239.3, 0.0, 41.3] SR:0 DR:82 LR:-247.1 LO:247.1);ALT=A[chr11:14541841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	22848934	+	chr11	22851256	+	.	31	0	4790244_1	74.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4790244_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:22848934(+)-11:22851256(-)__11_22834001_22859001D;SPAN=2322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:102 GQ:74.9 PL:[74.9, 0.0, 170.6] SR:0 DR:31 LR:-74.7 LO:76.84);ALT=T[chr11:22851256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32605476	+	chr11	32608555	+	.	70	18	4813771_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4813771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_32585001_32610001_63C;SPAN=3079;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:95 GQ:0.8 PL:[228.5, 0.0, 0.8] SR:18 DR:70 LR:-242.1 LO:242.1);ALT=G[chr11:32608555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32605482	+	chr11	32610136	+	.	52	0	4813773_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4813773_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:32605482(+)-11:32610136(-)__11_32585001_32610001D;SPAN=4654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:47 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=T[chr11:32610136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34460626	+	chr11	34470737	+	.	111	48	4819533_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4819533_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_34447001_34472001_46C;SPAN=10111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:124 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:48 DR:111 LR:-399.4 LO:399.4);ALT=G[chr11:34470737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35160917	+	chr11	35198121	+	.	59	53	4821704_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4821704_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35157501_35182501_184C;SPAN=37204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:201 GQ:99 PL:[315.5, 0.0, 170.3] SR:53 DR:59 LR:-317.5 LO:317.5);ALT=G[chr11:35198121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	36300213	+	chr11	36310910	+	.	33	0	4824914_1	95.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4824914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:36300213(+)-11:36310910(-)__11_36309001_36334001D;SPAN=10697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:52 GQ:29 PL:[95.0, 0.0, 29.0] SR:0 DR:33 LR:-96.6 LO:96.6);ALT=C[chr11:36310910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587286	+	chr11	44609022	+	.	35	11	4844335_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4844335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_44590001_44615001_66C;SPAN=21736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:11 DR:35 LR:-120.9 LO:120.9);ALT=G[chr11:44609022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587310	+	chr11	44616190	+	.	59	0	4844390_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4844390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:44587310(+)-11:44616190(-)__11_44614501_44639501D;SPAN=28880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:55 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=G[chr11:44616190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587324	+	chr11	44621707	+	.	36	0	4844391_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4844391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:44587324(+)-11:44621707(-)__11_44614501_44639501D;SPAN=34383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:65 GQ:55.1 PL:[101.3, 0.0, 55.1] SR:0 DR:36 LR:-101.9 LO:101.9);ALT=A[chr11:44621707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45429849	+	chr11	45431614	+	.	73	40	4846777_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCC;MAPQ=60;MATEID=4846777_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_45423001_45448001_5C;SPAN=1765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:23 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:40 DR:73 LR:-290.5 LO:290.5);ALT=C[chr11:45431614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47381644	+	chr11	47399859	+	.	51	0	4852587_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4852587_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:47381644(+)-11:47399859(-)__11_47383001_47408001D;SPAN=18215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:77 GQ:38.6 PL:[147.5, 0.0, 38.6] SR:0 DR:51 LR:-151.0 LO:151.0);ALT=G[chr11:47399859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47600711	+	chr11	47602077	+	GACTGGGCGACCCTCCGTTCTGTTGCTGCCGGTGAGGCGGGAGAGCGCCGGGGCCGACACGCGCC	60	55	4853543_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GACTGGGCGACCCTCCGTTCTGTTGCTGCCGGTGAGGCGGGAGAGCGCCGGGGCCGACACGCGCC;MAPQ=60;MATEID=4853543_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_47579001_47604001_182C;SPAN=1366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:127 DP:106 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:55 DR:60 LR:-376.3 LO:376.3);ALT=G[chr11:47602077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47660605	+	chr11	47663929	+	.	35	30	4853303_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4853303_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47652501_47677501_379C;SPAN=3324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:91 GQ:84.5 PL:[134.0, 0.0, 84.5] SR:30 DR:35 LR:-134.3 LO:134.3);ALT=T[chr11:47663929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	48600858	+	chr11	48604283	+	.	92	72	4856306_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=4856306_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_48583501_48608501_6C;SPAN=3425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:32 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:72 DR:92 LR:-373.0 LO:373.0);ALT=C[chr11:48604283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	48734780	+	chr11	48736949	+	.	58	11	4856572_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=TTCTCAGAAAGCTTCTTTCTAGTTTTTATTTGAAGATATTTCCTTTTT;MAPQ=60;MATEID=4856572_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_11_48730501_48755501_161C;SPAN=2169;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:15 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:11 DR:58 LR:-201.3 LO:201.3);ALT=T[chr11:48736949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57296438	+	chr11	57298129	+	.	32	0	4869172_1	83.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4869172_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57296438(+)-11:57298129(-)__11_57281001_57306001D;SPAN=1691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:80 GQ:83.9 PL:[83.9, 0.0, 110.3] SR:0 DR:32 LR:-83.96 LO:84.15);ALT=T[chr11:57298129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57322144	+	chr11	57335056	+	.	88	0	4869296_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4869296_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57322144(+)-11:57335056(-)__11_57330001_57355001D;SPAN=12912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:55 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:0 DR:88 LR:-260.8 LO:260.8);ALT=T[chr11:57335056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	58594188	+	chr11	58596020	+	.	90	62	4872674_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4872674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_58579501_58604501_80C;SPAN=1832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:30 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:62 DR:90 LR:-369.7 LO:369.7);ALT=T[chr11:58596020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59949216	+	chr11	59950451	+	.	111	16	4875786_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4875786_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59927001_59952001_152C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:114 DP:100 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:16 DR:111 LR:-336.7 LO:336.7);ALT=T[chr11:59950451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60681765	+	chr11	60687155	+	.	40	0	4877513_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4877513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:60681765(+)-11:60687155(-)__11_60686501_60711501D;SPAN=5390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:40 LR:-130.9 LO:130.9);ALT=G[chr11:60687155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61557426	+	chr11	61560024	+	.	87	0	4880064_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4880064_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61557426(+)-11:61560024(-)__11_61544001_61569001D;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:158 GQ:99 PL:[244.4, 0.0, 138.8] SR:0 DR:87 LR:-245.9 LO:245.9);ALT=T[chr11:61560024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61558075	+	chr11	61560027	+	.	36	50	4880068_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4880068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61544001_61569001_50C;SPAN=1952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:191 GQ:99 PL:[209.3, 0.0, 252.2] SR:50 DR:36 LR:-209.0 LO:209.3);ALT=C[chr11:61560027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61841813	+	chr14	81786774	+	C	43	42	5819167_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=5819167_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_81781001_81806001_356C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:32 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:42 DR:43 LR:-221.2 LO:221.2);ALT=G[chr14:81786774[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	62430848	+	chr11	62432600	+	.	31	0	4883105_1	80.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4883105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62430848(+)-11:62432600(-)__11_62426001_62451001D;SPAN=1752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:83 GQ:80 PL:[80.0, 0.0, 119.6] SR:0 DR:31 LR:-79.84 LO:80.32);ALT=C[chr11:62432600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62529157	+	chr11	62530336	+	.	69	0	4883505_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4883505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62529157(+)-11:62530336(-)__11_62524001_62549001D;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:112 GQ:72.2 PL:[197.6, 0.0, 72.2] SR:0 DR:69 LR:-200.5 LO:200.5);ALT=A[chr11:62530336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62555000	+	chr11	62556492	+	.	104	25	4883323_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4883323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62548501_62573501_83C;SPAN=1492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:94 GQ:30 PL:[330.0, 30.0, 0.0] SR:25 DR:104 LR:-330.1 LO:330.1);ALT=G[chr11:62556492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63304400	+	chr11	63312092	+	.	41	0	4885570_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4885570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63304400(+)-11:63312092(-)__11_63283501_63308501D;SPAN=7692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=C[chr11:63312092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63742267	+	chr11	63743696	+	.	138	160	4886969_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4886969_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63724501_63749501_182C;SPAN=1429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:260 DP:248 GQ:70.3 PL:[772.3, 70.3, 0.0] SR:160 DR:138 LR:-772.4 LO:772.4);ALT=G[chr11:63743696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63754008	+	chr11	63755818	+	.	44	0	4887026_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4887026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63754008(+)-11:63755818(-)__11_63749001_63774001D;SPAN=1810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:73 GQ:49.7 PL:[125.6, 0.0, 49.7] SR:0 DR:44 LR:-127.1 LO:127.1);ALT=T[chr11:63755818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63754037	+	chr11	63763998	+	.	35	0	4887027_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4887027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63754037(+)-11:63763998(-)__11_63749001_63774001D;SPAN=9961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:89 GQ:91.4 PL:[91.4, 0.0, 124.4] SR:0 DR:35 LR:-91.42 LO:91.7);ALT=G[chr11:63763998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64085861	+	chr11	64087204	+	.	104	121	4888484_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGGTG;MAPQ=60;MATEID=4888484_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_11_64067501_64092501_370C;SPAN=1343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:180 DP:176 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:121 DR:104 LR:-534.7 LO:534.7);ALT=G[chr11:64087204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64544099	+	chr11	64545834	+	.	111	93	4889559_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4889559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64533001_64558001_3C;SPAN=1735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:160 DP:106 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:93 DR:111 LR:-475.3 LO:475.3);ALT=C[chr11:64545834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64781744	+	chr11	64785836	+	.	114	21	4890441_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=4890441_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_64778001_64803001_34C;SPAN=4092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:88 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:21 DR:114 LR:-356.5 LO:356.5);ALT=T[chr11:64785836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65623714	+	chr11	65625567	+	.	195	41	4893129_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=4893129_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_11_65611001_65636001_75C;SPAN=1853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:218 DP:134 GQ:58.9 PL:[646.9, 58.9, 0.0] SR:41 DR:195 LR:-647.0 LO:647.0);ALT=C[chr11:65625567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65647456	+	chr11	65648875	+	.	68	0	4893284_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893284_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65647456(+)-11:65648875(-)__11_65635501_65660501D;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:116 GQ:87.5 PL:[193.1, 0.0, 87.5] SR:0 DR:68 LR:-195.1 LO:195.1);ALT=G[chr11:65648875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65820009	+	chr11	65822541	+	.	34	0	4893634_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65820009(+)-11:65822541(-)__11_65807001_65832001D;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:99 GQ:85.4 PL:[85.4, 0.0, 154.7] SR:0 DR:34 LR:-85.41 LO:86.51);ALT=A[chr11:65822541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66360771	+	chr11	66366584	+	TTGGAGTTCGCGGTGCAGATGACCTGTCAGAGCTGTGTGGACGCGGTGCGCAAATCCCTGCAAGGGGTGG	77	103	4895588_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CAGGT;INSERTION=TTGGAGTTCGCGGTGCAGATGACCTGTCAGAGCTGTGTGGACGCGGTGCGCAAATCCCTGCAAGGGGTGG;MAPQ=60;MATEID=4895588_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_66346001_66371001_169C;SPAN=5813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:115 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:103 DR:77 LR:-445.6 LO:445.6);ALT=G[chr11:66366584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66711541	+	chr11	66713342	+	.	31	0	4896993_1	89.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4896993_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66711541(+)-11:66713342(-)__11_66689001_66714001D;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=A[chr11:66713342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67250729	+	chr11	67254475	+	.	40	24	4898541_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4898541_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67252501_67277501_92C;SPAN=3746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:59 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:24 DR:40 LR:-174.9 LO:174.9);ALT=G[chr11:67254475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67374547	+	chr11	67375866	+	.	75	30	4898795_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4898795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67350501_67375501_24C;SPAN=1319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:44 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:30 DR:75 LR:-254.2 LO:254.2);ALT=G[chr11:67375866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67798253	+	chr11	67800388	+	.	93	0	4900683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4900683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67798253(+)-11:67800388(-)__11_67791501_67816501D;SPAN=2135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:89 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:93 LR:-274.0 LO:274.0);ALT=G[chr11:67800388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67798276	+	chr11	67799616	+	.	37	0	4900684_1	97.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4900684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67798276(+)-11:67799616(-)__11_67791501_67816501D;SPAN=1340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:91 GQ:97.7 PL:[97.7, 0.0, 120.8] SR:0 DR:37 LR:-97.48 LO:97.65);ALT=G[chr11:67799616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68582956	+	chr11	68609241	+	.	35	6	4903104_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=4903104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68575501_68600501_141C;SPAN=26285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:29 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:6 DR:35 LR:-108.9 LO:108.9);ALT=C[chr11:68609241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68664206	+	chr11	68671189	+	.	31	0	4903530_1	80.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4903530_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68664206(+)-11:68671189(-)__11_68649001_68674001D;SPAN=6983;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:79 GQ:80.9 PL:[80.9, 0.0, 110.6] SR:0 DR:31 LR:-80.93 LO:81.18);ALT=T[chr11:68671189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68665526	+	chr11	68671209	+	.	50	0	4903534_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4903534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68665526(+)-11:68671209(-)__11_68649001_68674001D;SPAN=5683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:82 GQ:53.9 PL:[143.0, 0.0, 53.9] SR:0 DR:50 LR:-144.9 LO:144.9);ALT=G[chr11:68671209[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77340946	+	chr11	77348635	+	.	69	108	4927236_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4927236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77346501_77371501_7C;SPAN=7689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:159 DP:52 GQ:43 PL:[472.0, 43.0, 0.0] SR:108 DR:69 LR:-472.0 LO:472.0);ALT=T[chr11:77348635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77532287	+	chr11	77553524	+	.	37	5	4927615_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4927615_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77542501_77567501_219C;SPAN=21237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:36 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:5 DR:37 LR:-118.8 LO:118.8);ALT=G[chr11:77553524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77784239	+	chr11	77790677	+	.	39	0	4928397_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4928397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:77784239(+)-11:77790677(-)__11_77787501_77812501D;SPAN=6438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:104 GQ:99 PL:[100.7, 0.0, 150.2] SR:0 DR:39 LR:-100.6 LO:101.1);ALT=T[chr11:77790677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111750349	+	chr11	111753087	+	.	34	0	5004468_1	90.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5004468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:111750349(+)-11:111753087(-)__11_111744501_111769501D;SPAN=2738;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:79 GQ:90.8 PL:[90.8, 0.0, 100.7] SR:0 DR:34 LR:-90.83 LO:90.86);ALT=T[chr11:111753087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111956197	+	chr11	111957359	+	.	67	0	5004916_1	99.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5004916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:111956197(+)-11:111957359(-)__11_111940501_111965501D;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:77 GQ:14.1 PL:[214.5, 14.1, 0.0] SR:0 DR:67 LR:-216.8 LO:216.8);ALT=A[chr11:111957359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	112025808	+	chr11	112034629	+	.	55	20	5005082_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=5005082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_112014001_112039001_261C;SPAN=8821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:20 DR:55 LR:-235.6 LO:235.6);ALT=G[chr11:112034629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	122347584	+	chr11	122349281	+	.	79	60	5031365_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAGAAAG;MAPQ=60;MATEID=5031365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_122328501_122353501_261C;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:42 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:60 DR:79 LR:-346.6 LO:346.6);ALT=G[chr11:122349281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	122931522	+	chr11	122932783	+	.	51	0	5033502_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5033502_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:122931522(+)-11:122932783(-)__11_122916501_122941501D;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:224 GQ:99 PL:[107.8, 0.0, 434.6] SR:0 DR:51 LR:-107.7 LO:118.9);ALT=A[chr11:122932783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6041904	+	chr12	6040782	+	.	58	0	5078888_1	99.0	.	DISC_MAPQ=6;EVDNC=DSCRD;IMPRECISE;MAPQ=6;MATEID=5078888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6040782(-)-12:6041904(+)__12_6027001_6052001D;SPAN=1122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:200 GQ:99 PL:[137.3, 0.0, 348.5] SR:0 DR:58 LR:-137.3 LO:142.3);ALT=]chr12:6041904]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	6241438	+	chr12	6248078	+	.	40	49	5079389_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5079389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6247501_6272501_101C;SPAN=6640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:30 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:49 DR:40 LR:-211.3 LO:211.3);ALT=G[chr12:6248078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6309731	+	chr12	6334591	+	.	56	58	5079338_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5079338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6296501_6321501_150C;SPAN=24860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:44 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:58 DR:56 LR:-267.4 LO:267.4);ALT=G[chr12:6334591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6547703	-	chr15	40331293	+	.	116	0	5930665_1	99.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=5930665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6547703(-)-15:40331293(-)__15_40327001_40352001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:70 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:0 DR:116 LR:-343.3 LO:343.3);ALT=[chr15:40331293[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	6644055	+	chr12	6645657	+	.	80	0	5080809_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5080809_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6644055(+)-12:6645657(-)__12_6639501_6664501D;SPAN=1602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:80 DP:119 GQ:56.9 PL:[231.8, 0.0, 56.9] SR:0 DR:80 LR:-237.8 LO:237.8);ALT=T[chr12:6645657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6762600	+	chr12	6772227	+	.	31	0	5081197_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5081197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6762600(+)-12:6772227(-)__12_6737501_6762501D;SPAN=9627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:1 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=G[chr12:6772227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9907908	+	chr12	9913431	+	.	73	0	5090940_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5090940_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:9907908(+)-12:9913431(-)__12_9898001_9923001D;SPAN=5523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:159 GQ:99 PL:[197.9, 0.0, 188.0] SR:0 DR:73 LR:-197.9 LO:197.9);ALT=A[chr12:9913431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9909015	+	chr12	9913353	+	.	111	36	5090943_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5090943_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TACTAC;SCTG=c_12_9898001_9923001_218C;SPAN=4338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:119 DP:166 GQ:33.3 PL:[264.8, 0.0, 33.3] SR:36 DR:111 LR:-276.8 LO:276.8);ALT=T[chr12:9913353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10010572	+	chr12	10021800	+	.	84	0	5091219_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5091219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:10010572(+)-12:10021800(-)__12_10020501_10045501D;SPAN=11228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:53 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=A[chr12:10021800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10124286	+	chr12	10131563	+	.	34	46	5091603_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5091603_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_10118501_10143501_313C;SPAN=7277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:91 GQ:54.8 PL:[163.7, 0.0, 54.8] SR:46 DR:34 LR:-166.3 LO:166.3);ALT=G[chr12:10131563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	12544867	+	chr12	12546626	-	.	44	0	5097666_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5097666_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:12544867(+)-12:12546626(+)__12_12519501_12544501D;SPAN=1759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:0 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:0 DR:44 LR:-128.7 LO:128.7);ALT=C]chr12:12546626];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	21800002	+	chr12	21810684	+	.	103	0	5120205_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5120205_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:21800002(+)-12:21810684(-)__12_21805001_21830001D;SPAN=10682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:77 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:0 DR:103 LR:-303.7 LO:303.7);ALT=A[chr12:21810684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21807612	+	chr12	21810685	+	.	132	33	5120215_1	99.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=C;MAPQ=56;MATEID=5120215_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_21805001_21830001_23C;SPAN=3073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:161 DP:131 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:33 DR:132 LR:-475.3 LO:475.3);ALT=C[chr12:21810685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	25956130	-	chr12	125801147	+	.	36	0	5382534_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=5382534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:25956130(-)-12:125801147(-)__12_125783001_125808001D;SPAN=99845017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:0 DR:36 LR:-112.2 LO:112.2);ALT=[chr12:125801147[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	27863891	+	chr12	27869221	+	.	37	0	5135005_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5135005_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:27863891(+)-12:27869221(-)__12_27856501_27881501D;SPAN=5330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:84 GQ:99 PL:[99.5, 0.0, 102.8] SR:0 DR:37 LR:-99.38 LO:99.39);ALT=G[chr12:27869221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49334973	+	chr12	49351092	+	.	44	21	5181180_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5181180_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_49318501_49343501_364C;SPAN=16119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:43 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:21 DR:44 LR:-161.7 LO:161.7);ALT=T[chr12:49351092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49523522	+	chr12	49525104	+	.	133	0	5182092_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=5182092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49523522(+)-12:49525104(-)__12_49514501_49539501D;SPAN=1582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:89 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:0 DR:133 LR:-392.8 LO:392.8);ALT=A[chr12:49525104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49580617	+	chr12	49582760	+	.	111	23	5182017_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;HOMSEQ=C;MAPQ=0;MATEID=5182017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_49563501_49588501_187C;SPAN=2143;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:127 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:23 DR:111 LR:-376.3 LO:376.3);ALT=C[chr12:49582760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49658948	+	chr12	49663245	+	.	56	0	5182254_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5182254_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49658948(+)-12:49663245(-)__12_49661501_49686501D;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:65 GQ:10.8 PL:[178.2, 10.8, 0.0] SR:0 DR:56 LR:-180.4 LO:180.4);ALT=C[chr12:49663245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50135437	+	chr12	50146749	+	.	59	0	5183524_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5183524_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:50135437(+)-12:50146749(-)__12_50127001_50152001D;SPAN=11312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:89 GQ:45.2 PL:[170.6, 0.0, 45.2] SR:0 DR:59 LR:-174.7 LO:174.7);ALT=G[chr12:50146749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50506085	+	chr12	50513817	+	.	115	14	5184885_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5184885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_50494501_50519501_396C;SPAN=7732;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:123 GQ:33 PL:[363.0, 33.0, 0.0] SR:14 DR:115 LR:-363.1 LO:363.1);ALT=G[chr12:50513817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51632705	+	chr12	51634125	+	.	68	24	5188897_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5188897_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_51621501_51646501_341C;SPAN=1420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:103 GQ:24.3 PL:[297.0, 24.3, 0.0] SR:24 DR:68 LR:-296.7 LO:296.7);ALT=G[chr12:51634125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51632744	+	chr12	51634652	+	.	58	0	5188898_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5188898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:51632744(+)-12:51634652(-)__12_51621501_51646501D;SPAN=1908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:118 GQ:99 PL:[159.5, 0.0, 126.5] SR:0 DR:58 LR:-159.7 LO:159.7);ALT=T[chr12:51634652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53594271	+	chr12	53600982	+	.	36	0	5194260_1	96.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5194260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53594271(+)-12:53600982(-)__12_53581501_53606501D;SPAN=6711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:84 GQ:96.2 PL:[96.2, 0.0, 106.1] SR:0 DR:36 LR:-96.08 LO:96.12);ALT=A[chr12:53600982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53689423	+	chr12	53691631	+	.	48	12	5194794_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=0;MATEID=5194794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53679501_53704501_127C;SECONDARY;SPAN=2208;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:174 GQ:99 PL:[141.2, 0.0, 279.8] SR:12 DR:48 LR:-141.0 LO:143.6);ALT=G[chr12:53691631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53835823	+	chr19	40449669	-	.	43	0	6815630_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6815630_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53835823(+)-19:40449669(+)__19_40449501_40474501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:34 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=C]chr19:40449669];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	53846160	+	chr12	53848508	+	.	36	71	5195674_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5195674_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_12_53826501_53851501_26C;SPAN=2348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:121 DP:197 GQ:99 PL:[346.1, 0.0, 131.6] SR:71 DR:36 LR:-351.3 LO:351.3);ALT=G[chr12:53848508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54063128	+	chr12	54066356	+	.	47	0	5196112_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5196112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54063128(+)-12:54066356(-)__12_54047001_54072001D;SPAN=3228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:102 GQ:99 PL:[127.7, 0.0, 117.8] SR:0 DR:47 LR:-127.5 LO:127.5);ALT=G[chr12:54066356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54719017	+	chr12	54737008	+	.	32	0	5198486_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5198486_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54719017(+)-12:54737008(-)__12_54708501_54733501D;SPAN=17991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:32 LR:-102.3 LO:102.3);ALT=G[chr12:54737008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56110415	+	chr12	56112873	+	.	81	0	5201743_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5201743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56110415(+)-12:56112873(-)__12_56105001_56130001D;SPAN=2458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:125 GQ:68.6 PL:[233.6, 0.0, 68.6] SR:0 DR:81 LR:-238.4 LO:238.4);ALT=T[chr12:56112873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56121170	+	chr12	56122734	+	.	117	0	5201784_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5201784_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56121170(+)-12:56122734(-)__12_56105001_56130001D;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:106 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:0 DR:117 LR:-346.6 LO:346.6);ALT=G[chr12:56122734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56194736	+	chr12	56211447	+	.	40	0	5202113_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=5202113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56194736(+)-12:56211447(-)__12_56203001_56228001D;SPAN=16711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:68 GQ:50.9 PL:[113.6, 0.0, 50.9] SR:0 DR:40 LR:-114.9 LO:114.9);ALT=T[chr12:56211447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56552242	+	chr12	56553365	+	.	89	0	5203588_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5203588_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56552242(+)-12:56553365(-)__12_56546001_56571001D;SPAN=1123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:116 GQ:18.2 PL:[262.4, 0.0, 18.2] SR:0 DR:89 LR:-274.8 LO:274.8);ALT=G[chr12:56553365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56552242	+	chr12	56553757	+	.	53	0	5203589_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5203589_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56552242(+)-12:56553757(-)__12_56546001_56571001D;SPAN=1515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:135 GQ:99 PL:[138.5, 0.0, 188.0] SR:0 DR:53 LR:-138.4 LO:138.8);ALT=G[chr12:56553757[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57066858	+	chr12	57081845	+	.	45	0	5205323_1	98.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5205323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57066858(+)-12:57081845(-)__12_57060501_57085501D;SPAN=14987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:184 GQ:98.9 PL:[98.9, 0.0, 346.4] SR:0 DR:45 LR:-98.7 LO:106.5);ALT=G[chr12:57081845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57911588	+	chr12	57914200	+	.	42	0	5208090_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5208090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57911588(+)-12:57914200(-)__12_57893501_57918501D;SPAN=2612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:66 GQ:38.3 PL:[120.8, 0.0, 38.3] SR:0 DR:42 LR:-123.0 LO:123.0);ALT=C[chr12:57914200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57929679	+	chr12	57940856	+	.	37	0	5207876_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5207876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57929679(+)-12:57940856(-)__12_57918001_57943001D;SPAN=11177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:110 GQ:92.3 PL:[92.3, 0.0, 174.8] SR:0 DR:37 LR:-92.34 LO:93.73);ALT=A[chr12:57940856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	62654287	+	chr12	62687959	+	.	48	14	5218937_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTA;MAPQ=60;MATEID=5218937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_62671001_62696001_165C;SPAN=33672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:33 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:14 DR:48 LR:-151.8 LO:151.8);ALT=A[chr12:62687959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66527651	+	chr12	66529877	+	.	70	36	5229088_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATGGTATTAATA;MAPQ=60;MATEID=5229088_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_66517501_66542501_131C;SPAN=2226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:30 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:36 DR:70 LR:-257.5 LO:257.5);ALT=A[chr12:66529877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66546210	+	chr12	66563674	+	.	42	0	5229007_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5229007_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:66546210(+)-12:66563674(-)__12_66542001_66567001D;SPAN=17464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:85 GQ:89.3 PL:[115.7, 0.0, 89.3] SR:0 DR:42 LR:-115.8 LO:115.8);ALT=T[chr12:66563674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66547229	+	chr12	66563635	+	.	50	16	5229008_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5229008_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_66542001_66567001_87C;SPAN=16406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:75 GQ:19.4 PL:[161.3, 0.0, 19.4] SR:16 DR:50 LR:-167.5 LO:167.5);ALT=C[chr12:66563635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69633487	+	chr12	69644906	+	.	34	6	5236722_1	98.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5236722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69629001_69654001_357C;SPAN=11419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:87 GQ:98.6 PL:[98.6, 0.0, 111.8] SR:6 DR:34 LR:-98.57 LO:98.62);ALT=G[chr12:69644906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69742325	+	chr12	69743888	+	.	121	189	5237477_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5237477_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_69727001_69752001_255C;SPAN=1563;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:271 DP:364 GQ:86.4 PL:[796.1, 0.0, 86.4] SR:189 DR:121 LR:-829.0 LO:829.0);ALT=G[chr12:69743888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69979351	+	chr12	69980529	+	.	38	0	5237729_1	98.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5237729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69979351(+)-12:69980529(-)__12_69972001_69997001D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:98 GQ:98.9 PL:[98.9, 0.0, 138.5] SR:0 DR:38 LR:-98.89 LO:99.26);ALT=C[chr12:69980529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70594864	+	chr12	70597578	+	.	63	36	5239429_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAAGTATGACACTTC;MAPQ=60;MATEID=5239429_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_70584501_70609501_34C;SPAN=2714;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:56 GQ:21 PL:[231.0, 21.0, 0.0] SR:36 DR:63 LR:-231.1 LO:231.1);ALT=C[chr12:70597578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	71602361	+	chr12	71604474	+	.	40	26	5241454_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TACT;MAPQ=60;MATEID=5241454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_71589001_71614001_136C;SPAN=2113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:43 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:26 DR:40 LR:-151.8 LO:151.8);ALT=T[chr12:71604474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	73239578	+	chr15	94888547	-	.	71	39	6044574_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=6044574_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_94864001_94889001_17C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:40 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:39 DR:71 LR:-293.8 LO:293.8);ALT=G]chr15:94888547];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	76462802	+	chr12	76478346	+	.	42	0	5252619_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=5252619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76462802(+)-12:76478346(-)__12_76440001_76465001D;SPAN=15544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:30 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=T[chr12:76478346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	82139719	+	chr12	82144320	+	.	31	17	5265170_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AACA;MAPQ=60;MATEID=5265170_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_82124001_82149001_249C;SPAN=4601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:69 GQ:50.6 PL:[116.6, 0.0, 50.6] SR:17 DR:31 LR:-118.1 LO:118.1);ALT=A[chr12:82144320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	89172969	+	chr12	89184607	+	G	53	33	5280301_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=5280301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_89180001_89205001_73C;SPAN=11638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:21 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:33 DR:53 LR:-214.6 LO:214.6);ALT=A[chr12:89184607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112451340	+	chr12	112457557	+	.	44	0	5341325_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5341325_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112451340(+)-12:112457557(-)__12_112430501_112455501D;SPAN=6217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:54 GQ:1.2 PL:[132.0, 1.2, 0.0] SR:0 DR:44 LR:-138.6 LO:138.6);ALT=T[chr12:112457557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112451340	+	chr20	50727569	-	.	64	0	5341326_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5341326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112451340(+)-20:50727569(+)__12_112430501_112455501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:54 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=T]chr20:50727569];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	113019463	+	chr12	113020507	+	.	36	0	5343078_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5343078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:113019463(+)-12:113020507(-)__12_113018501_113043501D;SPAN=1044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:54 GQ:25.1 PL:[104.3, 0.0, 25.1] SR:0 DR:36 LR:-106.8 LO:106.8);ALT=C[chr12:113020507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	87426048	+	chr12	117013730	+	.	94	0	5353875_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=5353875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:117013730(-)-16:87426048(+)__12_117012001_117037001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:57 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:0 DR:94 LR:-277.3 LO:277.3);ALT=]chr16:87426048]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	117086884	+	chr12	117088194	+	.	53	28	5354127_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGTGGCTCAGGCCTATAATCCCAGCACTT;MAPQ=60;MATEID=5354127_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_12_117085501_117110501_183C;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:35 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:28 DR:53 LR:-217.9 LO:217.9);ALT=T[chr12:117088194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120934030	+	chr12	120935873	+	.	41	0	5365557_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5365557_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:120934030(+)-12:120935873(-)__12_120932001_120957001D;SPAN=1843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:92 GQ:99 PL:[110.6, 0.0, 110.6] SR:0 DR:41 LR:-110.4 LO:110.4);ALT=C[chr12:120935873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121163734	+	chr12	121164827	+	.	37	9	5366604_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5366604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121152501_121177501_365C;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:78 GQ:87.8 PL:[101.0, 0.0, 87.8] SR:9 DR:37 LR:-101.0 LO:101.0);ALT=G[chr12:121164827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123006847	+	chr12	123011394	+	.	31	10	5373036_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5373036_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122990001_123015001_65C;SPAN=4547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:101 GQ:85.1 PL:[85.1, 0.0, 157.7] SR:10 DR:31 LR:-84.87 LO:86.14);ALT=C[chr12:123011394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124069363	+	chr12	124071292	+	.	31	57	5376855_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5376855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124068001_124093001_292C;SPAN=1929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:116 GQ:80.9 PL:[199.7, 0.0, 80.9] SR:57 DR:31 LR:-202.3 LO:202.3);ALT=G[chr12:124071292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	131131938	+	chr12	131133868	+	.	90	59	5396285_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=5396285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_131124001_131149001_414C;SPAN=1930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:32 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:59 DR:90 LR:-379.6 LO:379.6);ALT=C[chr12:131133868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133175151	+	chr12	133174003	+	.	32	0	5401927_1	87.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5401927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:133174003(-)-12:133175151(+)__12_133157501_133182501D;SPAN=1148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:68 GQ:77.3 PL:[87.2, 0.0, 77.3] SR:0 DR:32 LR:-87.24 LO:87.24);ALT=]chr12:133175151]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	46733823	+	chr13	46756246	+	.	72	18	5483770_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5483770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46721501_46746501_155C;SPAN=22423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:48 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:18 DR:72 LR:-237.7 LO:237.7);ALT=T[chr13:46756246[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47361294	+	chr13	47371239	+	.	79	0	5485768_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5485768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:47361294(+)-13:47371239(-)__13_47358501_47383501D;SPAN=9945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:125 GQ:75.2 PL:[227.0, 0.0, 75.2] SR:0 DR:79 LR:-231.0 LO:231.0);ALT=A[chr13:47371239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47365603	+	chr13	47371239	+	.	42	0	5485783_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5485783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:47365603(+)-13:47371239(-)__13_47358501_47383501D;SPAN=5636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:118 GQ:99 PL:[106.7, 0.0, 179.3] SR:0 DR:42 LR:-106.7 LO:107.7);ALT=A[chr13:47371239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51069350	+	chr13	51075079	+	.	103	63	5496294_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCTC;MAPQ=60;MATEID=5496294_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_51058001_51083001_85C;SPAN=5729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:33 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:63 DR:103 LR:-402.7 LO:402.7);ALT=C[chr13:51075079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51484620	+	chr13	51503593	+	.	35	0	5497401_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5497401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:51484620(+)-13:51503593(-)__13_51474501_51499501D;SPAN=18973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:35 LR:-115.2 LO:115.2);ALT=T[chr13:51503593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	31789766	-	chr17	46972515	+	.	75	0	6420812_1	99.0	.	DISC_MAPQ=5;EVDNC=DSCRD;IMPRECISE;MAPQ=5;MATEID=6420812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:31789766(-)-17:46972515(-)__17_46966501_46991501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:55 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:0 DR:75 LR:-221.2 LO:221.2);ALT=[chr17:46972515[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	32953311	+	chr14	32954349	+	.	39	0	5695354_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5695354_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:32953311(+)-14:32954349(-)__14_32952501_32977501D;SPAN=1038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:5 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:39 LR:-115.5 LO:115.5);ALT=T[chr14:32954349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35761736	+	chr14	35777196	+	.	33	0	5702629_1	96.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5702629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35761736(+)-14:35777196(-)__14_35770001_35795001D;SPAN=15460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:47 GQ:17 PL:[96.2, 0.0, 17.0] SR:0 DR:33 LR:-99.25 LO:99.25);ALT=C[chr14:35777196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	44248335	+	chr14	43824277	+	.	64	66	5722667_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAT;MAPQ=60;MATEID=5722667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_44247001_44272001_22C;SPAN=424058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:50 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:66 DR:64 LR:-303.7 LO:303.7);ALT=]chr14:44248335]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	45716582	+	chr14	45722236	+	.	38	10	5726228_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5726228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_45717001_45742001_332C;SPAN=5654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:10 DR:38 LR:-141.4 LO:141.4);ALT=T[chr14:45722236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	47117868	-	chr14	63226284	+	.	40	32	5729177_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=A;MAPQ=0;MATEID=5729177_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GGG;SCTG=c_14_47113501_47138501_134C;SECONDARY;SPAN=16108416;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:51 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:32 DR:40 LR:-191.4 LO:191.4);ALT=[chr14:63226284[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	49331368	+	chr14	49333935	+	.	92	82	5733830_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GCT;MAPQ=60;MATEID=5733830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_49318501_49343501_217C;SPAN=2567;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:40 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:82 DR:92 LR:-415.9 LO:415.9);ALT=T[chr14:49333935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	52456418	+	chr14	52458033	+	.	71	75	5742362_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5742362_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_52454501_52479501_323C;SPAN=1615;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:104 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:75 DR:71 LR:-389.5 LO:389.5);ALT=G[chr14:52458033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54710349	+	chr14	54713686	+	.	90	61	5748017_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGA;MAPQ=60;MATEID=5748017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54708501_54733501_165C;SPAN=3337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:33 GQ:33 PL:[363.0, 33.0, 0.0] SR:61 DR:90 LR:-363.1 LO:363.1);ALT=A[chr14:54713686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54897171	+	chr14	54907992	+	.	33	0	5748494_1	95.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5748494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54897171(+)-14:54907992(-)__14_54904501_54929501D;SPAN=10821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:48 GQ:20 PL:[95.9, 0.0, 20.0] SR:0 DR:33 LR:-98.67 LO:98.67);ALT=C[chr14:54907992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54898987	+	chr14	54907989	+	.	66	0	5748495_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5748495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54898987(+)-14:54907989(-)__14_54904501_54929501D;SPAN=9002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:42 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:0 DR:66 LR:-194.7 LO:194.7);ALT=A[chr14:54907989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54903155	+	chr14	54907965	+	.	36	23	5748496_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5748496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54904501_54929501_119C;SPAN=4810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:28 GQ:12 PL:[132.0, 12.0, 0.0] SR:23 DR:36 LR:-132.0 LO:132.0);ALT=T[chr14:54907965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55596062	+	chr14	55604760	+	.	51	0	5750397_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5750397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55596062(+)-14:55604760(-)__14_55590501_55615501D;SPAN=8698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:74 GQ:29.6 PL:[148.4, 0.0, 29.6] SR:0 DR:51 LR:-152.6 LO:152.6);ALT=G[chr14:55604760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56047074	+	chr14	56078736	+	.	40	16	5752052_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5752052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56056001_56081001_199C;SPAN=31662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:39 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:16 DR:40 LR:-148.5 LO:148.5);ALT=T[chr14:56078736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58711659	+	chr14	58718835	+	TATGACCTGTCAGCCTCTACATTCTCTCCTGACGGAAGAGTTTTTCAAGTTGAATATGCTATGAAGGCTGTGGAAAATAGT	41	22	5758570_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TATGACCTGTCAGCCTCTACATTCTCTCCTGACGGAAGAGTTTTTCAAGTTGAATATGCTATGAAGGCTGTGGAAAATAGT;MAPQ=60;MATEID=5758570_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_58702001_58727001_369C;SPAN=7176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:82 GQ:50.6 PL:[146.3, 0.0, 50.6] SR:22 DR:41 LR:-148.5 LO:148.5);ALT=G[chr14:58718835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65360396	+	chr14	65363541	+	.	76	52	5775303_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGAATTTTC;MAPQ=60;MATEID=5775303_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_14_65341501_65366501_300C;SPAN=3145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:33 GQ:27 PL:[297.0, 27.0, 0.0] SR:52 DR:76 LR:-297.1 LO:297.1);ALT=C[chr14:65363541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381253	+	chr14	65390708	+	.	87	8	5775401_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5775401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65390501_65415501_359C;SPAN=9455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:40 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:8 DR:87 LR:-267.4 LO:267.4);ALT=G[chr14:65390708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381279	+	chr14	65398853	+	.	36	0	5775402_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5775402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65381279(+)-14:65398853(-)__14_65390501_65415501D;SPAN=17574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:59 GQ:40.1 PL:[102.8, 0.0, 40.1] SR:0 DR:36 LR:-104.3 LO:104.3);ALT=C[chr14:65398853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381282	+	chr14	65392724	+	.	50	0	5775403_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5775403_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65381282(+)-14:65392724(-)__14_65390501_65415501D;SPAN=11442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:50 LR:-161.7 LO:161.7);ALT=G[chr14:65392724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	69853826	+	chr14	69864946	+	.	65	0	5786822_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=5786822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:69853826(+)-14:69864946(-)__14_69849501_69874501D;SPAN=11120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:114 GQ:91.4 PL:[183.8, 0.0, 91.4] SR:0 DR:65 LR:-185.3 LO:185.3);ALT=A[chr14:69864946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70796006	+	chr14	70826238	+	.	33	0	5789243_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5789243_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:70796006(+)-14:70826238(-)__14_70805001_70830001D;SPAN=30232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:61 GQ:53 PL:[92.6, 0.0, 53.0] SR:0 DR:33 LR:-92.9 LO:92.9);ALT=A[chr14:70826238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70809487	+	chr14	70826295	+	.	40	0	5789253_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5789253_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:70809487(+)-14:70826295(-)__14_70805001_70830001D;SPAN=16808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:97 GQ:99 PL:[105.8, 0.0, 128.9] SR:0 DR:40 LR:-105.8 LO:105.9);ALT=C[chr14:70826295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73525413	+	chr14	73538334	+	.	44	26	5795961_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5795961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73524501_73549501_277C;SPAN=12921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:96 GQ:79.7 PL:[152.3, 0.0, 79.7] SR:26 DR:44 LR:-153.4 LO:153.4);ALT=G[chr14:73538334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	90863578	+	chr14	90867602	+	CTGATCAGCTGACCGAAGAACAGATTGCT	39	211	5839807_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CTGATCAGCTGACCGAAGAACAGATTGCT;MAPQ=60;MATEID=5839807_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_90846001_90871001_177C;SPAN=4024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:232 DP:135 GQ:62.5 PL:[686.5, 62.5, 0.0] SR:211 DR:39 LR:-686.6 LO:686.6);ALT=G[chr14:90867602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	94546110	+	chr14	94547464	+	.	50	0	5850020_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5850020_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:94546110(+)-14:94547464(-)__14_94521001_94546001D;SPAN=1354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:0 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=T[chr14:94547464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	103800934	+	chr14	103801989	+	.	32	37	5874493_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5874493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_103782001_103807001_337C;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:37 DR:32 LR:-163.7 LO:163.7);ALT=G[chr14:103801989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104379095	+	chr14	104387803	+	.	75	0	5876590_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5876590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:104379095(+)-14:104387803(-)__14_104370001_104395001D;SPAN=8708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:176 GQ:99 PL:[200.0, 0.0, 226.4] SR:0 DR:75 LR:-199.9 LO:200.0);ALT=A[chr14:104387803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104381528	+	chr14	104387807	+	.	62	3	5876599_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5876599_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_104370001_104395001_319C;SPAN=6279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:241 GQ:99 PL:[146.2, 0.0, 436.7] SR:3 DR:62 LR:-146.0 LO:154.1);ALT=T[chr14:104387807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105219656	+	chr14	105221966	+	.	115	62	5878785_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5878785_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_105203001_105228001_34C;SPAN=2310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:81 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:62 DR:115 LR:-422.5 LO:422.5);ALT=G[chr14:105221966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105391327	+	chr14	105393476	+	.	45	9	5879068_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5879068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_105374501_105399501_235C;SPAN=2149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:87 GQ:55.7 PL:[154.7, 0.0, 55.7] SR:9 DR:45 LR:-157.2 LO:157.2);ALT=G[chr14:105393476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105417220	+	chr14	105418257	+	.	31	0	5879124_1	92.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5879124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105417220(+)-14:105418257(-)__14_105399001_105424001D;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=A[chr14:105418257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106227280	+	chr14	106082685	+	AC	35	63	5882176_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AC;MAPQ=35;MATEID=5882176_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_14_106207501_106232501_108C;SPAN=144595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:107 GQ:7.4 PL:[251.6, 0.0, 7.4] SR:63 DR:35 LR:-265.4 LO:265.4);ALT=]chr14:106227280]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106115778	+	chr14	106096963	+	.	84	0	5881616_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5881616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106096963(-)-14:106115778(+)__14_106085001_106110001D;SPAN=18815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:49 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=]chr14:106115778]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106346009	+	chr14	106386922	+	.	41	6	5882731_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=5882731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106379001_106404001_249C;SPAN=40913;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:56 GQ:8 PL:[126.8, 0.0, 8.0] SR:6 DR:41 LR:-132.8 LO:132.8);ALT=A[chr14:106386922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106374811	+	chr14	106386920	+	.	36	8	5882739_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5882739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106379001_106404001_2C;SPAN=12109;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:53 GQ:0.9 PL:[128.7, 0.9, 0.0] SR:8 DR:36 LR:-135.3 LO:135.3);ALT=G[chr14:106386920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	23671438	+	chr15	23675199	+	.	39	11	5901087_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=GGCACGGTGGCTCACGCCTGTAATCCCAGCACTTTGGGAGGCCAAGG;MAPQ=60;MATEID=5901087_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_23667001_23692001_111C;SPAN=3761;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:77 GQ:45.2 PL:[140.9, 0.0, 45.2] SR:11 DR:39 LR:-143.5 LO:143.5);ALT=G[chr15:23675199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	35529517	-	chr15	69113095	+	.	32	0	5979459_1	93.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5979459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:35529517(-)-15:69113095(-)__15_69090001_69115001D;SPAN=33583578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:44 GQ:11.3 PL:[93.8, 0.0, 11.3] SR:0 DR:32 LR:-97.22 LO:97.22);ALT=[chr15:69113095[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	39372395	+	chr15	39373461	+	.	43	34	5929389_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=TTCTCCTGCCTCAGCCTCCCGAGTAGCTGGGATTACAGGCA;MAPQ=60;MATEID=5929389_2;MATENM=5;NM=1;NUMPARTS=2;SCTG=c_15_39371501_39396501_138C;SPAN=1066;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:6 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:34 DR:43 LR:-221.2 LO:221.2);ALT=A[chr15:39373461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41576309	+	chr15	41577421	+	.	40	14	5933342_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5933342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41576501_41601501_263C;SPAN=1112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:31 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:14 DR:40 LR:-135.3 LO:135.3);ALT=G[chr15:41577421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41709512	+	chr15	41730517	+	.	44	56	5933821_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5933821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41699001_41724001_208C;SPAN=21005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:38 GQ:18 PL:[198.0, 18.0, 0.0] SR:56 DR:44 LR:-198.0 LO:198.0);ALT=G[chr15:41730517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	44084833	+	chr15	44085888	+	.	209	0	5938738_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5938738_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:44084833(+)-15:44085888(-)__15_44075501_44100501D;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:209 DP:77 GQ:56.5 PL:[620.5, 56.5, 0.0] SR:0 DR:209 LR:-620.6 LO:620.6);ALT=G[chr15:44085888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45927306	+	chr15	45951104	+	.	46	4	5942278_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5942278_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_15_45913001_45938001_146C;SPAN=23798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:4 DR:46 LR:-138.6 LO:138.6);ALT=G[chr15:45951104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55485033	+	chr15	55489006	+	.	79	49	5956087_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=23;MATEID=5956087_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_55468001_55493001_269C;SPAN=3973;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:85 GQ:27 PL:[297.0, 27.0, 0.0] SR:49 DR:79 LR:-297.1 LO:297.1);ALT=T[chr15:55489006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34188507	+	chr15	55489006	+	.	40	26	5956092_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5956092_2;MATENM=4;NM=0;NUMPARTS=2;REPSEQ=CC;SCTG=c_15_55468001_55493001_269C;SECONDARY;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:40 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:26 DR:40 LR:-174.9 LO:174.9);ALT=]chr17:34188507]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr15	59943023	+	chr15	59949602	+	.	56	0	5963454_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5963454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:59943023(+)-15:59949602(-)__15_59927001_59952001D;SPAN=6579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:61 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:56 LR:-178.2 LO:178.2);ALT=A[chr15:59949602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59944527	+	chr15	59949604	+	.	74	7	5963460_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5963460_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59927001_59952001_89C;SPAN=5077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:66 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:7 DR:74 LR:-224.5 LO:224.5);ALT=T[chr15:59949604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	62706095	+	chr15	62707793	+	.	73	50	5967651_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATT;MAPQ=60;MATEID=5967651_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_62695501_62720501_151C;SPAN=1698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:19 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:50 DR:73 LR:-303.7 LO:303.7);ALT=T[chr15:62707793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63447972	+	chr15	63449595	+	.	75	0	5969026_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=5969026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:63447972(+)-15:63449595(-)__15_63430501_63455501D;SPAN=1623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:70 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:0 DR:75 LR:-221.2 LO:221.2);ALT=G[chr15:63449595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64381051	+	chr15	64385852	+	ATAAACC	34	44	5970707_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=ATAAACC;MAPQ=60;MATEID=5970707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64361501_64386501_199C;SPAN=4801;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:63 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:44 DR:34 LR:-214.6 LO:214.6);ALT=C[chr15:64385852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64452451	+	chr15	64455048	+	.	112	0	5970813_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5970813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64452451(+)-15:64455048(-)__15_64435001_64460001D;SPAN=2597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:84 GQ:30 PL:[330.0, 30.0, 0.0] SR:0 DR:112 LR:-330.1 LO:330.1);ALT=A[chr15:64455048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64669154	+	chr15	64673556	+	.	86	0	5971195_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5971195_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64669154(+)-15:64673556(-)__15_64655501_64680501D;SPAN=4402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:55 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:0 DR:86 LR:-254.2 LO:254.2);ALT=C[chr15:64673556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66161963	+	chr15	66169668	+	.	82	13	5974226_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5974226_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_66150001_66175001_191C;SPAN=7705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:68 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:13 DR:82 LR:-260.8 LO:260.8);ALT=G[chr15:66169668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	68426020	+	chr15	68428928	+	.	56	40	5978453_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGAAATTTAGATTTTTA;MAPQ=60;MATEID=5978453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_68404001_68429001_49C;SPAN=2908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:33 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:40 DR:56 LR:-237.7 LO:237.7);ALT=A[chr15:68428928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69080263	+	chr15	69113048	+	.	52	0	5979461_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5979461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:69080263(+)-15:69113048(-)__15_69090001_69115001D;SPAN=32785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:37 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=A[chr15:69113048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69745360	+	chr15	69747508	+	.	39	9	5980559_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=54;MATEID=5980559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_69727001_69752001_96C;SPAN=2148;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:44 DP:911 GQ:99 PL:[0.0, 101.1, 2413.0] SR:9 DR:39 LR:101.6 LO:70.92);ALT=G[chr15:69747508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	70596153	+	chr15	70594649	+	.	39	0	5981768_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5981768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:70594649(-)-15:70596153(+)__15_70584501_70609501D;SPAN=1504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:69 GQ:57.2 PL:[110.0, 0.0, 57.2] SR:0 DR:39 LR:-110.9 LO:110.9);ALT=]chr15:70596153]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	71708609	+	chr15	71713691	+	ACC	69	42	5983513_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=ACC;MAPQ=60;MATEID=5983513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_71711501_71736501_121C;SPAN=5082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:14 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:42 DR:69 LR:-267.4 LO:267.4);ALT=A[chr15:71713691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72385978	+	chr15	72388159	+	.	43	32	5984719_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCCTGTAATCCCA;MAPQ=60;MATEID=5984719_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72373001_72398001_104C;SPAN=2181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:25 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:32 DR:43 LR:-191.4 LO:191.4);ALT=A[chr15:72388159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72509880	+	chr15	72523470	+	.	49	0	5984950_1	99.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5984950_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:72509880(+)-15:72523470(-)__15_72520001_72545001D;SPAN=13590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:60 GQ:0.2 PL:[145.4, 0.0, 0.2] SR:0 DR:49 LR:-154.5 LO:154.5);ALT=T[chr15:72523470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72511453	+	chr15	72523456	+	.	163	30	5984951_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5984951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72520001_72545001_92C;SPAN=12003;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:180 DP:27 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:30 DR:163 LR:-534.7 LO:534.7);ALT=T[chr15:72523456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74751238	+	chr15	74753377	+	.	36	5	5988963_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5988963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_74749501_74774501_206C;SPAN=2139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:64 GQ:48.8 PL:[104.9, 0.0, 48.8] SR:5 DR:36 LR:-105.8 LO:105.8);ALT=C[chr15:74753377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75147037	+	chr15	75165604	+	.	31	0	5989635_1	87.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5989635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75147037(+)-15:75165604(-)__15_75141501_75166501D;SPAN=18567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:56 GQ:47.6 PL:[87.2, 0.0, 47.6] SR:0 DR:31 LR:-87.74 LO:87.74);ALT=G[chr15:75165604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75221619	+	chr15	75230314	+	.	131	0	5990015_1	99.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5990015_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75221619(+)-15:75230314(-)__15_75215001_75240001D;SPAN=8695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:131 DP:119 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:0 DR:131 LR:-386.2 LO:386.2);ALT=T[chr15:75230314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76585042	+	chr15	76603688	+	.	46	2	5992866_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=5992866_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76587001_76612001_276C;SPAN=18646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:44 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:2 DR:46 LR:-138.6 LO:138.6);ALT=C[chr15:76603688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76588079	+	chr15	76603690	+	.	32	7	5992872_1	92.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=5992872_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_15_76587001_76612001_30C;SPAN=15611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:73 GQ:82.7 PL:[92.6, 0.0, 82.7] SR:7 DR:32 LR:-92.47 LO:92.47);ALT=C[chr15:76603690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78585673	+	chr15	78591902	+	.	43	0	5996096_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5996096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78585673(+)-15:78591902(-)__15_78571501_78596501D;SPAN=6229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:70 GQ:47 PL:[122.9, 0.0, 47.0] SR:0 DR:43 LR:-124.8 LO:124.8);ALT=G[chr15:78591902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78832908	+	chr15	78834820	+	.	118	0	5996829_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5996829_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78832908(+)-15:78834820(-)__15_78816501_78841501D;SPAN=1912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:85 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:0 DR:118 LR:-349.9 LO:349.9);ALT=C[chr15:78834820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83551631	+	chr15	83557671	+	.	72	41	6005337_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCAGCCACT;MAPQ=60;MATEID=6005337_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_15_83545001_83570001_155C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:33 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:41 DR:72 LR:-267.4 LO:267.4);ALT=T[chr15:83557671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85231035	+	chr15	85259255	+	.	77	0	6008921_1	99.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6008921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:85231035(+)-15:85259255(-)__15_85235501_85260501D;SPAN=28220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:54 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:0 DR:77 LR:-227.8 LO:227.8);ALT=A[chr15:85259255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85234879	+	chr15	85259256	+	.	92	30	6008899_1	99.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=CTGC;MAPQ=60;MATEID=6008899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_85211001_85236001_210C;SPAN=24377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:64 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:30 DR:92 LR:-287.2 LO:287.2);ALT=C[chr15:85259256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90774928	+	chr15	90777080	+	.	71	0	6029401_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6029401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:90774928(+)-15:90777080(-)__15_90772501_90797501D;SPAN=2152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:117 GQ:80.6 PL:[202.7, 0.0, 80.6] SR:0 DR:71 LR:-205.5 LO:205.5);ALT=G[chr15:90777080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90775618	+	chr15	90777093	+	.	101	0	6029407_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6029407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:90775618(+)-15:90777093(-)__15_90772501_90797501D;SPAN=1475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:101 DP:143 GQ:50.6 PL:[294.8, 0.0, 50.6] SR:0 DR:101 LR:-304.3 LO:304.3);ALT=T[chr15:90777093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90931628	+	chr15	90934006	+	.	47	32	6030140_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6030140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90919501_90944501_281C;SPAN=2378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:115 GQ:94.4 PL:[183.5, 0.0, 94.4] SR:32 DR:47 LR:-184.9 LO:184.9);ALT=T[chr15:90934006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91981580	+	chr15	91989266	+	.	49	34	6034063_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=6034063_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91973001_91998001_93C;SPAN=7686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:94 GQ:27.5 PL:[199.1, 0.0, 27.5] SR:34 DR:49 LR:-206.3 LO:206.3);ALT=A[chr15:91989266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91989617	+	chr15	91983461	+	A	35	27	6034067_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=6034067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91973001_91998001_397C;SPAN=6156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:27 DR:35 LR:-163.7 LO:163.7);ALT=]chr15:91989617]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	92674576	+	chr15	92677071	+	.	109	87	6036556_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6036556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_92659001_92684001_237C;SPAN=2495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:44 GQ:46 PL:[505.0, 46.0, 0.0] SR:87 DR:109 LR:-505.0 LO:505.0);ALT=T[chr15:92677071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	100416715	+	chr15	100423235	+	.	40	0	6062961_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6062961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100416715(+)-15:100423235(-)__15_100401001_100426001D;SPAN=6520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:63 GQ:35.9 PL:[115.1, 0.0, 35.9] SR:0 DR:40 LR:-117.1 LO:117.1);ALT=T[chr15:100423235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	104060	+	chr16	105457	+	.	31	31	6071216_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6071216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_98001_123001_130C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:115 GQ:99 PL:[120.8, 0.0, 157.1] SR:31 DR:31 LR:-120.7 LO:121.0);ALT=T[chr16:105457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	128332	+	chr16	129421	+	.	135	13	6071097_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6071097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_122501_147501_174C;SPAN=1089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:69 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:13 DR:135 LR:-409.3 LO:409.3);ALT=G[chr16:129421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1359775	+	chr16	1364019	+	.	45	27	6075526_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6075526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1347501_1372501_55C;SPAN=4244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:59 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:27 DR:45 LR:-174.9 LO:174.9);ALT=G[chr16:1364019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1359780	+	chr16	1364293	+	.	47	0	6075527_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6075527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1359780(+)-16:1364293(-)__16_1347501_1372501D;SPAN=4513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:61 GQ:6.8 PL:[138.8, 0.0, 6.8] SR:0 DR:47 LR:-145.3 LO:145.3);ALT=C[chr16:1364293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1402047	+	chr16	1411742	+	.	40	0	6075659_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6075659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1402047(+)-16:1411742(-)__16_1396501_1421501D;SPAN=9695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:73 GQ:62.9 PL:[112.4, 0.0, 62.9] SR:0 DR:40 LR:-112.9 LO:112.9);ALT=G[chr16:1411742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1422869	+	chr16	1424141	+	.	35	0	6075579_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6075579_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1422869(+)-16:1424141(-)__16_1421001_1446001D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:58 GQ:40.4 PL:[99.8, 0.0, 40.4] SR:0 DR:35 LR:-101.2 LO:101.2);ALT=T[chr16:1424141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1828661	+	chr16	1832500	+	.	53	0	6076854_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6076854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1828661(+)-16:1832500(-)__16_1813001_1838001D;SPAN=3839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:75 GQ:26 PL:[154.7, 0.0, 26.0] SR:0 DR:53 LR:-159.7 LO:159.7);ALT=C[chr16:1832500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1833085	+	chr16	1836560	+	.	40	0	6076861_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6076861_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1833085(+)-16:1836560(-)__16_1813001_1838001D;SPAN=3475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:0 DR:40 LR:-109.9 LO:109.9);ALT=G[chr16:1836560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2009755	+	chr16	2011152	+	.	74	122	6077699_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6077699_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2009001_2034001_286C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:168 DP:155 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:122 DR:74 LR:-498.4 LO:498.4);ALT=G[chr16:2011152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2564183	+	chr16	2569218	+	.	84	185	6080032_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6080032_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2548001_2573001_120C;SPAN=5035;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:233 DP:187 GQ:62.8 PL:[689.8, 62.8, 0.0] SR:185 DR:84 LR:-689.9 LO:689.9);ALT=G[chr16:2569218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2802856	+	chr16	2806334	+	.	51	21	6080818_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6080818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2793001_2818001_240C;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:127 GQ:99 PL:[153.8, 0.0, 153.8] SR:21 DR:51 LR:-153.8 LO:153.8);ALT=G[chr16:2806334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4391643	+	chr16	4401230	+	.	48	0	6086527_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6086527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4391643(+)-16:4401230(-)__16_4385501_4410501D;SPAN=9587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:79 GQ:54.5 PL:[137.0, 0.0, 54.5] SR:0 DR:48 LR:-139.0 LO:139.0);ALT=C[chr16:4401230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18800442	+	chr16	18801566	+	.	38	19	6138794_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=54;MATEID=6138794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_144C;SPAN=1124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:146 GQ:99 PL:[112.4, 0.0, 241.1] SR:19 DR:38 LR:-112.3 LO:114.9);ALT=T[chr16:18801566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18809410	+	chr16	18812805	+	.	33	0	6138826_1	73.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6138826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:18809410(+)-16:18812805(-)__16_18791501_18816501D;SPAN=3395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:132 GQ:73.4 PL:[73.4, 0.0, 245.0] SR:0 DR:33 LR:-73.17 LO:78.46);ALT=T[chr16:18812805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18810157	+	chr16	18812752	+	.	79	25	6138829_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6138829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_205C;SPAN=2595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:112 GQ:16.8 PL:[303.6, 16.8, 0.0] SR:25 DR:79 LR:-308.5 LO:308.5);ALT=C[chr16:18812752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21170099	+	chr16	21172295	+	.	38	0	6147051_1	98.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6147051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:21170099(+)-16:21172295(-)__16_21168001_21193001D;SPAN=2196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:101 GQ:98.3 PL:[98.3, 0.0, 144.5] SR:0 DR:38 LR:-98.08 LO:98.61);ALT=G[chr16:21172295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21594442	+	chr16	22710751	-	ATG	48	34	6154760_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=ATG;MAPQ=60;MATEID=6154760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_22687001_22712001_390C;SPAN=1116309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:50 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:34 DR:48 LR:-204.7 LO:204.7);ALT=C]chr16:22710751];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	21964777	+	chr16	21968555	+	.	63	15	6150819_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6150819_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21952001_21977001_384C;SPAN=3778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:98 GQ:9.8 PL:[227.6, 0.0, 9.8] SR:15 DR:63 LR:-239.6 LO:239.6);ALT=G[chr16:21968555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23047775	+	chr16	23049532	+	GATTCT	50	32	6155842_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GATTCT;MAPQ=60;MATEID=6155842_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23030001_23055001_306C;SPAN=1757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:74 GQ:16.5 PL:[211.2, 16.5, 0.0] SR:32 DR:50 LR:-211.3 LO:211.3);ALT=A[chr16:23049532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23598642	+	chr16	23607442	+	.	69	90	6157996_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6157996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23593501_23618501_192C;SPAN=8800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:134 GQ:19.5 PL:[363.0, 19.5, 0.0] SR:90 DR:69 LR:-369.8 LO:369.8);ALT=T[chr16:23607442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30075855	+	chr16	30078767	+	.	40	0	6182052_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6182052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30075855(+)-16:30078767(-)__16_30061501_30086501D;SPAN=2912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:103 GQ:99 PL:[104.3, 0.0, 143.9] SR:0 DR:40 LR:-104.1 LO:104.5);ALT=A[chr16:30078767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30075855	+	chr16	30078550	+	.	100	0	6182051_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6182051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30075855(+)-16:30078550(-)__16_30061501_30086501D;SPAN=2695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:158 GQ:95.9 PL:[287.3, 0.0, 95.9] SR:0 DR:100 LR:-292.5 LO:292.5);ALT=A[chr16:30078550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30077166	+	chr16	30078769	+	.	44	0	6182055_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6182055_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30077166(+)-16:30078769(-)__16_30061501_30086501D;SPAN=1603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:252 GQ:77.2 PL:[77.2, 0.0, 532.7] SR:0 DR:44 LR:-76.97 LO:96.82);ALT=C[chr16:30078769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30077249	+	chr16	30078551	+	.	100	74	6182056_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAGG;MAPQ=60;MATEID=6182056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30061501_30086501_297C;SPAN=1302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:211 GQ:99 PL:[405.2, 0.0, 104.8] SR:74 DR:100 LR:-414.6 LO:414.6);ALT=G[chr16:30078551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30195046	+	chr16	30197917	+	AATGAGCCGGCAGGTGGTCCGCTCCAGCAAGTTCCGCCACGTGTTTGGACAGCCGGCCAAGGCCGACCAGTGCTATGAAGATGTGCGCGTCTCACAGACCACCTGGGACAGTGGCTTCTGTGCTGTCAACCCTAAGTTTGTGGCCCTGATCTGTGAGGCCAGCGGGGGAGGGGCCTTCCTGGTGCTGCCCCTGGGCA	41	109	6182552_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AATGAGCCGGCAGGTGGTCCGCTCCAGCAAGTTCCGCCACGTGTTTGGACAGCCGGCCAAGGCCGACCAGTGCTATGAAGATGTGCGCGTCTCACAGACCACCTGGGACAGTGGCTTCTGTGCTGTCAACCCTAAGTTTGTGGCCCTGATCTGTGAGGCCAGCGGGGGAGGGGCCTTCCTGGTGCTGCCCCTGGGCA;MAPQ=60;MATEID=6182552_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_30184001_30209001_269C;SPAN=2871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:110 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:109 DR:41 LR:-369.7 LO:369.7);ALT=G[chr16:30197917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30195046	+	chr16	30196527	+	.	163	22	6182551_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=6182551_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GACGAC;SCTG=c_16_30184001_30209001_269C;SPAN=1481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:171 DP:137 GQ:45.8 PL:[397.9, 45.8, 0.0] SR:22 DR:163 LR:-397.9 LO:397.9);ALT=G[chr16:30196527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30435905	+	chr16	30441102	+	.	31	0	6183824_1	75.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6183824_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30435905(+)-16:30441102(-)__16_30429001_30454001D;SPAN=5197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:100 GQ:75.2 PL:[75.2, 0.0, 167.6] SR:0 DR:31 LR:-75.24 LO:77.17);ALT=G[chr16:30441102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31102666	+	chr16	31105876	+	.	32	20	6186471_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=6186471_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_31090501_31115501_120C;SPAN=3210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:119 GQ:99 PL:[103.1, 0.0, 185.6] SR:20 DR:32 LR:-103.1 LO:104.4);ALT=G[chr16:31105876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31104787	+	chr16	31105872	+	.	51	0	6186478_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6186478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:31104787(+)-16:31105872(-)__16_31090501_31115501D;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:105 GQ:99 PL:[140.0, 0.0, 113.6] SR:0 DR:51 LR:-140.0 LO:140.0);ALT=A[chr16:31105872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31191548	+	chr16	31193832	+	ATTATACCCAACAAGCAACCCAA	86	25	6186845_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ATTATACCCAACAAGCAACCCAA;MAPQ=60;MATEID=6186845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_31188501_31213501_357C;SPAN=2284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:121 GQ:13.7 PL:[277.7, 0.0, 13.7] SR:25 DR:86 LR:-291.4 LO:291.4);ALT=G[chr16:31193832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	32600335	+	chr16	32601844	+	.	40	17	6192885_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGGCCTATGGTGACAAACTGAATATCCCCAGATAA;MAPQ=60;MATEID=6192885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_32585001_32610001_34C;SPAN=1509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:83 GQ:43.7 PL:[155.9, 0.0, 43.7] SR:17 DR:40 LR:-159.1 LO:159.1);ALT=A[chr16:32601844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	33238416	+	chr16	33237191	+	.	32	0	6197586_1	34.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=6197586_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:33237191(-)-16:33238416(+)__16_33222001_33247001D;SPAN=1225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:263 GQ:34.6 PL:[34.6, 0.0, 602.3] SR:0 DR:32 LR:-34.38 LO:64.95);ALT=]chr16:33238416]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	33374049	+	chr16	33379406	+	TTTAGGT	46	28	6198019_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;INSERTION=TTTAGGT;MAPQ=60;MATEID=6198019_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_16_33369001_33394001_144C;SPAN=5357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:149 GQ:99 PL:[184.1, 0.0, 177.5] SR:28 DR:46 LR:-184.1 LO:184.1);ALT=C[chr16:33379406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57725395	+	chr16	57727847	+	.	83	50	6221380_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6221380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57722001_57747001_146C;SPAN=2452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:22 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:50 DR:83 LR:-340.0 LO:340.0);ALT=G[chr16:57727847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58624545	+	chr16	58663331	+	CCAG	69	33	6223031_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=CCAG;MAPQ=60;MATEID=6223031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_58653001_58678001_43C;SPAN=38786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:11 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:33 DR:69 LR:-254.2 LO:254.2);ALT=T[chr16:58663331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66586696	+	chr16	66596974	+	.	32	3	6234080_1	92.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6234080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66566501_66591501_200C;SPAN=10278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:59 GQ:50 PL:[92.9, 0.0, 50.0] SR:3 DR:32 LR:-93.63 LO:93.63);ALT=G[chr16:66596974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66586697	+	chr16	66592092	+	.	55	61	6234081_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6234081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66566501_66591501_80C;SPAN=5395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:56 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:61 DR:55 LR:-283.9 LO:283.9);ALT=G[chr16:66592092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67261164	+	chr16	67262255	+	.	54	0	6235464_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6235464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67261164(+)-16:67262255(-)__16_67252501_67277501D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:58 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:54 LR:-171.6 LO:171.6);ALT=A[chr16:67262255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69761829	-	chr16	69762896	+	.	41	41	6241149_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TCAAG;MAPQ=60;MATEID=6241149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69751501_69776501_123C;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:56 GQ:18 PL:[198.0, 18.0, 0.0] SR:41 DR:41 LR:-198.0 LO:198.0);ALT=[chr16:69762896[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	74330817	+	chr16	74334009	+	.	31	0	6249585_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6249585_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:74330817(+)-16:74334009(-)__16_74333001_74358001D;SPAN=3192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=C[chr16:74334009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75600418	+	chr16	75601934	+	AACACAGATGCGTGGAGTCCGCGAAGATTCGAGCGAAATATCCCGACAGGGTTCC	71	99	6252445_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GGTGA;INSERTION=AACACAGATGCGTGGAGTCCGCGAAGATTCGAGCGAAATATCCCGACAGGGTTCC;MAPQ=60;MATEID=6252445_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_75582501_75607501_157C;SPAN=1516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:62 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:99 DR:71 LR:-409.3 LO:409.3);ALT=G[chr16:75601934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	83841728	+	chr16	83842910	+	GCAGACACTCCTGCAGCAGATGCAAGATAAATTTCAGACCATGTCTGACCAGATCATTGGGAGAA	73	137	6265376_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=GCAGACACTCCTGCAGCAGATGCAAGATAAATTTCAGACCATGTCTGACCAGATCATTGGGAGAA;MAPQ=60;MATEID=6265376_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_83839001_83864001_27C;SPAN=1182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:192 DP:83 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:137 DR:73 LR:-567.7 LO:567.7);ALT=T[chr16:83842910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	84623920	+	chr16	84651442	+	.	37	0	6266910_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6266910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:84623920(+)-16:84651442(-)__16_84647501_84672501D;SPAN=27522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:70 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.6 LO:103.6);ALT=G[chr16:84651442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85302493	+	chr16	85304391	+	.	52	33	6267974_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6267974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85284501_85309501_134C;SPAN=1898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:17 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:33 DR:52 LR:-224.5 LO:224.5);ALT=G[chr16:85304391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85833358	+	chr16	85834808	+	.	37	29	6269443_1	75.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6269443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85823501_85848501_176C;SPAN=1450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:333 GQ:75 PL:[75.0, 0.0, 731.9] SR:29 DR:37 LR:-74.83 LO:106.4);ALT=G[chr16:85834808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85833409	+	chr16	85838538	+	.	186	0	6269447_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6269447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85833409(+)-16:85838538(-)__16_85823501_85848501D;SPAN=5129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:186 DP:114 GQ:50.2 PL:[551.2, 50.2, 0.0] SR:0 DR:186 LR:-551.2 LO:551.2);ALT=G[chr16:85838538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85932830	+	chr16	85936619	+	.	31	3	6269352_1	88.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6269352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85921501_85946501_15C;SPAN=3789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:63 GQ:62.3 PL:[88.7, 0.0, 62.3] SR:3 DR:31 LR:-88.77 LO:88.77);ALT=G[chr16:85936619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	86622031	+	chr16	86621014	+	.	50	0	6270611_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6270611_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:86621014(-)-16:86622031(+)__16_86607501_86632501D;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:72 GQ:26.9 PL:[145.7, 0.0, 26.9] SR:0 DR:50 LR:-149.9 LO:149.9);ALT=]chr16:86622031]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	87773402	+	chr16	87771949	+	.	59	0	6272747_1	99.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=6272747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:87771949(-)-16:87773402(+)__16_87759001_87784001D;SPAN=1453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:67 GQ:14.7 PL:[191.4, 14.7, 0.0] SR:0 DR:59 LR:-192.0 LO:192.0);ALT=]chr16:87773402]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	88876967	+	chr16	88878227	+	CGATGTAGTCGATGCGGCCCCCGTGGGTCGCCTTCAGGTGTCGCGCCAGGAGGCCGATGGCGGCGCGGAAGGAGGCGGGGTCCTTCAGGACGGGCGAGATGTC	120	166	6275057_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=CGATGTAGTCGATGCGGCCCCCGTGGGTCGCCTTCAGGTGTCGCGCCAGGAGGCCGATGGCGGCGCGGAAGGAGGCGGGGTCCTTCAGGACGGGCGAGATGTC;MAPQ=60;MATEID=6275057_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_88861501_88886501_194C;SPAN=1260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:222 DP:91 GQ:59.8 PL:[656.8, 59.8, 0.0] SR:166 DR:120 LR:-656.9 LO:656.9);ALT=G[chr16:88878227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88923634	+	chr16	88925024	+	.	40	0	6274707_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6274707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88923634(+)-16:88925024(-)__16_88910501_88935501D;SPAN=1390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:40 LR:-118.8 LO:118.8);ALT=C[chr16:88925024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88923634	+	chr16	88926070	+	.	34	0	6274708_1	96.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6274708_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88923634(+)-16:88926070(-)__16_88910501_88935501D;SPAN=2436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:59 GQ:46.7 PL:[96.2, 0.0, 46.7] SR:0 DR:34 LR:-97.17 LO:97.17);ALT=C[chr16:88926070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89967871	+	chr16	89969134	+	.	55	19	6277041_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAGGGGCTGTGAGGGGTGAGGGTGAAATCCCTCCTTAAGACGGGCCTCC;MAPQ=60;MATEID=6277041_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_16_89964001_89989001_53C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:13 GQ:18 PL:[198.0, 18.0, 0.0] SR:19 DR:55 LR:-198.0 LO:198.0);ALT=C[chr16:89969134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	20626	+	chr17	21729	+	.	56	0	6277629_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6277629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:20626(+)-17:21729(-)__17_1_25001D;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:42 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:56 LR:-165.0 LO:165.0);ALT=G[chr17:21729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	862402	-	chr19	5680466	+	.	35	0	6708496_1	97.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6708496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:862402(-)-19:5680466(-)__19_5659501_5684501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:67 GQ:64.4 PL:[97.4, 0.0, 64.4] SR:0 DR:35 LR:-97.72 LO:97.72);ALT=[chr19:5680466[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr17	1268383	+	chr17	1303387	+	.	97	0	6282326_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6282326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1268383(+)-17:1303387(-)__17_1298501_1323501D;SPAN=35004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:45 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:0 DR:97 LR:-287.2 LO:287.2);ALT=C[chr17:1303387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	2719930	+	chr17	2721218	+	.	58	42	6287557_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6287557_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_2719501_2744501_109C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:42 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:42 DR:58 LR:-237.7 LO:237.7);ALT=T[chr17:2721218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3568093	+	chr17	3571782	+	.	34	4	6289413_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6289413_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CC;SCTG=c_17_3552501_3577501_138C;SPAN=3689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:61 GQ:46.4 PL:[99.2, 0.0, 46.4] SR:4 DR:34 LR:-99.92 LO:99.92);ALT=C[chr17:3571782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3620138	+	chr17	3627014	+	.	41	0	6290312_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6290312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:3620138(+)-17:3627014(-)__17_3626001_3651001D;SPAN=6876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:49 GQ:3.3 PL:[125.4, 3.3, 0.0] SR:0 DR:41 LR:-130.5 LO:130.5);ALT=A[chr17:3627014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3623698	+	chr17	3626982	+	.	58	24	6290314_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6290314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_3626001_3651001_6C;SPAN=3284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:41 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:24 DR:58 LR:-194.7 LO:194.7);ALT=T[chr17:3626982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4337462	+	chr17	4342948	+	.	52	102	6292535_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGCAGG;MAPQ=60;MATEID=6292535_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_4336501_4361501_356C;SPAN=5486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:119 DP:140 GQ:14.7 PL:[369.6, 14.7, 0.0] SR:102 DR:52 LR:-381.1 LO:381.1);ALT=G[chr17:4342948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4614078	+	chr17	4619704	+	.	54	0	6293607_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6293607_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:4614078(+)-17:4619704(-)__17_4606001_4631001D;SPAN=5626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:96 GQ:79.7 PL:[152.3, 0.0, 79.7] SR:0 DR:54 LR:-153.4 LO:153.4);ALT=G[chr17:4619704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4863843	+	chr17	4871015	+	CTTTTACGAAACTCCACTTTCTGTTGTTTCTCTTGCTCTTGTAGTTTCTTCAGGCGGGCGGCCTGTT	49	23	6294571_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTTTTACGAAACTCCACTTTCTGTTGTTTCTCTTGCTCTTGTAGTTTCTTCAGGCGGGCGGCCTGTT;MAPQ=60;MATEID=6294571_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_4851001_4876001_106C;SPAN=7172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:103 GQ:68 PL:[180.2, 0.0, 68.0] SR:23 DR:49 LR:-182.7 LO:182.7);ALT=C[chr17:4871015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5323605	+	chr17	5324612	+	.	43	0	6296485_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6296485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5323605(+)-17:5324612(-)__17_5316501_5341501D;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:81 GQ:74 PL:[120.2, 0.0, 74.0] SR:0 DR:43 LR:-120.5 LO:120.5);ALT=C[chr17:5324612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7144278	+	chr17	7145471	+	.	49	0	6301878_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6301878_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7144278(+)-17:7145471(-)__17_7129501_7154501D;SPAN=1193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:98 GQ:99 PL:[135.2, 0.0, 102.2] SR:0 DR:49 LR:-135.4 LO:135.4);ALT=A[chr17:7145471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7211075	+	chr17	7212929	+	.	111	0	6302549_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6302549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7211075(+)-17:7212929(-)__17_7203001_7228001D;SPAN=1854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:107 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:111 LR:-326.8 LO:326.8);ALT=A[chr17:7212929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7211432	+	chr17	7212932	+	.	51	7	6302550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6302550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_7203001_7228001_234C;SPAN=1500;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:108 GQ:99 PL:[149.0, 0.0, 112.7] SR:7 DR:51 LR:-149.3 LO:149.3);ALT=G[chr17:7212932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7336437	+	chr17	7337683	+	.	44	0	6302286_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6302286_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7336437(+)-17:7337683(-)__17_7325501_7350501D;SPAN=1246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:30 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:0 DR:44 LR:-128.7 LO:128.7);ALT=C[chr17:7337683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8065086	+	chr17	8066194	+	CATCCACCTGGGCCTGGGTCTGCTGCAGTCTCCTGTTACTGGTGAGGTTTGGAGGGGGTGCAGGGGGACCACCCTCCCCAGCCGGGGCAGCAGGGGGGGCCGTGGCAGCGGTAGCAG	81	92	6305596_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=CATCCACCTGGGCCTGGGTCTGCTGCAGTCTCCTGTTACTGGTGAGGTTTGGAGGGGGTGCAGGGGGACCACCCTCCCCAGCCGGGGCAGCAGGGGGGGCCGTGGCAGCGGTAGCAG;MAPQ=60;MATEID=6305596_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_8060501_8085501_71C;SPAN=1108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:107 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:92 DR:81 LR:-389.5 LO:389.5);ALT=T[chr17:8066194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8246645	+	chr17	8247969	+	.	63	11	6306144_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GCTAATTTTTGTATTTTTAGTAGAGACGGGGTTT;MAPQ=60;MATEID=6306144_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_17_8232001_8257001_352C;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:37 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:11 DR:63 LR:-208.0 LO:208.0);ALT=T[chr17:8247969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	9460847	+	chr17	9471688	+	.	31	24	6309664_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6309664_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_9457001_9482001_247C;SPAN=10841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:90 GQ:99 PL:[110.9, 0.0, 107.6] SR:24 DR:31 LR:-111.0 LO:111.0);ALT=T[chr17:9471688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25536553	+	chr17	25540382	+	.	38	22	6349875_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAATTCACATGGCA;MAPQ=60;MATEID=6349875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25529001_25554001_137C;SPAN=3829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:92 GQ:71 PL:[150.2, 0.0, 71.0] SR:22 DR:38 LR:-151.5 LO:151.5);ALT=A[chr17:25540382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25958358	+	chr17	25967595	+	.	89	0	6351234_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6351234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:25958358(+)-17:25967595(-)__17_25945501_25970501D;SPAN=9237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:75 GQ:24 PL:[264.0, 24.0, 0.0] SR:0 DR:89 LR:-264.1 LO:264.1);ALT=C[chr17:25967595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27216047	+	chr17	27224543	+	.	32	19	6355115_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6355115_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_27195001_27220001_204C;SPAN=8496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:19 DR:32 LR:-112.2 LO:112.2);ALT=G[chr17:27224543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29632650	+	chr17	29640997	+	.	94	5	6363310_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6363310_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_29620501_29645501_208C;SPAN=8347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:93 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:5 DR:94 LR:-277.3 LO:277.3);ALT=T[chr17:29640997[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30677349	+	chr17	30678804	+	.	33	44	6366796_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTAT;MAPQ=60;MATEID=6366796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30674001_30699001_163C;SECONDARY;SPAN=1455;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:92 GQ:11.6 PL:[209.6, 0.0, 11.6] SR:44 DR:33 LR:-219.6 LO:219.6);ALT=T[chr17:30678804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34136609	+	chr17	34147025	+	.	71	0	6376454_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6376454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34136609(+)-17:34147025(-)__17_34128501_34153501D;SPAN=10416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:89 GQ:5.6 PL:[210.2, 0.0, 5.6] SR:0 DR:71 LR:-222.0 LO:222.0);ALT=A[chr17:34147025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34205643	+	chr17	34207234	+	.	48	22	6376754_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6376754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_34202001_34227001_212C;SPAN=1591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:106 GQ:93.5 PL:[162.8, 0.0, 93.5] SR:22 DR:48 LR:-163.7 LO:163.7);ALT=T[chr17:34207234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34416157	+	chr17	34417331	+	.	49	0	6377628_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6377628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34416157(+)-17:34417331(-)__17_34398001_34423001D;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:94 GQ:90.2 PL:[136.4, 0.0, 90.2] SR:0 DR:49 LR:-136.7 LO:136.7);ALT=A[chr17:34417331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40149261	+	chr17	40169357	+	GGCTTTTGTATAATAATTATAAGCTTCATTGTAATCTTTCTTGGCATAGTATGCATTTCCTTGTTCCTTGAAAGTCTCTGCTTC	33	39	6397494_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GGCTTTTGTATAATAATTATAAGCTTCATTGTAATCTTTCTTGGCATAGTATGCATTTCCTTGTTCCTTGAAAGTCTCTGCTTC;MAPQ=60;MATEID=6397494_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_17_40155501_40180501_306C;SPAN=20096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:39 DR:33 LR:-155.1 LO:155.1);ALT=T[chr17:40169357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40282608	+	chr17	40306911	+	.	115	8	6397962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6397962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40302501_40327501_150C;SPAN=24303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:40 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:8 DR:115 LR:-340.0 LO:340.0);ALT=A[chr17:40306911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41150578	+	chr17	41151947	+	.	51	0	6401112_1	99.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6401112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41150578(+)-17:41151947(-)__17_41135501_41160501D;SPAN=1369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:121 GQ:99 PL:[135.8, 0.0, 155.6] SR:0 DR:51 LR:-135.6 LO:135.7);ALT=C[chr17:41151947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42422703	+	chr17	42426522	+	.	48	2	6405863_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GCAGG;MAPQ=60;MATEID=6405863_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42409501_42434501_444C;SPAN=3819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:207 GQ:99 PL:[214.7, 0.0, 287.3] SR:2 DR:48 LR:-214.6 LO:215.2);ALT=G[chr17:42426522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42422754	+	chr17	42426787	+	.	52	0	6405866_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6405866_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:42422754(+)-17:42426787(-)__17_42409501_42434501D;SPAN=4033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:98 GQ:92.3 PL:[145.1, 0.0, 92.3] SR:0 DR:52 LR:-145.7 LO:145.7);ALT=C[chr17:42426787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46654382	+	chr17	46667487	+	.	38	10	6419627_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=6419627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46648001_46673001_284C;SPAN=13105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:86 GQ:98.9 PL:[108.8, 0.0, 98.9] SR:10 DR:38 LR:-108.8 LO:108.8);ALT=A[chr17:46667487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46667953	+	chr17	46677808	+	.	45	58	6419669_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6419669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46648001_46673001_154C;SPAN=9855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:46 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:58 DR:45 LR:-241.0 LO:241.0);ALT=T[chr17:46677808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46908490	+	chr17	46925425	+	.	31	0	6420392_1	88.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6420392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46908490(+)-17:46925425(-)__17_46917501_46942501D;SPAN=16935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:50 GQ:32.6 PL:[88.7, 0.0, 32.6] SR:0 DR:31 LR:-90.21 LO:90.21);ALT=T[chr17:46925425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46908493	+	chr17	46919058	+	.	54	0	6420394_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6420394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46908493(+)-17:46919058(-)__17_46917501_46942501D;SPAN=10565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:51 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=A[chr17:46919058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49231056	+	chr17	49233010	+	.	63	0	6428431_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6428431_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49231056(+)-17:49233010(-)__17_49220501_49245501D;SPAN=1954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:92 GQ:38 PL:[183.2, 0.0, 38.0] SR:0 DR:63 LR:-188.2 LO:188.2);ALT=G[chr17:49233010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49231067	+	chr17	49237338	+	.	60	0	6428433_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6428433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49231067(+)-17:49237338(-)__17_49220501_49245501D;SPAN=6271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:109 GQ:95.9 PL:[168.5, 0.0, 95.9] SR:0 DR:60 LR:-169.6 LO:169.6);ALT=A[chr17:49237338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55089757	+	chr17	55092846	+	.	54	0	6442414_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6442414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55089757(+)-17:55092846(-)__17_55076001_55101001D;SPAN=3089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:5 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=T[chr17:55092846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55687811	+	chr17	55689915	+	.	70	45	6444031_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6444031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_55688501_55713501_320C;SPAN=2104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:33 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:45 DR:70 LR:-254.2 LO:254.2);ALT=T[chr17:55689915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66508689	+	chr17	66511532	+	.	56	12	6478114_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6478114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_66493001_66518001_366C;SPAN=2843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:106 GQ:86.9 PL:[169.4, 0.0, 86.9] SR:12 DR:56 LR:-170.7 LO:170.7);ALT=G[chr17:66511532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72462909	+	chr17	72469670	+	.	35	0	6494684_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6494684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:72462909(+)-17:72469670(-)__17_72446501_72471501D;SPAN=6761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:0 DR:35 LR:-91.97 LO:92.16);ALT=C[chr17:72469670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73038393	+	chr17	73043018	+	.	43	0	6496664_1	99.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6496664_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73038393(+)-17:73043018(-)__17_73034501_73059501D;SPAN=4625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:105 GQ:99 PL:[113.6, 0.0, 140.0] SR:0 DR:43 LR:-113.5 LO:113.7);ALT=A[chr17:73043018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	114953559	+	chr17	73178992	+	.	40	0	7503369_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=7503369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73178992(-)-23:114953559(+)__23_114929501_114954501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:40 LR:-125.4 LO:125.4);ALT=]chrX:114953559]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	73389847	+	chr17	73401569	+	.	74	43	6497987_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6497987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73377501_73402501_60C;SPAN=11722;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:138 GQ:74.9 PL:[259.7, 0.0, 74.9] SR:43 DR:74 LR:-265.3 LO:265.3);ALT=C[chr17:73401569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76164798	+	chr17	76166897	+	.	87	22	6507342_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6507342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76146001_76171001_95C;SPAN=2099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:81 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:22 DR:87 LR:-277.3 LO:277.3);ALT=T[chr17:76166897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76972290	+	chr17	76975909	+	.	48	0	6510173_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6510173_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76972290(+)-17:76975909(-)__17_76954501_76979501D;SPAN=3619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:89 GQ:81.5 PL:[134.3, 0.0, 81.5] SR:0 DR:48 LR:-135.0 LO:135.0);ALT=C[chr17:76975909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	77393690	+	chr17	77365465	+	.	49	28	6511543_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6511543_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_77371001_77396001_104C;SPAN=28225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:51 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:28 DR:49 LR:-181.5 LO:181.5);ALT=]chr17:77393690]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	79213492	+	chr17	79214785	+	.	39	0	6516554_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6516554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79213492(+)-17:79214785(-)__17_79208501_79233501D;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:85 GQ:99 PL:[105.8, 0.0, 99.2] SR:0 DR:39 LR:-105.7 LO:105.7);ALT=G[chr17:79214785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79827834	+	chr17	79829171	+	.	112	58	6518996_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=6518996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79821001_79846001_191C;SPAN=1337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:94 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:58 DR:112 LR:-373.0 LO:373.0);ALT=C[chr17:79829171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79849982	+	chr17	79851427	+	.	129	6	6518761_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6518761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79845501_79870501_198C;SPAN=1445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:81 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:6 DR:129 LR:-399.4 LO:399.4);ALT=G[chr17:79851427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79849998	+	chr17	79857795	+	.	63	0	6518763_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6518763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79849998(+)-17:79857795(-)__17_79845501_79870501D;SPAN=7797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:124 GQ:99 PL:[174.5, 0.0, 125.0] SR:0 DR:63 LR:-174.8 LO:174.8);ALT=T[chr17:79857795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79977306	+	chr17	79980693	+	.	66	0	6519076_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6519076_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79977306(+)-17:79980693(-)__17_79968001_79993001D;SPAN=3387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:83 GQ:4.1 PL:[195.5, 0.0, 4.1] SR:0 DR:66 LR:-206.2 LO:206.2);ALT=C[chr17:79980693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80009882	+	chr17	80011740	+	.	36	0	6519314_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6519314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80009882(+)-17:80011740(-)__17_79992501_80017501D;SPAN=1858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:45 GQ:1.1 PL:[106.7, 0.0, 1.1] SR:0 DR:36 LR:-112.7 LO:112.7);ALT=C[chr17:80011740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80059743	+	chr17	80064146	+	.	48	6	6519145_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6519145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80041501_80066501_279C;SPAN=4403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:78 GQ:41.6 PL:[147.2, 0.0, 41.6] SR:6 DR:48 LR:-150.5 LO:150.5);ALT=C[chr17:80064146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9102815	+	chr19	53727935	-	.	59	0	6862571_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6862571_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:9102815(+)-19:53727935(+)__19_53704001_53729001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:56 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=G]chr19:53727935];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr18	9475691	+	chr18	9512986	+	.	41	30	6537869_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=6537869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_9506001_9531001_226C;SPAN=37295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:56 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:30 DR:41 LR:-171.6 LO:171.6);ALT=T[chr18:9512986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9914330	+	chr18	9931807	+	.	33	0	6538777_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6538777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:9914330(+)-18:9931807(-)__18_9922501_9947501D;SPAN=17477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:39 GQ:3.9 PL:[102.3, 3.9, 0.0] SR:0 DR:33 LR:-105.5 LO:105.5);ALT=A[chr18:9931807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	10222280	+	chr18	10223605	+	.	59	46	6539080_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=6539080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_10216501_10241501_211C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:42 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:46 DR:59 LR:-267.4 LO:267.4);ALT=A[chr18:10223605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21903397	+	chr18	21904597	+	.	75	0	6562722_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6562722_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:21903397(+)-18:21904597(-)__18_21903001_21928001D;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:182 GQ:99 PL:[198.5, 0.0, 241.4] SR:0 DR:75 LR:-198.3 LO:198.5);ALT=C[chr18:21904597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21990742	+	chr18	21992048	+	.	68	50	6562677_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6562677_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_18_21976501_22001501_37C;SPAN=1306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:44 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:50 DR:68 LR:-267.4 LO:267.4);ALT=C[chr18:21992048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43671855	+	chr18	43678166	+	.	100	0	6609467_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6609467_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:43671855(+)-18:43678166(-)__18_43659001_43684001D;SPAN=6311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:91 GQ:27 PL:[297.0, 27.0, 0.0] SR:0 DR:100 LR:-297.1 LO:297.1);ALT=T[chr18:43678166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47329225	+	chr18	47339836	+	.	32	8	6619096_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=6619096_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_47334001_47359001_192C;SPAN=10611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:8 DR:32 LR:-115.5 LO:115.5);ALT=T[chr18:47339836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	54946737	+	chr18	54948718	+	.	53	46	6635909_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=6635909_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_54929001_54954001_164C;SPAN=1981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:40 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:46 DR:53 LR:-244.3 LO:244.3);ALT=A[chr18:54948718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	57567467	+	chr18	57569876	+	.	34	43	6642667_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6642667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_57550501_57575501_291C;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:83 GQ:20.6 PL:[179.0, 0.0, 20.6] SR:43 DR:34 LR:-185.9 LO:185.9);ALT=G[chr18:57569876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	75266998	+	chr18	75268160	+	.	59	41	6681908_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6681908_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_75264001_75289001_115C;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:42 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:41 DR:59 LR:-250.9 LO:250.9);ALT=T[chr18:75268160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76202137	+	chr18	76203341	+	.	45	34	6683978_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAGATTGATCAAGG;MAPQ=60;MATEID=6683978_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_76195001_76220001_177C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:39 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:34 DR:45 LR:-204.7 LO:204.7);ALT=G[chr18:76203341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76295468	+	chr18	76296725	+	.	61	38	6684283_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=6684283_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_18_76293001_76318001_81C;SPAN=1257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:39 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:38 DR:61 LR:-241.0 LO:241.0);ALT=C[chr18:76296725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	77309950	+	chr18	77312062	+	.	76	18	6686927_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GACAAAGCCTCACAGACCCCCAGACAGGG;MAPQ=60;MATEID=6686927_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_18_77297501_77322501_163C;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:35 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:18 DR:76 LR:-260.8 LO:260.8);ALT=G[chr18:77312062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	572701	+	chr19	579502	+	CT	101	22	6690845_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CT;MAPQ=60;MATEID=6690845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_563501_588501_54C;SPAN=6801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:75 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:22 DR:101 LR:-323.5 LO:323.5);ALT=G[chr19:579502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	692052	+	chr19	695350	+	.	110	0	6691099_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691099_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:692052(+)-19:695350(-)__19_686001_711001D;SPAN=3298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:122 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:0 DR:110 LR:-359.8 LO:359.8);ALT=G[chr19:695350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	902618	+	chr19	913104	+	.	65	0	6691503_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:902618(+)-19:913104(-)__19_882001_907001D;SPAN=10486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:33 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=C[chr19:913104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1026723	+	chr19	1031069	+	.	78	21	6692493_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6692493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1029001_1054001_204C;SPAN=4346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:40 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:21 DR:78 LR:-250.9 LO:250.9);ALT=G[chr19:1031069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1104126	+	chr19	1105184	+	.	173	16	6692418_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6692418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1102501_1127501_158C;SPAN=1058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:184 DP:119 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:16 DR:173 LR:-544.6 LO:544.6);ALT=G[chr19:1105184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1269410	+	chr19	1270926	+	.	55	12	6692834_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6692834_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1249501_1274501_58C;SPAN=1516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:94 GQ:53.9 PL:[172.7, 0.0, 53.9] SR:12 DR:55 LR:-175.9 LO:175.9);ALT=G[chr19:1270926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1269417	+	chr19	1271135	+	.	116	0	6692835_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6692835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1269417(+)-19:1271135(-)__19_1249501_1274501D;SPAN=1718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:127 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:0 DR:116 LR:-376.3 LO:376.3);ALT=C[chr19:1271135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1383993	+	chr19	1388541	+	.	85	0	6693399_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6693399_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1383993(+)-19:1388541(-)__19_1372001_1397001D;SPAN=4548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:120 GQ:43.4 PL:[248.0, 0.0, 43.4] SR:0 DR:85 LR:-256.3 LO:256.3);ALT=G[chr19:1388541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1383995	+	chr19	1390866	+	.	37	0	6693400_1	94.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6693400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1383995(+)-19:1390866(-)__19_1372001_1397001D;SPAN=6871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:103 GQ:94.4 PL:[94.4, 0.0, 153.8] SR:0 DR:37 LR:-94.23 LO:95.06);ALT=A[chr19:1390866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1598263	+	chr19	1605361	+	.	61	0	6694010_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6694010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1598263(+)-19:1605361(-)__19_1592501_1617501D;SPAN=7098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:91 GQ:41.6 PL:[176.9, 0.0, 41.6] SR:0 DR:61 LR:-181.2 LO:181.2);ALT=G[chr19:1605361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1599560	+	chr19	1605358	+	.	75	24	6694017_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6694017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1592501_1617501_289C;SPAN=5798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:114 GQ:25.4 PL:[249.8, 0.0, 25.4] SR:24 DR:75 LR:-260.2 LO:260.2);ALT=C[chr19:1605358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2236932	+	chr19	2243377	+	.	46	0	6696056_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6696056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2236932(+)-19:2243377(-)__19_2229501_2254501D;SPAN=6445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:75 GQ:49.1 PL:[131.6, 0.0, 49.1] SR:0 DR:46 LR:-133.5 LO:133.5);ALT=C[chr19:2243377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2269744	+	chr19	2271779	+	.	34	4	6696469_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6696469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2254001_2279001_360C;SPAN=2035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:216 GQ:99 PL:[109.9, 0.0, 413.6] SR:4 DR:34 LR:-109.8 LO:119.8);ALT=G[chr19:2271779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2270247	+	chr19	2271381	+	.	111	0	6696475_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6696475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2270247(+)-19:2271381(-)__19_2254001_2279001D;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:195 GQ:99 PL:[313.7, 0.0, 158.6] SR:0 DR:111 LR:-316.3 LO:316.3);ALT=G[chr19:2271381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2349583	+	chr19	2348175	+	.	44	0	6696649_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6696649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2348175(-)-19:2349583(+)__19_2327501_2352501D;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:73 GQ:49.7 PL:[125.6, 0.0, 49.7] SR:0 DR:44 LR:-127.1 LO:127.1);ALT=]chr19:2349583]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	2737680	+	chr19	2739942	+	.	58	0	6697898_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6697898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2737680(+)-19:2739942(-)__19_2719501_2744501D;SPAN=2262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:81 GQ:24.5 PL:[169.7, 0.0, 24.5] SR:0 DR:58 LR:-175.4 LO:175.4);ALT=T[chr19:2739942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3474996	+	chr19	3478417	+	.	51	6	6700826_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6700826_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_3454501_3479501_216C;SPAN=3421;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:81 GQ:27.8 PL:[166.4, 0.0, 27.8] SR:6 DR:51 LR:-171.5 LO:171.5);ALT=T[chr19:3478417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3762816	+	chr19	3765160	+	.	83	45	6701650_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAG;MAPQ=60;MATEID=6701650_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_3748501_3773501_150C;SPAN=2344;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:100 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:45 DR:83 LR:-303.7 LO:303.7);ALT=G[chr19:3765160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3983336	+	chr19	3985399	+	.	75	0	6702679_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6702679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3983336(+)-19:3985399(-)__19_3969001_3994001D;SPAN=2063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:245 GQ:99 PL:[181.3, 0.0, 412.4] SR:0 DR:75 LR:-181.2 LO:186.2);ALT=G[chr19:3985399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3984349	+	chr19	3985372	+	.	161	23	6702686_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCACC;MAPQ=60;MATEID=6702686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3969001_3994001_329C;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:168 DP:110 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:23 DR:161 LR:-498.4 LO:498.4);ALT=C[chr19:3985372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4665004	+	chr19	4670171	+	.	37	0	6704965_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6704965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4665004(+)-19:4670171(-)__19_4655001_4680001D;SPAN=5167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:80 GQ:93.8 PL:[100.4, 0.0, 93.8] SR:0 DR:37 LR:-100.5 LO:100.5);ALT=C[chr19:4670171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4668715	+	chr19	4670269	+	.	57	0	6704978_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6704978_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4668715(+)-19:4670269(-)__19_4655001_4680001D;SPAN=1554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:75 GQ:12.8 PL:[167.9, 0.0, 12.8] SR:0 DR:57 LR:-175.5 LO:175.5);ALT=A[chr19:4670269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4860074	+	chr19	4867619	+	.	62	0	6705652_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6705652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4860074(+)-19:4867619(-)__19_4851001_4876001D;SPAN=7545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:101 GQ:65.3 PL:[177.5, 0.0, 65.3] SR:0 DR:62 LR:-180.0 LO:180.0);ALT=G[chr19:4867619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5896795	+	chr19	5903677	+	.	47	0	6709409_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6709409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:5896795(+)-19:5903677(-)__19_5880001_5905001D;SPAN=6882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:132 GQ:99 PL:[119.6, 0.0, 198.8] SR:0 DR:47 LR:-119.4 LO:120.5);ALT=G[chr19:5903677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6373036	+	chr19	6374213	+	.	67	89	6711229_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6711229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_6370001_6395001_254C;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:137 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:89 DR:67 LR:-406.0 LO:406.0);ALT=G[chr19:6374213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7702112	+	chr19	7704615	+	.	35	0	6715787_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6715787_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7702112(+)-19:7704615(-)__19_7693001_7718001D;SPAN=2503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:90 GQ:91.1 PL:[91.1, 0.0, 127.4] SR:0 DR:35 LR:-91.15 LO:91.48);ALT=G[chr19:7704615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7745936	+	chr19	7747126	+	.	115	7	6715859_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6715859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_7742001_7767001_141C;SPAN=1190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:120 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:7 DR:115 LR:-356.5 LO:356.5);ALT=G[chr19:7747126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8056718	+	chr19	8070379	+	.	52	20	6717081_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6717081_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8060501_8085501_245C;SPAN=13661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:6 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:20 DR:52 LR:-178.2 LO:178.2);ALT=G[chr19:8070379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8381530	+	chr19	8386192	+	GCTTGGAGATCTCCTGGTAGCGTAGCTGCAGCTTCCCCTGCAGGTCATG	74	28	6718260_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GCTTGGAGATCTCCTGGTAGCGTAGCTGCAGCTTCCCCTGCAGGTCATG;MAPQ=60;MATEID=6718260_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8379001_8404001_277C;SPAN=4662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:99 GQ:6.9 PL:[254.1, 6.9, 0.0] SR:28 DR:74 LR:-264.3 LO:264.3);ALT=C[chr19:8386192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8455340	+	chr19	8464745	+	.	85	4	6718532_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6718532_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8452501_8477501_184C;SPAN=9405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:94 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:4 DR:85 LR:-277.3 LO:277.3);ALT=G[chr19:8464745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8509995	+	chr19	8520288	+	.	41	16	6718641_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6718641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8501501_8526501_363C;SPAN=10293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:89 GQ:88.1 PL:[127.7, 0.0, 88.1] SR:16 DR:41 LR:-128.1 LO:128.1);ALT=G[chr19:8520288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8564665	+	chr19	8567448	+	.	53	4	6718945_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6718945_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_8550501_8575501_130C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:106 GQ:99 PL:[152.9, 0.0, 103.4] SR:4 DR:53 LR:-153.3 LO:153.3);ALT=C[chr19:8567448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9274508	+	chr19	9042090	+	.	36	0	6721691_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6721691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:9042090(-)-19:9274508(+)__19_9261001_9286001D;SPAN=232418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:16 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=]chr19:9274508]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	9946079	+	chr19	9949109	+	.	97	4	6725345_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6725345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_9922501_9947501_61C;SPAN=3030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:54 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:4 DR:97 LR:-290.5 LO:290.5);ALT=G[chr19:9949109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10229453	+	chr19	10230513	+	.	35	0	6726433_1	80.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6726433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10229453(+)-19:10230513(-)__19_10216501_10241501D;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:132 GQ:80 PL:[80.0, 0.0, 238.4] SR:0 DR:35 LR:-79.77 LO:84.27);ALT=C[chr19:10230513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10291618	+	chr19	10305517	+	.	70	0	6726615_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6726615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10291618(+)-19:10305517(-)__19_10290001_10315001D;SPAN=13899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:89 GQ:8.9 PL:[206.9, 0.0, 8.9] SR:0 DR:70 LR:-217.9 LO:217.9);ALT=A[chr19:10305517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10506882	+	chr19	10514053	+	.	144	67	6727689_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6727689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10486001_10511001_172C;SPAN=7171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:178 DP:60 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:67 DR:144 LR:-528.1 LO:528.1);ALT=G[chr19:10514053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77359862	+	chr19	12670380	+	.	134	0	7455522_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=7455522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12670380(-)-23:77359862(+)__23_77346501_77371501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:50 GQ:36 PL:[396.0, 36.0, 0.0] SR:0 DR:134 LR:-396.1 LO:396.1);ALT=]chrX:77359862]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	12694884	+	chr19	12698931	+	.	89	76	6735358_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=GCCTCCCA;MAPQ=0;MATEID=6735358_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12691001_12716001_27C;SPAN=4047;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:32 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:76 DR:89 LR:-415.9 LO:415.9);ALT=A[chr19:12698931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13041565	+	chr19	13044362	+	.	41	19	6736517_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6736517_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_13034001_13059001_196C;SPAN=2797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:95 GQ:99 PL:[129.5, 0.0, 99.8] SR:19 DR:41 LR:-129.6 LO:129.6);ALT=T[chr19:13044362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13056774	+	chr19	13058660	+	.	82	0	6736751_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6736751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:13056774(+)-19:13058660(-)__19_13058501_13083501D;SPAN=1886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:38 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=C[chr19:13058660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13885521	+	chr19	13888864	+	.	105	63	6739548_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6739548_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_19_13867001_13892001_36C;SPAN=3343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:121 GQ:37.7 PL:[327.7, 37.7, 0.0] SR:63 DR:105 LR:-327.7 LO:327.7);ALT=G[chr19:13888864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14492357	+	chr19	14499261	+	.	65	33	6742295_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=G;MAPQ=58;MATEID=6742295_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_19_14479501_14504501_10C;SPAN=6904;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:106 GQ:21.9 PL:[300.3, 21.9, 0.0] SR:33 DR:65 LR:-302.1 LO:302.1);ALT=G[chr19:14499261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14499260	-	chr19	14887590	+	.	47	0	6742323_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6742323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14499260(-)-19:14887590(-)__19_14479501_14504501D;SPAN=388330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:55 GQ:8.1 PL:[148.5, 8.1, 0.0] SR:0 DR:47 LR:-150.8 LO:150.8);ALT=[chr19:14887590[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	14524083	+	chr19	14530081	+	.	37	0	6742376_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6742376_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14524083(+)-19:14530081(-)__19_14528501_14553501D;SPAN=5998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:64 GQ:48.8 PL:[104.9, 0.0, 48.8] SR:0 DR:37 LR:-105.8 LO:105.8);ALT=G[chr19:14530081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14732345	+	chr19	14734127	+	.	63	36	6743190_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TAAAACTCCTGGACTT;MAPQ=60;MATEID=6743190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14724501_14749501_298C;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:127 GQ:54.8 PL:[252.8, 0.0, 54.8] SR:36 DR:63 LR:-259.9 LO:259.9);ALT=T[chr19:14734127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16254586	+	chr19	16259529	+	.	66	14	6747887_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCCAGGT;MAPQ=60;MATEID=6747887_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16243501_16268501_339C;SPAN=4943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:136 GQ:99 PL:[200.9, 0.0, 128.3] SR:14 DR:66 LR:-201.7 LO:201.7);ALT=T[chr19:16259529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16254627	+	chr19	16263361	+	.	67	0	6747889_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6747889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16254627(+)-19:16263361(-)__19_16243501_16268501D;SPAN=8734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:118 GQ:96.8 PL:[189.2, 0.0, 96.8] SR:0 DR:67 LR:-190.8 LO:190.8);ALT=G[chr19:16263361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16308881	+	chr19	16314268	+	.	37	20	6748229_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6748229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16292501_16317501_235C;SPAN=5387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:84 GQ:69.8 PL:[132.5, 0.0, 69.8] SR:20 DR:37 LR:-133.4 LO:133.4);ALT=T[chr19:16314268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16435814	+	chr19	16437665	+	.	31	19	6748677_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTGAG;MAPQ=60;MATEID=6748677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16415001_16440001_342C;SPAN=1851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:108 GQ:99 PL:[129.2, 0.0, 132.5] SR:19 DR:31 LR:-129.2 LO:129.2);ALT=G[chr19:16437665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17378336	+	chr19	17379601	+	.	84	3	6752067_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6752067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_17370501_17395501_112C;SPAN=1265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:81 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:3 DR:84 LR:-247.6 LO:247.6);ALT=G[chr19:17379601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18043908	+	chr19	18053462	+	.	40	0	6754374_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6754374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18043908(+)-19:18053462(-)__19_18032001_18057001D;SPAN=9554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:0 DR:40 LR:-109.9 LO:109.9);ALT=C[chr19:18053462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18284783	+	chr19	18285848	+	.	82	66	6755349_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6755349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18277001_18302001_56C;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:118 DP:152 GQ:18.5 PL:[348.5, 0.0, 18.5] SR:66 DR:82 LR:-365.7 LO:365.7);ALT=G[chr19:18285848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18420721	+	chr19	18433825	+	.	79	0	6755900_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6755900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18420721(+)-19:18433825(-)__19_18424001_18449001D;SPAN=13104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:49 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=C[chr19:18433825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18423569	+	chr19	18433825	+	.	93	0	6755769_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6755769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18423569(+)-19:18433825(-)__19_18399501_18424501D;SPAN=10256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:31 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:93 LR:-274.0 LO:274.0);ALT=C[chr19:18433825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18652807	+	chr19	18654295	+	.	137	12	6756974_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6756974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18644501_18669501_231C;SPAN=1488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:97 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:12 DR:137 LR:-422.5 LO:422.5);ALT=T[chr19:18654295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18668772	+	chr19	18675678	+	.	53	0	6757075_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6757075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18668772(+)-19:18675678(-)__19_18669001_18694001D;SPAN=6906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:53 LR:-161.7 LO:161.7);ALT=A[chr19:18675678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18682766	+	chr19	18685677	+	.	35	0	6757135_1	55.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6757135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18682766(+)-19:18685677(-)__19_18669001_18694001D;SPAN=2911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:220 GQ:55.9 PL:[55.9, 0.0, 478.4] SR:0 DR:35 LR:-55.93 LO:75.45);ALT=G[chr19:18685677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19021941	+	chr19	19030031	+	.	90	0	6758114_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6758114_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19021941(+)-19:19030031(-)__19_19012001_19037001D;SPAN=8090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:93 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:90 LR:-274.0 LO:274.0);ALT=G[chr19:19030031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19023906	+	chr19	19030103	+	.	81	0	6758130_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6758130_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19023906(+)-19:19030103(-)__19_19012001_19037001D;SPAN=6197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:85 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:0 DR:81 LR:-250.9 LO:250.9);ALT=C[chr19:19030103[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19049859	+	chr19	19051859	+	.	34	8	6758350_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6758350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_19036501_19061501_239C;SPAN=2000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:61 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:8 DR:34 LR:-107.1 LO:107.1);ALT=C[chr19:19051859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19627142	+	chr19	19636990	+	.	87	42	6760414_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6760414_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_19_19624501_19649501_44C;SPAN=9848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:173 DP:102 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:42 DR:87 LR:-511.6 LO:511.6);ALT=G[chr19:19636990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24595035	+	chr19	24596046	+	.	38	23	6775996_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTCTTTTTGTAGAATCT;MAPQ=60;MATEID=6775996_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_19_24573501_24598501_452C;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:72 GQ:13.7 PL:[158.9, 0.0, 13.7] SR:23 DR:38 LR:-165.6 LO:165.6);ALT=T[chr19:24596046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	30388804	+	chr19	30393101	+	.	80	41	6783648_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TAATTTTTATTTTT;MAPQ=60;MATEID=6783648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_30380001_30405001_173C;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:78 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:41 DR:80 LR:-277.3 LO:277.3);ALT=T[chr19:30393101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35645772	+	chr19	35648322	+	ATGTCGCCCTCTGGTCGCCTGTGTCTTCTCACCATCGTTGGCCTGATTCTCCCCACCAG	73	73	6798452_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGTCGCCCTCTGGTCGCCTGTGTCTTCTCACCATCGTTGGCCTGATTCTCCCCACCAG;MAPQ=60;MATEID=6798452_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_19_35623001_35648001_50C;SPAN=2550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:53 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:73 DR:73 LR:-432.4 LO:432.4);ALT=G[chr19:35648322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36139306	+	chr19	36145472	+	ATTCAGCACCATGGCGGAAGACATGGAGACCAAAATCAAGAACTACAAGACCGCCCCTTTTGACAGCCGCTTCCCCAACCAGAACCAGACTAGAAACTGCTGGCAGAACTACCTG	97	188	6800245_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATTCAGCACCATGGCGGAAGACATGGAGACCAAAATCAAGAACTACAAGACCGCCCCTTTTGACAGCCGCTTCCCCAACCAGAACCAGACTAGAAACTGCTGGCAGAACTACCTG;MAPQ=60;MATEID=6800245_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36137501_36162501_282C;SPAN=6166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:266 DP:218 GQ:71.8 PL:[788.8, 71.8, 0.0] SR:188 DR:97 LR:-788.9 LO:788.9);ALT=G[chr19:36145472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36139306	+	chr19	36142133	+	.	56	9	6800244_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6800244_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_36137501_36162501_282C;SPAN=2827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:159 GQ:79.1 PL:[306.8, 0.0, 79.1] SR:9 DR:56 LR:-314.3 LO:314.3);ALT=G[chr19:36142133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36232120	+	chr19	36233290	+	.	77	0	6799896_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6799896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36232120(+)-19:36233290(-)__19_36211001_36236001D;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:87 GQ:20.1 PL:[250.8, 20.1, 0.0] SR:0 DR:77 LR:-251.3 LO:251.3);ALT=C[chr19:36233290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36637217	+	chr19	36640713	+	CCTTCAAATCTCTTGACAAAGATGGCACTGGACAAATCCAGGTGAACATCCAGG	32	35	6801457_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCTTCAAATCTCTTGACAAAGATGGCACTGGACAAATCCAGGTGAACATCCAGG;MAPQ=60;MATEID=6801457_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_19_36627501_36652501_378C;SPAN=3496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:90 GQ:71.3 PL:[147.2, 0.0, 71.3] SR:35 DR:32 LR:-148.7 LO:148.7);ALT=G[chr19:36640713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38800319	+	chr19	38806356	+	.	80	0	6810009_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6810009_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:38800319(+)-19:38806356(-)__19_38783501_38808501D;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:97 GQ:3 PL:[240.9, 3.0, 0.0] SR:0 DR:80 LR:-253.2 LO:253.2);ALT=C[chr19:38806356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39109979	+	chr19	39114716	+	.	81	0	6811129_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6811129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39109979(+)-19:39114716(-)__19_39102001_39127001D;SPAN=4737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:125 GQ:68.6 PL:[233.6, 0.0, 68.6] SR:0 DR:81 LR:-238.4 LO:238.4);ALT=G[chr19:39114716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39820312	+	chr19	39826613	+	.	45	0	6813754_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6813754_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39820312(+)-19:39826613(-)__19_39812501_39837501D;SPAN=6301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:176 GQ:99 PL:[101.0, 0.0, 325.4] SR:0 DR:45 LR:-100.9 LO:107.5);ALT=A[chr19:39826613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39824149	+	chr19	39826613	+	.	67	0	6813771_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6813771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39824149(+)-19:39826613(-)__19_39812501_39837501D;SPAN=2464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:170 GQ:99 PL:[175.1, 0.0, 237.8] SR:0 DR:67 LR:-175.1 LO:175.6);ALT=G[chr19:39826613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39924437	+	chr19	39926494	+	.	78	0	6814131_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6814131_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39924437(+)-19:39926494(-)__19_39910501_39935501D;SPAN=2057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:123 GQ:72.5 PL:[224.3, 0.0, 72.5] SR:0 DR:78 LR:-228.3 LO:228.3);ALT=C[chr19:39926494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40331430	+	chr19	40336930	+	.	186	12	6815089_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6815089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40327001_40352001_248C;SPAN=5500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:193 DP:91 GQ:52 PL:[571.0, 52.0, 0.0] SR:12 DR:186 LR:-571.0 LO:571.0);ALT=G[chr19:40336930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40854678	+	chr19	40871458	+	.	38	2	6817119_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=6817119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40841501_40866501_234C;SPAN=16780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:2 DR:38 LR:-120.9 LO:120.9);ALT=A[chr19:40871458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40964455	+	chr19	40971516	+	.	85	41	6817279_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6817279_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40964001_40989001_233C;SPAN=7061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:102 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:41 DR:85 LR:-303.7 LO:303.7);ALT=G[chr19:40971516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41903840	+	chr19	41916550	+	CACCCCCA	37	10	6820662_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CACCCCCA;MAPQ=60;MATEID=6820662_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41895001_41920001_221C;SPAN=12710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:97 GQ:99 PL:[109.1, 0.0, 125.6] SR:10 DR:37 LR:-109.1 LO:109.1);ALT=T[chr19:41916550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44118603	+	chr19	44123709	+	.	87	0	6827570_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6827570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:44118603(+)-19:44123709(-)__19_44100001_44125001D;SPAN=5106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:88 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:0 DR:87 LR:-260.8 LO:260.8);ALT=G[chr19:44123709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45668229	+	chr19	45681392	+	.	77	3	6832621_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6832621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45643501_45668501_27C;SPAN=13163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:61 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:3 DR:77 LR:-234.4 LO:234.4);ALT=C[chr19:45681392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45668453	+	chr19	45681392	+	.	33	9	6832761_1	81.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6832761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45668001_45693001_348C;SPAN=12939;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:115 GQ:81.2 PL:[81.2, 0.0, 196.7] SR:9 DR:33 LR:-81.08 LO:83.78);ALT=C[chr19:45681392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46191011	+	chr19	46195142	+	.	32	0	6834934_1	60.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6834934_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46191011(+)-19:46195142(-)__19_46182501_46207501D;SPAN=4131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:166 GQ:60.8 PL:[60.8, 0.0, 341.3] SR:0 DR:32 LR:-60.66 LO:71.95);ALT=A[chr19:46195142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46191852	+	chr19	46195141	+	.	139	0	6834939_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6834939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46191852(+)-19:46195141(-)__19_46182501_46207501D;SPAN=3289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:158 GQ:32.8 PL:[448.9, 32.8, 0.0] SR:0 DR:139 LR:-452.2 LO:452.2);ALT=G[chr19:46195141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47104695	+	chr19	47111451	+	CTGACCAGCTGACTGAGGAGCAGATTG	95	58	6837877_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTGACCAGCTGACTGAGGAGCAGATTG;MAPQ=60;MATEID=6837877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47089001_47114001_115C;SPAN=6756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:78 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:58 DR:95 LR:-346.6 LO:346.6);ALT=G[chr19:47111451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47342909	+	chr19	47354019	+	.	87	0	6839008_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6839008_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:47342909(+)-19:47354019(-)__19_47334001_47359001D;SPAN=11110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:91 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:0 DR:87 LR:-267.4 LO:267.4);ALT=T[chr19:47354019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47349400	+	chr19	47354021	+	.	108	18	6839035_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6839035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47334001_47359001_269C;SPAN=4621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:104 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:18 DR:108 LR:-340.0 LO:340.0);ALT=C[chr19:47354021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48828868	+	chr19	48830086	+	.	43	72	6844163_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6844163_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48804001_48829001_26C;SPAN=1218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:115 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:72 DR:43 LR:-340.0 LO:340.0);ALT=G[chr19:48830086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49404124	+	chr19	49407602	+	.	44	0	6847145_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847145_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49404124(+)-19:49407602(-)__19_49392001_49417001D;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:130 GQ:99 PL:[110.0, 0.0, 205.7] SR:0 DR:44 LR:-110.0 LO:111.6);ALT=T[chr19:49407602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49839044	+	chr19	49840165	+	.	46	113	6849161_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6849161_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_49833001_49858001_283C;SPAN=1121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:129 DP:184 GQ:69.1 PL:[376.1, 0.0, 69.1] SR:113 DR:46 LR:-387.8 LO:387.8);ALT=G[chr19:49840165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50180613	+	chr19	50185162	+	.	53	0	6850109_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6850109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50180613(+)-19:50185162(-)__19_50176001_50201001D;SPAN=4549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:69 GQ:11 PL:[156.2, 0.0, 11.0] SR:0 DR:53 LR:-163.7 LO:163.7);ALT=T[chr19:50185162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50840933	+	chr19	50847929	+	.	124	15	6852589_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6852589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50837501_50862501_102C;SPAN=6996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:99 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:15 DR:124 LR:-382.9 LO:382.9);ALT=C[chr19:50847929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50979916	+	chr19	50982213	+	CTGGGGCGGAAGGTCGAGAGGGCGAGGCCTGTGGCACGGTGGGGCTGCTGCTGGAGCACTCATTTGAGATC	41	67	6852878_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTGGGGCGGAAGGTCGAGAGGGCGAGGCCTGTGGCACGGTGGGGCTGCTGCTGGAGCACTCATTTGAGATC;MAPQ=60;MATEID=6852878_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_50960001_50985001_164C;SPAN=2297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:102 GQ:17.4 PL:[280.5, 17.4, 0.0] SR:67 DR:41 LR:-283.6 LO:283.6);ALT=G[chr19:50982213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51302260	+	chr19	51305475	+	.	54	0	6855161_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6855161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51302260(+)-19:51305475(-)__19_51278501_51303501D;SPAN=3215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:41 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=C[chr19:51305475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51856597	+	chr19	51869525	+	.	54	0	6857157_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6857157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51856597(+)-19:51869525(-)__19_51866501_51891501D;SPAN=12928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:56 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:54 LR:-165.0 LO:165.0);ALT=A[chr19:51869525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51857564	+	chr19	51869524	+	.	143	30	6857158_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6857158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51866501_51891501_197C;SPAN=11960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:55 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:30 DR:143 LR:-429.1 LO:429.1);ALT=T[chr19:51869524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52175937	+	chr19	52177514	+	.	60	30	6857843_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAATTTTC;MAPQ=60;MATEID=6857843_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_19_52160501_52185501_270C;SPAN=1577;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:31 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:30 DR:60 LR:-244.3 LO:244.3);ALT=C[chr19:52177514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52693419	+	chr19	52709211	+	.	50	0	6859425_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6859425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52693419(+)-19:52709211(-)__19_52675001_52700001D;SPAN=15792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:43 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=G[chr19:52709211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52693427	+	chr19	52705195	+	.	48	32	6859426_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6859426_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52675001_52700001_321C;SPAN=11768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:39 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:32 DR:48 LR:-181.5 LO:181.5);ALT=G[chr19:52705195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53096022	+	chr19	53097609	+	.	94	28	6860645_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTAATTTTGTATTTTT;MAPQ=60;MATEID=6860645_2;MATENM=2;NM=5;NUMPARTS=2;SCTG=c_19_53091501_53116501_68C;SPAN=1587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:25 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:28 DR:94 LR:-320.2 LO:320.2);ALT=T[chr19:53097609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53422211	+	chr19	53424207	+	.	66	20	6862139_1	84.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAA;MAPQ=60;MATEID=6862139_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_53410001_53435001_234C;SPAN=1996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:640 GQ:84.1 PL:[84.1, 0.0, 1470.0] SR:20 DR:66 LR:-84.09 LO:158.4);ALT=A[chr19:53424207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54371200	+	chr19	54376781	+	CTCTTACAGCCTGTTCCAAGTGTGGCTTAATCCGTCTCCACCACCAGATCTTTCTCCGTGGATTCCTCTGCTAAGACCGCT	114	46	6865218_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTCTTACAGCCTGTTCCAAGTGTGGCTTAATCCGTCTCCACCACCAGATCTTTCTCCGTGGATTCCTCTGCTAAGACCGCT;MAPQ=60;MATEID=6865218_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54365501_54390501_220C;SPAN=5581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:157 GQ:32.5 PL:[445.6, 32.5, 0.0] SR:46 DR:114 LR:-448.7 LO:448.7);ALT=G[chr19:54376781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54373092	+	chr19	54376781	+	.	44	41	6865225_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6865225_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54365501_54390501_220C;SPAN=3689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:105 GQ:11.3 PL:[242.3, 0.0, 11.3] SR:41 DR:44 LR:-254.6 LO:254.6);ALT=G[chr19:54376781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54428719	+	chr19	54426619	+	.	41	0	6865939_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6865939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54426619(-)-19:54428719(+)__19_54414501_54439501D;SPAN=2100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:130 GQ:99 PL:[100.1, 0.0, 215.6] SR:0 DR:41 LR:-100.1 LO:102.4);ALT=]chr19:54428719]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54606496	+	chr19	54609240	+	.	37	49	6866525_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6866525_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54586001_54611001_271C;SPAN=2744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:132 GQ:99 PL:[212.0, 0.0, 106.4] SR:49 DR:37 LR:-213.6 LO:213.6);ALT=G[chr19:54609240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54606545	+	chr19	54610112	+	.	64	0	6866526_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6866526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54606545(+)-19:54610112(-)__19_54586001_54611001D;SPAN=3567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:134 GQ:99 PL:[175.1, 0.0, 148.7] SR:0 DR:64 LR:-175.1 LO:175.1);ALT=C[chr19:54610112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54872898	+	chr19	54876380	+	.	46	0	6867202_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6867202_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54872898(+)-19:54876380(-)__19_54855501_54880501D;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:103 GQ:99 PL:[124.1, 0.0, 124.1] SR:0 DR:46 LR:-123.9 LO:123.9);ALT=A[chr19:54876380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	55967857	+	chr19	55972879	+	.	41	19	6871088_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6871088_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_55958001_55983001_289C;SPAN=5022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:106 GQ:99 PL:[123.2, 0.0, 133.1] SR:19 DR:41 LR:-123.1 LO:123.2);ALT=C[chr19:55972879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56111826	+	chr19	56113436	+	.	33	0	6871337_1	89.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6871337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:56111826(+)-19:56113436(-)__19_56105001_56130001D;SPAN=1610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:72 GQ:83 PL:[89.6, 0.0, 83.0] SR:0 DR:33 LR:-89.43 LO:89.43);ALT=A[chr19:56113436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56186801	+	chr19	56189891	+	.	36	33	6871691_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6871691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_56178501_56203501_40C;SPAN=3090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:93 GQ:80.6 PL:[143.3, 0.0, 80.6] SR:33 DR:36 LR:-144.0 LO:144.0);ALT=G[chr19:56189891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58898735	+	chr19	58904339	+	.	57	0	6880845_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6880845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:58898735(+)-19:58904339(-)__19_58898001_58923001D;SPAN=5604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:149 GQ:99 PL:[147.8, 0.0, 213.8] SR:0 DR:57 LR:-147.8 LO:148.5);ALT=A[chr19:58904339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	59063806	+	chr19	59065411	+	.	45	58	6880793_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6880793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_59045001_59070001_254C;SPAN=1605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:110 GQ:16.4 PL:[250.7, 0.0, 16.4] SR:58 DR:45 LR:-263.1 LO:263.1);ALT=C[chr19:59065411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1389146	+	chr20	1390815	+	.	67	38	6886506_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=6886506_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_20_1372001_1397001_298C;SPAN=1669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:94 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:38 DR:67 LR:-277.3 LO:277.3);ALT=A[chr20:1390815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2446514	+	chr20	2451333	+	.	49	0	6890323_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6890323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:2446514(+)-20:2451333(-)__20_2450001_2475001D;SPAN=4819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:58 GQ:5.7 PL:[151.8, 5.7, 0.0] SR:0 DR:49 LR:-156.5 LO:156.5);ALT=G[chr20:2451333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2448405	+	chr20	2451334	+	.	118	27	6890324_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6890324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2450001_2475001_216C;SPAN=2929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:59 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:27 DR:118 LR:-373.0 LO:373.0);ALT=C[chr20:2451334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2803162	+	chr20	2806410	+	.	49	34	6891520_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAGAACTTGATTT;MAPQ=60;MATEID=6891520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2793001_2818001_85C;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:87 GQ:2.9 PL:[207.5, 0.0, 2.9] SR:34 DR:49 LR:-219.6 LO:219.6);ALT=T[chr20:2806410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3184065	+	chr20	3185183	+	.	37	17	6893221_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6893221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3160501_3185501_215C;SPAN=1118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:125 GQ:99 PL:[118.1, 0.0, 184.1] SR:17 DR:37 LR:-118.0 LO:118.8);ALT=G[chr20:3185183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3190265	+	chr20	3193813	+	.	40	12	6893356_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=6893356_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_3185001_3210001_191C;SPAN=3548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:113 GQ:99 PL:[108.2, 0.0, 164.3] SR:12 DR:40 LR:-108.0 LO:108.7);ALT=T[chr20:3193813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3740835	+	chr20	3748309	+	.	32	11	6895379_1	82.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6895379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3724001_3749001_394C;SPAN=7474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:99 GQ:82.1 PL:[82.1, 0.0, 158.0] SR:11 DR:32 LR:-82.11 LO:83.43);ALT=T[chr20:3748309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16710805	+	chr20	16712805	+	.	38	0	6938933_1	94.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6938933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:16710805(+)-20:16712805(-)__20_16709001_16734001D;SPAN=2000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:114 GQ:94.7 PL:[94.7, 0.0, 180.5] SR:0 DR:38 LR:-94.55 LO:96.07);ALT=C[chr20:16712805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	17550857	+	chr20	17581382	+	.	38	14	6941437_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6941437_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_20_17542001_17567001_402C;SECONDARY;SPAN=30525;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:45 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:14 DR:38 LR:-151.8 LO:151.8);ALT=G[chr20:17581382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	18191155	+	chr20	18189739	+	.	34	0	6944072_1	90.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6944072_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:18189739(-)-20:18191155(+)__20_18179001_18204001D;SPAN=1416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:80 GQ:90.5 PL:[90.5, 0.0, 103.7] SR:0 DR:34 LR:-90.56 LO:90.61);ALT=]chr20:18191155]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	18548240	+	chr20	18549881	+	.	78	50	6945633_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6945633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_18546501_18571501_261C;SPAN=1641;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:151 GQ:74.9 PL:[289.4, 0.0, 74.9] SR:50 DR:78 LR:-296.0 LO:296.0);ALT=G[chr20:18549881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	20336634	+	chr20	20335485	+	.	32	0	6951625_1	75.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6951625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:20335485(-)-20:20336634(+)__20_20335001_20360001D;SPAN=1149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:112 GQ:75.5 PL:[75.5, 0.0, 194.3] SR:0 DR:32 LR:-75.29 LO:78.28);ALT=]chr20:20336634]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	21284111	+	chr20	21306915	+	.	87	22	6954551_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6954551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_21290501_21315501_193C;SPAN=22804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:57 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:22 DR:87 LR:-270.7 LO:270.7);ALT=G[chr20:21306915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	21286127	+	chr20	21288773	+	.	98	40	6954360_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCATGTTGGCCAGGCTGGTCTCGAACTCCTGACCTCA;MAPQ=60;MATEID=6954360_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_20_21266001_21291001_41C;SPAN=2646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:29 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:40 DR:98 LR:-382.9 LO:382.9);ALT=A[chr20:21288773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31316016	+	chr20	31331112	+	.	130	0	6979298_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6979298_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31316016(+)-20:31331112(-)__20_31311001_31336001D;SPAN=15096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:130 DP:126 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:0 DR:130 LR:-386.2 LO:386.2);ALT=G[chr20:31331112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32581940	+	chr20	32659871	+	.	34	4	6985114_1	97.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6985114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32658501_32683501_315C;SPAN=77931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:79 GQ:94.1 PL:[97.4, 0.0, 94.1] SR:4 DR:34 LR:-97.44 LO:97.44);ALT=G[chr20:32659871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32581942	+	chr20	32619327	+	.	40	53	6984726_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGAG;MAPQ=60;MATEID=6984726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32560501_32585501_62C;SPAN=37385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:60 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:53 DR:40 LR:-208.0 LO:208.0);ALT=G[chr20:32619327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32815938	+	chr20	32819226	+	.	78	25	6985680_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAGAACTTTC;MAPQ=60;MATEID=6985680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32805501_32830501_34C;SPAN=3288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:109 DP:610 GQ:99 PL:[194.6, 0.0, 1287.0] SR:25 DR:78 LR:-194.5 LO:241.1);ALT=C[chr20:32819226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32883392	+	chr20	32891049	+	.	91	15	6985741_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6985741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32879001_32904001_160C;SPAN=7657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:109 GQ:19.5 PL:[303.6, 19.5, 0.0] SR:15 DR:91 LR:-307.6 LO:307.6);ALT=C[chr20:32891049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33104318	+	chr20	33122429	+	.	61	0	6987147_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6987147_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33104318(+)-20:33122429(-)__20_33099501_33124501D;SPAN=18111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:113 GQ:99 PL:[170.9, 0.0, 101.6] SR:0 DR:61 LR:-171.6 LO:171.6);ALT=A[chr20:33122429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34220846	+	chr20	34252682	+	.	72	17	6991850_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6991850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34202001_34227001_425C;SPAN=31836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:76 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:17 DR:72 LR:-227.8 LO:227.8);ALT=C[chr20:34252682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47836079	+	chr20	47837987	+	.	48	17	7042751_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7042751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47824001_47849001_305C;SPAN=1908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:127 GQ:99 PL:[143.9, 0.0, 163.7] SR:17 DR:48 LR:-143.8 LO:143.9);ALT=G[chr20:47837987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47895263	+	chr20	47897021	+	.	43	0	7043046_1	87.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7043046_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:47895263(+)-20:47897021(-)__20_47873001_47898001D;SPAN=1758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:203 GQ:87.1 PL:[87.1, 0.0, 404.0] SR:0 DR:43 LR:-86.95 LO:98.67);ALT=C[chr20:47897021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	54434623	+	chr20	54440617	+	.	66	46	7068164_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AATAAATTTGTGG;MAPQ=60;MATEID=7068164_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_20_54439001_54464001_8C;SPAN=5994;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:66 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:46 DR:66 LR:-260.8 LO:260.8);ALT=G[chr20:54440617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55043829	+	chr20	55049727	+	.	53	0	7069985_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7069985_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:55043829(+)-20:55049727(-)__20_55027001_55052001D;SPAN=5898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:132 GQ:99 PL:[139.4, 0.0, 179.0] SR:0 DR:53 LR:-139.2 LO:139.5);ALT=G[chr20:55049727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	60714967	+	chr20	60718262	+	AGGCCATGCAGACGTTGTCATCCAAAGCACAGATCTTCCGCACTGTTCTTTCATCCTGCAGTTTGGCCACTGACTTCTTCTCCACACCAAGAACAACAATGTCTCTTCCTCGAACACCA	91	133	7089945_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGGCCATGCAGACGTTGTCATCCAAAGCACAGATCTTCCGCACTGTTCTTTCATCCTGCAGTTTGGCCACTGACTTCTTCTCCACACCAAGAACAACAATGTCTCTTCCTCGAACACCA;MAPQ=60;MATEID=7089945_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_60711001_60736001_226C;SPAN=3295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:179 DP:153 GQ:48.4 PL:[531.4, 48.4, 0.0] SR:133 DR:91 LR:-531.4 LO:531.4);ALT=A[chr20:60718262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	60716001	+	chr20	60718262	+	.	118	39	7089949_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=7089949_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_20_60711001_60736001_226C;SPAN=2261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:142 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:39 DR:118 LR:-419.2 LO:419.2);ALT=C[chr20:60718262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62596231	+	chr20	62597441	+	.	41	0	7096127_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7096127_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62596231(+)-20:62597441(-)__20_62573001_62598001D;SPAN=1210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:59 GQ:23.6 PL:[119.3, 0.0, 23.6] SR:0 DR:41 LR:-123.0 LO:123.0);ALT=G[chr20:62597441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62612669	+	chr20	62614399	+	.	42	36	7096555_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7096555_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62597501_62622501_283C;SPAN=1730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:113 GQ:99 PL:[167.6, 0.0, 104.9] SR:36 DR:42 LR:-168.2 LO:168.2);ALT=G[chr20:62614399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40383249	+	chr21	40386577	+	.	35	2	7178258_1	95.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=7178258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40376001_40401001_274C;SPAN=3328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:88 GQ:95 PL:[95.0, 0.0, 118.1] SR:2 DR:35 LR:-95.0 LO:95.14);ALT=G[chr21:40386577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	17770350	+	chr22	17779109	+	C	88	83	7208307_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=7208307_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_17762501_17787501_215C;SPAN=8759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:32 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:83 DR:88 LR:-425.8 LO:425.8);ALT=C[chr22:17779109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18057770	+	chr22	18060458	+	.	91	18	7210196_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=ATTCTCCTGCCTCAGCCTCC;MAPQ=60;MATEID=7210196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18032001_18057001_398C;SPAN=2688;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:0 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:18 DR:91 LR:-310.3 LO:310.3);ALT=C[chr22:18060458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18226825	+	chr22	18257142	+	.	55	0	7211033_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7211033_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:18226825(+)-22:18257142(-)__22_18203501_18228501D;SPAN=30317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:66 GQ:4.5 PL:[168.3, 4.5, 0.0] SR:0 DR:55 LR:-174.7 LO:174.7);ALT=G[chr22:18257142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19420131	+	chr22	19422257	+	CTTCTGGGAACTTGGCAGACGCAGCTTAGAGAGACTCACCAGCGAGCGTCATTGTTGTCTTTCTGGGAACTCATTCCCATG	33	28	7216473_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTTCTGGGAACTTGGCAGACGCAGCTTAGAGAGACTCACCAGCGAGCGTCATTGTTGTCTTTCTGGGAACTCATTCCCATG;MAPQ=60;MATEID=7216473_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_19404001_19429001_151C;SPAN=2126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:112 GQ:99 PL:[128.3, 0.0, 141.5] SR:28 DR:33 LR:-128.1 LO:128.2);ALT=G[chr22:19422257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19929420	+	chr22	19948720	+	.	43	21	7218375_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7218375_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19918501_19943501_29C;SPAN=19300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:21 DR:43 LR:-158.4 LO:158.4);ALT=G[chr22:19948720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19948812	+	chr22	19950048	+	.	42	72	7218265_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7218265_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19943001_19968001_172C;SPAN=1236;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:119 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:72 DR:42 LR:-353.2 LO:353.2);ALT=G[chr22:19950048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20105351	+	chr22	20106529	+	.	52	0	7219105_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7219105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:20105351(+)-22:20106529(-)__22_20090001_20115001D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:86 GQ:59.3 PL:[148.4, 0.0, 59.3] SR:0 DR:52 LR:-150.4 LO:150.4);ALT=G[chr22:20106529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20950623	+	chr22	20953840	+	.	54	41	7222288_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7222288_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_20947501_20972501_293C;SPAN=3217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:75 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:41 DR:54 LR:-241.0 LO:241.0);ALT=C[chr22:20953840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24195941	+	chr22	24198506	+	.	44	51	7237519_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=GAAAAAAA;MAPQ=60;MATEID=7237519_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_22_24181501_24206501_422C;SPAN=2565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:72 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:51 DR:44 LR:-237.7 LO:237.7);ALT=A[chr22:24198506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24276436	+	chr22	24279226	+	.	102	97	7238239_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CG;MAPQ=60;MATEID=7238239_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_24255001_24280001_53C;SPAN=2790;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:40 GQ:46 PL:[505.0, 46.0, 0.0] SR:97 DR:102 LR:-505.0 LO:505.0);ALT=G[chr22:24279226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24952039	+	chr22	24953624	+	.	97	14	7240580_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7240580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24941001_24966001_110C;SPAN=1585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:112 GQ:30 PL:[330.0, 30.0, 0.0] SR:14 DR:97 LR:-330.1 LO:330.1);ALT=G[chr22:24953624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24952066	+	chr22	24963945	+	.	54	0	7240581_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7240581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:24952066(+)-22:24963945(-)__22_24941001_24966001D;SPAN=11879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:116 GQ:99 PL:[146.9, 0.0, 133.7] SR:0 DR:54 LR:-146.9 LO:146.9);ALT=G[chr22:24963945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	29195143	+	chr22	29196285	+	.	55	81	7256402_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7256402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_29179501_29204501_262C;SPAN=1142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:162 GQ:99 PL:[286.4, 0.0, 104.9] SR:81 DR:55 LR:-290.7 LO:290.7);ALT=T[chr22:29196285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30163537	+	chr22	30165666	+	.	138	112	7260691_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7260691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30159501_30184501_288C;SPAN=2129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:208 DP:226 GQ:61 PL:[670.0, 61.0, 0.0] SR:112 DR:138 LR:-670.1 LO:670.1);ALT=G[chr22:30165666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36745302	+	chr22	36783850	+	.	51	38	7287002_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=7287002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36774501_36799501_117C;SPAN=38548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:38 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:38 DR:51 LR:-208.0 LO:208.0);ALT=T[chr22:36783850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36920837	+	chr22	36925120	+	.	38	0	7287919_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7287919_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36920837(+)-22:36925120(-)__22_36897001_36922001D;SPAN=4283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:38 LR:-115.5 LO:115.5);ALT=A[chr22:36925120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36921808	+	chr22	36925122	+	.	51	0	7287926_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7287926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36921808(+)-22:36925122(-)__22_36897001_36922001D;SPAN=3314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:51 LR:-158.4 LO:158.4);ALT=C[chr22:36925122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36922181	+	chr22	36925123	+	.	97	17	7287927_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7287927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36897001_36922001_308C;SPAN=2942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:0 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:17 DR:97 LR:-303.7 LO:303.7);ALT=G[chr22:36925123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37143176	+	chr22	37147896	+	.	83	49	7288674_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGTAGCT;MAPQ=60;MATEID=7288674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37117501_37142501_166C;SPAN=4720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:0 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:49 DR:83 LR:-340.0 LO:340.0);ALT=T[chr22:37147896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37415952	+	chr22	37420230	+	.	31	0	7289659_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7289659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37415952(+)-22:37420230(-)__22_37411501_37436501D;SPAN=4278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:93 GQ:77.3 PL:[77.3, 0.0, 146.6] SR:0 DR:31 LR:-77.14 LO:78.38);ALT=G[chr22:37420230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37628082	+	chr22	37640178	+	.	53	0	7290446_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7290446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37628082(+)-22:37640178(-)__22_37632001_37657001D;SPAN=12096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:112 GQ:99 PL:[144.8, 0.0, 125.0] SR:0 DR:53 LR:-144.7 LO:144.7);ALT=T[chr22:37640178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37637699	+	chr22	37640153	+	.	81	58	7290464_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=7290464_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_22_37632001_37657001_39C;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:157 GQ:99 PL:[277.7, 0.0, 102.8] SR:58 DR:81 LR:-282.0 LO:282.0);ALT=C[chr22:37640153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37967989	+	chr22	37975965	+	.	73	0	7292182_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7292182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37967989(+)-22:37975965(-)__22_37975001_38000001D;SPAN=7976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:98 GQ:23 PL:[214.4, 0.0, 23.0] SR:0 DR:73 LR:-223.4 LO:223.4);ALT=C[chr22:37975965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38245490	+	chr22	38247284	+	CGGCTTATGACCCCTACGCTTATCCCAGCGACTATGATATGCACA	126	42	7293202_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CGGCTTATGACCCCTACGCTTATCCCAGCGACTATGATATGCACA;MAPQ=60;MATEID=7293202_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_38244501_38269501_180C;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:196 DP:191 GQ:52.9 PL:[580.9, 52.9, 0.0] SR:42 DR:126 LR:-580.9 LO:580.9);ALT=G[chr22:38247284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38349814	+	chr22	38355351	+	TTTTGATGGCGACGACTTTGATGATGTGGAGGAGGATGAAGGGCTAGATGACTTGGAGAATGCCGAAG	41	42	7293627_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TTTTGATGGCGACGACTTTGATGATGTGGAGGAGGATGAAGGGCTAGATGACTTGGAGAATGCCGAAG;MAPQ=60;MATEID=7293627_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_38342501_38367501_184C;SPAN=5537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:122 GQ:99 PL:[175.1, 0.0, 119.0] SR:42 DR:41 LR:-175.4 LO:175.4);ALT=A[chr22:38355351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39294108	+	chr22	39298685	+	.	90	81	7297678_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAAA;MAPQ=60;MATEID=7297678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39298001_39323001_190C;SPAN=4577;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:20 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:81 DR:90 LR:-399.4 LO:399.4);ALT=A[chr22:39298685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39746114	+	chr22	39770320	+	.	41	12	7299716_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7299716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39763501_39788501_68C;SPAN=24206;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:65 GQ:25.4 PL:[131.0, 0.0, 25.4] SR:12 DR:41 LR:-134.8 LO:134.8);ALT=G[chr22:39770320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39925974	+	chr22	39928691	+	.	62	0	7300478_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7300478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39925974(+)-22:39928691(-)__22_39910501_39935501D;SPAN=2717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:108 GQ:86.3 PL:[175.4, 0.0, 86.3] SR:0 DR:62 LR:-177.0 LO:177.0);ALT=A[chr22:39928691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347483	+	chr22	41363802	+	.	34	0	7306462_1	98.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7306462_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347483(+)-22:41363802(-)__22_41331501_41356501D;SPAN=16319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:50 GQ:22.7 PL:[98.6, 0.0, 22.7] SR:0 DR:34 LR:-101.4 LO:101.4);ALT=T[chr22:41363802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347803	+	chr22	41349555	+	.	44	0	7306464_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7306464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347803(+)-22:41349555(-)__22_41331501_41356501D;SPAN=1752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:127 GQ:99 PL:[110.9, 0.0, 196.7] SR:0 DR:44 LR:-110.8 LO:112.2);ALT=G[chr22:41349555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347899	+	chr22	41360048	+	.	59	0	7306466_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7306466_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347899(+)-22:41360048(-)__22_41331501_41356501D;SPAN=12149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:69 GQ:8.7 PL:[184.8, 8.7, 0.0] SR:0 DR:59 LR:-189.4 LO:189.4);ALT=C[chr22:41360048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42071233	+	chr22	42084796	+	.	61	0	7310094_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7310094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42071233(+)-22:42084796(-)__22_42066501_42091501D;SPAN=13563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:152 GQ:99 PL:[160.4, 0.0, 206.6] SR:0 DR:61 LR:-160.2 LO:160.5);ALT=T[chr22:42084796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42076369	+	chr22	42084798	+	.	36	8	7310127_1	72.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7310127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42066501_42091501_397C;SPAN=8429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:170 GQ:72.8 PL:[72.8, 0.0, 340.1] SR:8 DR:36 LR:-72.78 LO:82.6);ALT=C[chr22:42084798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42475958	+	chr22	42477929	+	.	40	84	7311743_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=7311743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42458501_42483501_304C;SPAN=1971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:104 DP:159 GQ:85.7 PL:[300.2, 0.0, 85.7] SR:84 DR:40 LR:-306.8 LO:306.8);ALT=A[chr22:42477929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43027507	+	chr22	43045300	+	.	41	0	7313859_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7313859_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43027507(+)-22:43045300(-)__22_43022001_43047001D;SPAN=17793;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:54 GQ:8.6 PL:[120.8, 0.0, 8.6] SR:0 DR:41 LR:-126.2 LO:126.2);ALT=A[chr22:43045300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43032853	+	chr22	43045301	+	.	50	7	7313877_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7313877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43022001_43047001_196C;SPAN=12448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:85 GQ:56.3 PL:[148.7, 0.0, 56.3] SR:7 DR:50 LR:-150.8 LO:150.8);ALT=C[chr22:43045301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43547662	+	chr22	43557055	+	.	45	0	7316166_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7316166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43547662(+)-22:43557055(-)__22_43536501_43561501D;SPAN=9393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:149 GQ:99 PL:[108.2, 0.0, 253.4] SR:0 DR:45 LR:-108.2 LO:111.4);ALT=G[chr22:43557055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43547662	+	chr22	43555214	+	.	140	0	7316165_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7316165_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43547662(+)-22:43555214(-)__22_43536501_43561501D;SPAN=7552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:186 GQ:38.8 PL:[411.8, 0.0, 38.8] SR:0 DR:140 LR:-429.7 LO:429.7);ALT=G[chr22:43555214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44420331	+	chr22	44489807	+	.	39	22	7319655_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7319655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44467501_44492501_36C;SPAN=69476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:67 GQ:51.2 PL:[110.6, 0.0, 51.2] SR:22 DR:39 LR:-111.7 LO:111.7);ALT=G[chr22:44489807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	45049189	+	chr22	45048157	+	.	31	0	7322063_1	69.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7322063_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:45048157(-)-22:45049189(+)__22_45031001_45056001D;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:123 GQ:69.2 PL:[69.2, 0.0, 227.6] SR:0 DR:31 LR:-69.01 LO:73.83);ALT=]chr22:45049189]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	50624455	+	chr22	50631472	+	.	37	0	7342490_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7342490_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:50624455(+)-22:50631472(-)__22_50617001_50642001D;SPAN=7017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:60 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:0 DR:37 LR:-107.5 LO:107.5);ALT=C[chr22:50631472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	15756524	+	chrX	15768091	+	.	37	0	7370718_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7370718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:15756524(+)-23:15768091(-)__23_15753501_15778501D;SPAN=11567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:68 GQ:60.8 PL:[103.7, 0.0, 60.8] SR:0 DR:37 LR:-104.3 LO:104.3);ALT=A[chrX:15768091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19854401	+	chrX	19905425	+	.	41	67	7377322_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7377322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19894001_19919001_262C;SPAN=51024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:28 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:67 DR:41 LR:-250.9 LO:250.9);ALT=C[chrX:19905425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47441921	+	chrX	47444333	+	.	82	0	7415622_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7415622_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47441921(+)-23:47444333(-)__23_47432001_47457001D;SPAN=2412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:116 GQ:41.3 PL:[239.3, 0.0, 41.3] SR:0 DR:82 LR:-247.1 LO:247.1);ALT=G[chrX:47444333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47441924	+	chrX	47444601	+	.	35	0	7415624_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47441924(+)-23:47444601(-)__23_47432001_47457001D;SPAN=2677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:97 GQ:89.3 PL:[89.3, 0.0, 145.4] SR:0 DR:35 LR:-89.26 LO:90.01);ALT=T[chrX:47444601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47487972	+	chrX	47488982	+	.	51	0	7415543_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7415543_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47487972(+)-23:47488982(-)__23_47481001_47506001D;SPAN=1010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:94 GQ:83.6 PL:[143.0, 0.0, 83.6] SR:0 DR:51 LR:-143.7 LO:143.7);ALT=G[chrX:47488982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47517090	+	chrX	47518288	+	.	55	0	7415834_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47517090(+)-23:47518288(-)__23_47505501_47530501D;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:97 GQ:79.4 PL:[155.3, 0.0, 79.4] SR:0 DR:55 LR:-156.6 LO:156.6);ALT=G[chrX:47518288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48380297	+	chrX	48382086	+	.	60	3	7417402_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=7417402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48363001_48388001_60C;SPAN=1789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:74 GQ:0 PL:[178.2, 0.0, 0.0] SR:3 DR:60 LR:-188.7 LO:188.7);ALT=T[chrX:48382086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49028443	+	chrX	49029476	+	.	102	154	7418806_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=7418806_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TATTAT;SCTG=c_23_49024501_49049501_63C;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:225 DP:175 GQ:60.5 PL:[525.3, 60.5, 0.0] SR:154 DR:102 LR:-525.4 LO:525.4);ALT=T[chrX:49029476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	51279677	+	chrX	51966036	-	.	32	0	7423313_1	86.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=7423313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:51279677(+)-23:51966036(+)__23_51964501_51989501D;SPAN=686359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:72 GQ:86.3 PL:[86.3, 0.0, 86.3] SR:0 DR:32 LR:-86.13 LO:86.13);ALT=C]chrX:51966036];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	53459404	+	chrX	53461264	+	.	44	0	7425680_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7425680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:53459404(+)-23:53461264(-)__23_53459001_53484001D;SPAN=1860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:76 GQ:58.7 PL:[124.7, 0.0, 58.7] SR:0 DR:44 LR:-125.9 LO:125.9);ALT=C[chrX:53461264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70129274	-	chrX	70140010	+	.	42	0	7444682_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7444682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:70129274(-)-23:70140010(-)__23_70119001_70144001D;SPAN=10736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:39 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=[chrX:70140010[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	70503594	+	chrX	70510476	+	.	41	0	7445461_1	99.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=7445461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:70503594(+)-23:70510476(-)__23_70486501_70511501D;SPAN=6882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:41 LR:-132.0 LO:132.0);ALT=T[chrX:70510476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77121417	+	chrX	77123867	+	.	70	27	7455196_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTCACGCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=60;MATEID=7455196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_77101501_77126501_63C;SPAN=2450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:20 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:27 DR:70 LR:-267.4 LO:267.4);ALT=C[chrX:77123867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77155090	+	chrX	77158137	+	.	80	45	7455258_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AAG;MAPQ=60;MATEID=7455258_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_77150501_77175501_297C;SPAN=3047;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:86 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:45 DR:80 LR:-333.4 LO:333.4);ALT=G[chrX:77158137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77359865	+	chrX	77369238	+	.	45	0	7455545_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7455545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:77359865(+)-23:77369238(-)__23_77346501_77371501D;SPAN=9373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:97 GQ:99 PL:[122.3, 0.0, 112.4] SR:0 DR:45 LR:-122.3 LO:122.3);ALT=G[chrX:77369238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	106957980	+	chrX	106959920	+	ATGGCCTGTTCGATCTTGTTGTCTATGGCCACCACGCTGGCTCCGGAGGCA	65	165	7492976_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATGGCCTGTTCGATCTTGTTGTCTATGGCCACCACGCTGGCTCCGGAGGCA;MAPQ=60;MATEID=7492976_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_106942501_106967501_92C;SPAN=1940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:198 DP:123 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:165 DR:65 LR:-587.5 LO:587.5);ALT=C[chrX:106959920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	133594368	+	chrX	133607388	+	.	50	11	7530656_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7530656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_133574001_133599001_157C;SPAN=13020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:30 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:11 DR:50 LR:-151.8 LO:151.8);ALT=G[chrX:133607388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	133594407	+	chrX	133609208	+	.	77	0	7530657_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7530657_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:133594407(+)-23:133609208(-)__23_133574001_133599001D;SPAN=14801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:17 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:0 DR:77 LR:-227.8 LO:227.8);ALT=C[chrX:133609208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	148735758	+	chrX	148830979	-	.	41	0	7552645_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7552645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:148735758(+)-23:148830979(+)__23_148813001_148838001D;SPAN=95221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:24 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=T]chrX:148830979];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	150293942	+	chrX	150295716	+	.	39	34	7554681_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAA;MAPQ=60;MATEID=7554681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_150283001_150308001_38C;SPAN=1774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:15 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:34 DR:39 LR:-174.9 LO:174.9);ALT=A[chrX:150295716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	150565833	+	chrX	150572100	+	.	35	19	7555028_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7555028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_150552501_150577501_214C;SPAN=6267;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:46 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:19 DR:35 LR:-148.5 LO:148.5);ALT=G[chrX:150572100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
