chr12	42555568	+	chr12	42631400	+	.	0	9	5164396_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5164396_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_42532001_42557001_244C;SPAN=75832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:9 DR:0 LR:-19.41 LO:21.15);ALT=C[chr12:42631400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	42697871	+	chr12	42700094	+	.	16	6	5165043_1	53.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CCTCGGCCTCCCAAAGTGCTGGGATTGCAGGCATGAGCC;MAPQ=60;MATEID=5165043_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_42679001_42704001_313C;SPAN=2223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:61 GQ:53 PL:[53.0, 0.0, 92.6] SR:6 DR:16 LR:-52.8 LO:53.46);ALT=C[chr12:42700094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	42717928	+	chr12	42719815	+	.	17	0	5165271_1	29.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=5165271_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:42717928(+)-12:42719815(-)__12_42703501_42728501D;SPAN=1887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:100 GQ:29 PL:[29.0, 0.0, 213.8] SR:0 DR:17 LR:-29.02 LO:37.19);ALT=T[chr12:42719815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	42720070	+	chr12	42729683	+	.	8	0	5165276_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5165276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:42720070(+)-12:42729683(-)__12_42703501_42728501D;SPAN=9613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=C[chr12:42729683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	42729777	+	chr12	42748963	+	.	0	9	5164811_1	6.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5164811_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_42728001_42753001_48C;SPAN=19186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:9 DR:0 LR:-6.139 LO:17.59);ALT=G[chr12:42748963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
