chr7	121878660	+	chr7	121924954	-	.	15	0	3558604_1	28.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3558604_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:121878660(+)-7:121924954(+)__7_121912001_121937001D;SPAN=46294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:77 GQ:28.7 PL:[28.7, 0.0, 157.4] SR:0 DR:15 LR:-28.65 LO:33.8);ALT=A]chr7:121924954];VARTYPE=BND:INV-hh;JOINTYPE=hh
