chr6	122768152	+	chr6	122772809	+	GAATAAAATACACACAACAAAAAGAGAATTAGTCCTATAATTCCTTGAGCATGCCACCACTGGACTGACTGCCCTTCCTTTGGGACAGTGCTTGTTGTATTGTAGCCAATTATGCTTAGTAGACTTGGGTTGCAATTTGTTT	3	8	3010067_1	22.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GAATAAAATACACACAACAAAAAGAGAATTAGTCCTATAATTCCTTGAGCATGCCACCACTGGACTGACTGCCCTTCCTTTGGGACAGTGCTTGTTGTATTGTAGCCAATTATGCTTAGTAGACTTGGGTTGCAATTTGTTT;MAPQ=60;MATEID=3010067_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_122745001_122770001_107C;SPAN=4657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:8 DR:3 LR:-22.44 LO:23.91);ALT=G[chr6:122772809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	122768413	+	chr6	122772809	+	.	2	5	3009964_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=3009964_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_6_122769501_122794501_279C;SPAN=4396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:34 GQ:10.7 PL:[10.7, 0.0, 70.1] SR:5 DR:2 LR:-10.59 LO:13.23);ALT=G[chr6:122772809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	122779827	+	chr6	122792844	+	.	15	6	3009988_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3009988_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_122769501_122794501_20C;SPAN=13017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:87 GQ:32.6 PL:[32.6, 0.0, 177.8] SR:6 DR:15 LR:-32.55 LO:38.33);ALT=C[chr6:122792844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	122931681	+	chr6	122954427	+	.	6	7	3010361_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3010361_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_122941001_122966001_194C;SPAN=22746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:7 DR:6 LR:-19.68 LO:21.27);ALT=G[chr6:122954427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	123039108	+	chr6	123046271	+	.	11	10	3010660_1	49.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3010660_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_123014501_123039501_96C;SPAN=7163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:36 GQ:36.5 PL:[49.7, 0.0, 36.5] SR:10 DR:11 LR:-49.75 LO:49.75);ALT=G[chr6:123046271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
