chr1	36733250	+	chr1	36734642	-	TTT	64	86	185156_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TTT;MAPQ=60;MATEID=185156_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36725501_36750501_65C;SPAN=1392;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:143 DP:95 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:86 DR:64 LR:-422.5 LO:422.5);ALT=A]chr1:36734642];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	36873709	-	chr1	36874937	+	.	8	0	186113_1	1.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=186113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36873709(-)-1:36874937(-)__1_36872501_36897501D;SPAN=1228;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=[chr1:36874937[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	37424238	+	chr1	37425749	+	.	69	27	188802_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CCTGTGTGCCCTGTGAGCCTGTGTGCCCTGTGA;MAPQ=60;MATEID=188802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_37411501_37436501_318C;SPAN=1511;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:90 DP:95 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:27 DR:69 LR:-280.6 LO:280.6);ALT=A[chr1:37425749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
