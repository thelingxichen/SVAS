chr9	30674468	+	chr7	88091360	+	.	7	26	5028083_1	84.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TTTTTTTTT;MAPQ=18;MATEID=5028083_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_88077501_88102501_60C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:29 DP:40 GQ:12.2 PL:[84.8, 0.0, 12.2] SR:26 DR:7 LR:-88.02 LO:88.02);ALT=]chr9:30674468]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	88518949	+	chr7	88516540	+	CTTTTTTCATATACTTCTTAGCTGCA	0	65	5029752_1	99.0	.	EVDNC=ASSMB;INSERTION=CTTTTTTCATATACTTCTTAGCTGCA;MAPQ=60;MATEID=5029752_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_88494001_88519001_319C;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:65 DP:135 GQ:99 PL:[178.1, 0.0, 148.4] SR:65 DR:0 LR:-178.1 LO:178.1);ALT=]chr7:88518949]T;VARTYPE=BND:DUP-th;JOINTYPE=th
