chr4	14846795	+	chr7	27506295	+	.	91	162	4645411_1	99.0	.	DISC_MAPQ=1;EVDNC=DSCRD;IMPRECISE;MAPQ=0;MATEID=4645411_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GGG;SCTG=c_7_27489001_27514001_16C;SECONDARY;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:192 DP:71 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:162 DR:91 LR:-567.7 LO:567.7);ALT=G[chr7:27506295[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	15706264	+	chr4	15705109	+	.	35	0	2640110_1	91.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2640110_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:15705109(-)-4:15706264(+)__4_15704501_15729501D;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:35 DP:91 GQ:91.1 PL:[91.1, 0.0, 127.4] SR:0 DR:35 LR:-90.88 LO:91.26);ALT=]chr4:15706264]C;VARTYPE=BND:DUP-th;JOINTYPE=th
