chr5	156721866	+	chr5	156723678	+	.	0	23	2622054_1	57.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2622054_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_156702001_156727001_47C;SPAN=1812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:68 GQ:57.5 PL:[57.5, 0.0, 107.0] SR:23 DR:0 LR:-57.5 LO:58.33);ALT=C[chr5:156723678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	157158641	+	chr5	157159875	+	.	0	15	2622721_1	31.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=2622721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_157143001_157168001_25C;SPAN=1234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:66 GQ:31.7 PL:[31.7, 0.0, 127.4] SR:15 DR:0 LR:-31.63 LO:34.94);ALT=T[chr5:157159875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	157244555	+	chr5	157285938	+	.	20	17	2623027_1	82.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=2623027_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_157265501_157290501_4C;SPAN=41383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:33 GQ:2.1 PL:[82.5, 2.1, 0.0] SR:17 DR:20 LR:-85.19 LO:85.19);ALT=G[chr5:157285938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
