chr8	24151708	+	chr8	24157484	+	.	7	4	3783403_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=3783403_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_24132501_24157501_136C;SPAN=5776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:98 GQ:3.3 PL:[0.0, 3.3, 244.2] SR:4 DR:7 LR:3.444 LO:12.5);ALT=G[chr8:24157484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	25066685	+	chr8	25070653	+	.	63	42	3786017_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGCTCAG;MAPQ=60;MATEID=3786017_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_25063501_25088501_45C;SPAN=3968;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:76 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:42 DR:63 LR:-257.5 LO:257.5);ALT=G[chr8:25070653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
