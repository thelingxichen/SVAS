chr8	113795705	+	chr13	39943737	-	.	6	7	4028420_1	28.0	.	DISC_MAPQ=9;EVDNC=ASDIS;HOMSEQ=TTCCTTCCTTCCTTCCTTCCTTCCTTCCTTCCT;MAPQ=19;MATEID=4028420_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_113778001_113803001_343C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:29 GQ:28.4 PL:[28.4, 0.0, 41.6] SR:7 DR:6 LR:-28.45 LO:28.6);ALT=A]chr13:39943737];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	129939978	+	chr11	129979322	+	.	53	37	5050273_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5050273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_129972501_129997501_227C;SPAN=39344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:55 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:37 DR:53 LR:-211.3 LO:211.3);ALT=G[chr11:129979322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	129979497	+	chr11	129990600	+	ATGTATCCAGAGCTACAGATCACAAATGTGATGGAGGCAAACCAGCGGGTTAGTATTGACAACTGGTGCCGGAGGGACAAAAAGCAATGCAAGAGTCGCTTTGTTACACCTTTCAAGTGTCTC	4	64	5050288_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGTATCCAGAGCTACAGATCACAAATGTGATGGAGGCAAACCAGCGGGTTAGTATTGACAACTGGTGCCGGAGGGACAAAAAGCAATGCAAGAGTCGCTTTGTTACACCTTTCAAGTGTCTC;MAPQ=60;MATEID=5050288_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_129972501_129997501_60C;SPAN=11103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:88 GQ:22.4 PL:[190.7, 0.0, 22.4] SR:64 DR:4 LR:-198.4 LO:198.4);ALT=G[chr11:129990600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	129980556	+	chr11	129990600	+	.	5	45	5050290_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5050290_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_11_129972501_129997501_60C;SPAN=10044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:105 GQ:99 PL:[133.4, 0.0, 120.2] SR:45 DR:5 LR:-133.3 LO:133.3);ALT=G[chr11:129990600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	129980556	+	chr11	129991507	+	TGGGTGAATTTGTAAGTGATGTCCTGCTAGTTCCAGAAAAGTGCCAGTTTTTCCACAAAGAGCGGATGGAGGTGTGTGAGAATCACCAGCACTGGCACACGGTAGTCAAAG	18	118	5050291_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TGGGTGAATTTGTAAGTGATGTCCTGCTAGTTCCAGAAAAGTGCCAGTTTTTCCACAAAGAGCGGATGGAGGTGTGTGAGAATCACCAGCACTGGCACACGGTAGTCAAAG;MAPQ=60;MATEID=5050291_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_129972501_129997501_191C;SPAN=10951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:109 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:118 DR:18 LR:-373.0 LO:373.0);ALT=G[chr11:129991507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130003623	+	chr11	130005457	+	.	2	4	5050370_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5050370_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_129997001_130022001_280C;SPAN=1834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:81 GQ:1.8 PL:[0.0, 1.8, 198.0] SR:4 DR:2 LR:2.139 LO:10.82);ALT=G[chr11:130005457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130005611	+	chr11	130010291	+	.	6	6	5050373_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=5050373_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_129997001_130022001_326C;SPAN=4680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:6 DR:6 LR:-4.292 LO:19.12);ALT=G[chr11:130010291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130005611	+	chr11	130011392	+	ATCTGGAGTGGGAGAGCAGGATGGGGGACTGATCGGTGCCGAAGAGAAAGTGATTAACAGTAAGAATAAAGTGGATGAAAACAT	0	12	5050374_1	18.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=ATCTGGAGTGGGAGAGCAGGATGGGGGACTGATCGGTGCCGAAGAGAAAGTGATTAACAGTAAGAATAAAGTGGATGAAAACAT;MAPQ=60;MATEID=5050374_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_129997001_130022001_326C;SPAN=5781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:12 DR:0 LR:-18.21 LO:25.61);ALT=G[chr11:130011392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130010380	+	chr11	130011392	+	.	2	10	5050384_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=5050384_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_129997001_130022001_326C;SPAN=1012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:81 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:2 LR:-11.07 LO:20.36);ALT=T[chr11:130011392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130011971	+	chr11	130013240	+	.	11	11	5050393_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5050393_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_129997001_130022001_51C;SPAN=1269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:92 GQ:31.4 PL:[31.4, 0.0, 189.8] SR:11 DR:11 LR:-31.19 LO:37.87);ALT=T[chr11:130013240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	130184499	+	chr11	130193784	+	.	2	2	5051033_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=7;MATEID=5051033_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_130168501_130193501_20C;SPAN=9285;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:30 GQ:5 PL:[5.0, 0.0, 67.7] SR:2 DR:2 LR:-5.076 LO:8.289);ALT=G[chr11:130193784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	131126739	+	chr11	130625844	+	.	13	0	5053428_1	37.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=5053428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:130625844(-)-11:131126739(+)__11_131124001_131149001D;SPAN=500895;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:21 GQ:11 PL:[37.4, 0.0, 11.0] SR:0 DR:13 LR:-37.82 LO:37.82);ALT=]chr11:131126739]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	131930304	+	chr11	131924268	+	CT	68	50	5055148_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CT;MAPQ=60;MATEID=5055148_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_131908001_131933001_347C;SPAN=6036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:82 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:50 DR:68 LR:-310.3 LO:310.3);ALT=]chr11:131930304]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	132305095	-	chr11	132306477	+	.	9	0	5055836_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5055836_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:132305095(-)-11:132306477(-)__11_132300001_132325001D;SPAN=1382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:0 DR:9 LR:-9.119 LO:18.15);ALT=[chr11:132306477[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	132496166	+	chr13	40801815	+	.	2	3	5056329_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCAC;MAPQ=60;MATEID=5056329_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_132496001_132521001_241C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:50 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:3 DR:2 LR:0.3422 LO:7.35);ALT=C[chr13:40801815[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr13	36910015	+	chr13	36920388	+	.	12	0	5456847_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5456847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:36910015(+)-13:36920388(-)__13_36897001_36922001D;SPAN=10373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:0 DR:12 LR:-17.4 LO:25.39);ALT=T[chr13:36920388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37007359	+	chr13	37011764	+	.	3	5	5457069_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5457069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_36995001_37020001_39C;SPAN=4405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:5 DR:3 LR:1.055 LO:10.95);ALT=G[chr13:37011764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37546173	+	chr13	37559764	+	.	2	4	5458702_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5458702_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_37534001_37559001_269C;SPAN=13591;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:37 GQ:3.2 PL:[3.2, 0.0, 85.7] SR:4 DR:2 LR:-3.18 LO:7.9);ALT=T[chr13:37559764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37567812	+	chr13	37569562	+	TCTCTTCTCTAGATAGCTCAGAGCTTCATCCATCATCACAGGCA	0	24	5458624_1	52.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TCTCTTCTCTAGATAGCTCAGAGCTTCATCCATCATCACAGGCA;MAPQ=60;MATEID=5458624_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_37558501_37583501_242C;SPAN=1750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:101 GQ:52.1 PL:[52.1, 0.0, 190.7] SR:24 DR:0 LR:-51.86 LO:56.45);ALT=G[chr13:37569562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37569734	+	chr13	37573372	+	.	38	3	5458632_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5458632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_37558501_37583501_223C;SPAN=3638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:110 GQ:99 PL:[105.5, 0.0, 161.6] SR:3 DR:38 LR:-105.5 LO:106.2);ALT=C[chr13:37573372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37575008	+	chr13	37577070	+	.	10	0	5458644_1	9.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5458644_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:37575008(+)-13:37577070(-)__13_37558501_37583501D;SPAN=2062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:0 DR:10 LR:-9.44 LO:20.03);ALT=A[chr13:37577070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37575009	+	chr13	37580055	+	.	10	0	5458646_1	11.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5458646_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:37575009(+)-13:37580055(-)__13_37558501_37583501D;SPAN=5046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:81 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.07 LO:20.36);ALT=G[chr13:37580055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37577145	+	chr13	37580056	+	AATTTGCAGCACCATCAACAGATGCCCCTGATAAAGGATACGTT	0	22	5458653_1	50.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATTTGCAGCACCATCAACAGATGCCCCTGATAAAGGATACGTT;MAPQ=60;MATEID=5458653_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_37558501_37583501_279C;SPAN=2911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:84 GQ:50 PL:[50.0, 0.0, 152.3] SR:22 DR:0 LR:-49.86 LO:52.83);ALT=G[chr13:37580056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	37621740	+	chr13	37625625	+	TCCACTTGATAGGTATTTCCTTTTAGGAGGTCTCTGTCGGGCACTTTCAATGACATACTCTGCACGATCCAAAGCTAGTTCTAAAGCTTGTTG	0	15	5458886_1	26.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCCACTTGATAGGTATTTCCTTTTAGGAGGTCTCTGTCGGGCACTTTCAATGACATACTCTGCACGATCCAAAGCTAGTTCTAAAGCTTGTTG;MAPQ=60;MATEID=5458886_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_37607501_37632501_356C;SPAN=3885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:15 DR:0 LR:-26.49 LO:33.08);ALT=T[chr13:37625625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	38071943	+	chr13	38085578	+	.	35	30	5459969_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5459969_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_13_38048501_38073501_114C;SPAN=13635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:36 GQ:15 PL:[165.0, 15.0, 0.0] SR:30 DR:35 LR:-165.0 LO:165.0);ALT=T[chr13:38085578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	39057319	+	chr13	39060202	+	.	63	39	5462292_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGAA;MAPQ=60;MATEID=5462292_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_39053001_39078001_160C;SPAN=2883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:20 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:39 DR:63 LR:-247.6 LO:247.6);ALT=A[chr13:39060202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41341170	+	chr13	41345120	+	.	12	13	5468330_1	29.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5468330_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_41331501_41356501_366C;SPAN=3950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:100 GQ:29 PL:[29.0, 0.0, 213.8] SR:13 DR:12 LR:-29.02 LO:37.19);ALT=C[chr13:41345120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41515907	+	chr13	41516916	+	.	8	0	5468948_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5468948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:41515907(+)-13:41516916(-)__13_41503001_41528001D;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:112 GQ:3.6 PL:[0.0, 3.6, 277.2] SR:0 DR:8 LR:3.936 LO:14.29);ALT=C[chr13:41516916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41517281	+	chr13	41523941	+	CTTTCCATCTTTGTTTTTCTTCTTCACAGATATATTTGGCGTAGTGGCTGGGGAATCTGGTCGTGGTGGTTTAGTTTTTCTT	7	18	5468952_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTTTCCATCTTTGTTTTTCTTCTTCACAGATATATTTGGCGTAGTGGCTGGGGAATCTGGTCGTGGTGGTTTAGTTTTTCTT;MAPQ=60;MATEID=5468952_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_41503001_41528001_236C;SPAN=6660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:88 GQ:48.8 PL:[48.8, 0.0, 164.3] SR:18 DR:7 LR:-48.78 LO:52.31);ALT=C[chr13:41523941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41524109	+	chr13	41525465	+	.	0	58	5468966_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5468966_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_41503001_41528001_78C;SPAN=1356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:106 GQ:93.5 PL:[162.8, 0.0, 93.5] SR:58 DR:0 LR:-163.7 LO:163.7);ALT=T[chr13:41525465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41525575	+	chr13	41532972	+	.	0	29	5468968_1	81.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5468968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_41503001_41528001_15C;SPAN=7397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:52 GQ:42.2 PL:[81.8, 0.0, 42.2] SR:29 DR:0 LR:-82.23 LO:82.23);ALT=G[chr13:41532972[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41533155	+	chr13	41556119	+	.	23	34	5468992_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=5468992_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_41552001_41577001_96C;SPAN=22964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:51 GQ:3.6 PL:[128.7, 3.6, 0.0] SR:34 DR:23 LR:-132.8 LO:132.8);ALT=G[chr13:41556119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41556420	+	chr13	41593363	+	.	74	8	5469132_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5469132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_41576501_41601501_28C;SPAN=36943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:47 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:8 DR:74 LR:-221.2 LO:221.2);ALT=T[chr13:41593363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	41574761	+	chr13	41593364	+	.	13	4	5469053_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5469053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_41552001_41577001_181C;SPAN=18603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:56 GQ:34.4 PL:[34.4, 0.0, 100.4] SR:4 DR:13 LR:-34.34 LO:36.19);ALT=T[chr13:41593364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	42041103	+	chr13	42044613	+	.	15	0	5470889_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5470889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:42041103(+)-13:42044613(-)__13_42042001_42067001D;SPAN=3510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:52 GQ:35.6 PL:[35.6, 0.0, 88.4] SR:0 DR:15 LR:-35.43 LO:36.77);ALT=T[chr13:42044613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	42042977	+	chr13	42044614	+	.	4	7	5470891_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTA;MAPQ=60;MATEID=5470891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_42042001_42067001_106C;SPAN=1637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:96 GQ:7.1 PL:[7.1, 0.0, 224.9] SR:7 DR:4 LR:-7.001 LO:19.58);ALT=A[chr13:42044614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	42949866	+	chr13	42947370	+	.	9	28	5473084_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5473084_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_42948501_42973501_71C;SPAN=2496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:29 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:28 DR:9 LR:-92.42 LO:92.42);ALT=]chr13:42949866]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	42947426	+	chr13	42949870	+	GAAAATGAGG	14	23	5473085_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;INSERTION=GAAAATGAGG;MAPQ=60;MATEID=5473085_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_13_42948501_42973501_301C;SPAN=2444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:23 DR:14 LR:-89.12 LO:89.12);ALT=T[chr13:42949870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43539809	+	chr13	43541448	+	.	99	58	5474803_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAAAATCAGCTGGAG;MAPQ=60;MATEID=5474803_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_43536501_43561501_178C;SPAN=1639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:44 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:58 DR:99 LR:-382.9 LO:382.9);ALT=G[chr13:43541448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43597833	+	chr13	43652747	+	.	20	0	5475010_1	54.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5475010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:43597833(+)-13:43652747(-)__13_43634501_43659501D;SPAN=54914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:44 GQ:50.9 PL:[54.2, 0.0, 50.9] SR:0 DR:20 LR:-54.1 LO:54.1);ALT=C[chr13:43652747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43597840	+	chr13	43643059	+	.	47	0	5475011_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5475011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:43597840(+)-13:43643059(-)__13_43634501_43659501D;SPAN=45219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=G[chr13:43643059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43597872	+	chr13	43639821	+	.	24	28	5475012_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5475012_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_43634501_43659501_189C;SPAN=41949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:40 GQ:4.2 PL:[105.6, 4.2, 0.0] SR:28 DR:24 LR:-108.9 LO:108.9);ALT=T[chr13:43639821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43643139	+	chr13	43652748	+	.	0	46	5475034_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5475034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_43634501_43659501_209C;SPAN=9609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:92 GQ:94.1 PL:[127.1, 0.0, 94.1] SR:46 DR:0 LR:-127.1 LO:127.1);ALT=T[chr13:43652748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	43652824	+	chr13	43681312	+	CCCATCTGCTGGCAAGGCTAAGATTAGAACAGCTCATAGGAGAGTCATGATTTTGAATCACCCAGATAA	0	62	5475053_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=CCCATCTGCTGGCAAGGCTAAGATTAGAACAGCTCATAGGAGAGTCATGATTTTGAATCACCCAGATAA;MAPQ=60;MATEID=5475053_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_43634501_43659501_5C;SPAN=28488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:56 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:62 DR:0 LR:-181.5 LO:181.5);ALT=G[chr13:43681312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
