chr5	46144219	+	chr5	46145991	+	GTGAAAAA	43	27	2466655_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GTGAAAAA;MAPQ=60;MATEID=2466655_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_5_46133501_46158501_50C;SPAN=1772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:18 GQ:15 PL:[165.0, 15.0, 0.0] SR:27 DR:43 LR:-165.0 LO:165.0);ALT=G[chr5:46145991[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
