chr20	57464410	+	chr20	57470667	+	.	0	12	7078919_1	15.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=7078919_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_57452501_57477501_57C;SPAN=6257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:89 GQ:15.5 PL:[15.5, 0.0, 200.3] SR:12 DR:0 LR:-15.5 LO:24.93);ALT=T[chr20:57470667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57466922	+	chr20	57470666	+	.	0	8	7078924_1	11.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7078924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_57452501_57477501_210C;SPAN=3744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:8 DR:0 LR:-11.51 LO:16.91);ALT=T[chr20:57470666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57466969	+	chr20	57478582	+	.	14	0	7079080_1	28.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7079080_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57466969(+)-20:57478582(-)__20_57477001_57502001D;SPAN=11613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:66 GQ:28.4 PL:[28.4, 0.0, 130.7] SR:0 DR:14 LR:-28.33 LO:32.13);ALT=G[chr20:57478582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57470739	+	chr20	57478727	+	TGAGAAGGCAACCAAAGTGCAGGACATCAAAAACAACCTGAAAGAGGCGATTGAA	3	19	7079083_1	54.0	.	DISC_MAPQ=18;EVDNC=TSI_G;INSERTION=TGAGAAGGCAACCAAAGTGCAGGACATCAAAAACAACCTGAAAGAGGCGATTGAA;MAPQ=60;MATEID=7079083_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_57477001_57502001_230C;SPAN=7988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:67 GQ:54.5 PL:[54.5, 0.0, 107.3] SR:19 DR:3 LR:-54.47 LO:55.44);ALT=A[chr20:57478727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57478847	+	chr20	57480438	+	.	14	15	7079089_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=7079089_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_20_57477001_57502001_168C;SPAN=1591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:117 GQ:37.7 PL:[37.7, 0.0, 245.6] SR:15 DR:14 LR:-37.62 LO:46.49);ALT=G[chr20:57480438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57478891	+	chr20	57484216	+	.	10	0	7079091_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7079091_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57478891(+)-20:57484216(-)__20_57477001_57502001D;SPAN=5325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:134 GQ:3 PL:[0.0, 3.0, 330.0] SR:0 DR:10 LR:3.294 LO:18.06);ALT=A[chr20:57484216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57480535	+	chr20	57484401	+	CTTCCTGGACAAGATCGACGTGATCAAGCAGGCTGACTATGTGCCGAGCGA	2	21	7079098_1	41.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TCAGG;INSERTION=CTTCCTGGACAAGATCGACGTGATCAAGCAGGCTGACTATGTGCCGAGCGA;MAPQ=60;MATEID=7079098_2;MATENM=97;NM=0;NUMPARTS=3;SCTG=c_20_57477001_57502001_69C;SPAN=3866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:116 GQ:41.3 PL:[41.3, 0.0, 239.3] SR:21 DR:2 LR:-41.2 LO:49.29);ALT=A[chr20:57484401[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57520581	+	chr20	57522011	-	.	8	0	7079346_1	1.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=7079346_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57520581(+)-20:57522011(+)__20_57501501_57526501D;SPAN=1430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:0 DR:8 LR:-1.212 LO:14.96);ALT=G]chr20:57522011];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr20	57556448	+	chr20	57561144	+	.	11	0	7079391_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7079391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57556448(+)-20:57561144(-)__20_57550501_57575501D;SPAN=4696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:61 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-19.78 LO:24.38);ALT=C[chr20:57561144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57562872	+	chr20	57563967	+	.	2	4	7079416_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7079416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_57550501_57575501_187C;SPAN=1095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:89 GQ:7.5 PL:[0.0, 7.5, 231.0] SR:4 DR:2 LR:7.607 LO:8.395);ALT=G[chr20:57563967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57572809	+	chr20	57576520	+	.	11	17	7079459_1	66.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7079459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_57575001_57600001_424C;SPAN=3711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:46 GQ:43.7 PL:[66.8, 0.0, 43.7] SR:17 DR:11 LR:-66.99 LO:66.99);ALT=C[chr20:57576520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57576700	+	chr20	57581377	+	.	9	6	7079470_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7079470_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_57575001_57600001_405C;SPAN=4677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:98 GQ:16.4 PL:[16.4, 0.0, 221.0] SR:6 DR:9 LR:-16.36 LO:26.91);ALT=C[chr20:57581377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57603917	+	chr20	57607273	+	.	54	0	7079564_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=7079564_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57603917(+)-20:57607273(-)__20_57599501_57624501D;SPAN=3356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:125 GQ:99 PL:[144.5, 0.0, 157.7] SR:0 DR:54 LR:-144.4 LO:144.4);ALT=C[chr20:57607273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57605496	+	chr20	57607273	+	.	72	0	7079567_1	99.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=7079567_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:57605496(+)-20:57607273(-)__20_57599501_57624501D;SPAN=1777;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:142 GQ:99 PL:[199.4, 0.0, 143.3] SR:0 DR:72 LR:-199.6 LO:199.6);ALT=T[chr20:57607273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	57613689	+	chr20	57617754	+	.	25	4	7079591_1	61.0	.	DISC_MAPQ=40;EVDNC=ASDIS;MAPQ=32;MATEID=7079591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_57599501_57624501_331C;SPAN=4065;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:91 GQ:61.4 PL:[61.4, 0.0, 157.1] SR:4 DR:25 LR:-61.17 LO:63.6);ALT=G[chr20:57617754[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
