chr13	30215837	+	chr13	30221845	+	.	30	26	7978746_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAGAACTACTTTTT;MAPQ=60;MATEID=7978746_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_13_30208501_30233501_304C;SPAN=6008;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:80 GQ:44.3 PL:[149.9, 0.0, 44.3] SR:26 DR:30 LR:-153.2 LO:153.2);ALT=T[chr13:30221845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
