chr7	75992937	-	chr7	75994455	+	.	9	0	4978465_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4978465_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:75992937(-)-7:75994455(-)__7_75974501_75999501D;SPAN=1518;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:111 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.3636 LO:16.59);ALT=[chr7:75994455[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
