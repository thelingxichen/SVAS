chr4	25916044	+	chr4	25930774	+	AGAAGGAACAAGCTATAAATCGGGCTGGAATTGTTCAAGAGGATGTGCAGCCACC	12	21	1925776_1	82.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AGAAGGAACAAGCTATAAATCGGGCTGGAATTGTTCAAGAGGATGTGCAGCCACC;MAPQ=60;MATEID=1925776_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_25896501_25921501_47C;SPAN=14730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:31 GQ:4.8 PL:[82.5, 4.8, 0.0] SR:21 DR:12 LR:-82.81 LO:82.81);ALT=A[chr4:25930774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	26290469	+	chr4	26295386	+	.	25	17	1926423_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=1926423_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_4_26288501_26313501_85C;SPAN=4917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:29 GQ:9 PL:[99.0, 9.0, 0.0] SR:17 DR:25 LR:-99.02 LO:99.02);ALT=C[chr4:26295386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
