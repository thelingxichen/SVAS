chr13	23632400	+	chr13	23637302	+	.	31	0	5418686_1	85.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5418686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:23632400(+)-13:23637302(-)__13_23618001_23643001D;SPAN=4902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:64 GQ:68.6 PL:[85.1, 0.0, 68.6] SR:0 DR:31 LR:-85.06 LO:85.06);ALT=G[chr13:23637302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	23935641	-	chr13	23937007	+	.	2	3	5419301_1	0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAGCCACCATG;MAPQ=0;MATEID=5419301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_23912001_23937001_251C;SPAN=1366;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:85 GQ:6.3 PL:[0.0, 6.3, 217.8] SR:3 DR:2 LR:6.524 LO:8.497);ALT=[chr13:23937007[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
