chr1	6086520	+	chr1	6132804	+	.	19	0	17234_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=17234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6086520(+)-1:6132804(-)__1_6125001_6150001D;SPAN=46284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:42 GQ:48.2 PL:[51.5, 0.0, 48.2] SR:0 DR:19 LR:-51.34 LO:51.34);ALT=C[chr1:6132804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6086527	+	chr1	6100573	+	.	25	0	17292_1	73.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=17292_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6086527(+)-1:6100573(-)__1_6100501_6125501D;SPAN=14046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:33 GQ:4.4 PL:[73.7, 0.0, 4.4] SR:0 DR:25 LR:-76.89 LO:76.89);ALT=T[chr1:6100573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6100706	+	chr1	6133792	+	AACCTGGGCAAGTCTGGCCTGCGGGTCTCCTGCCTGGGACTT	2	33	17238_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AACCTGGGCAAGTCTGGCCTGCGGGTCTCCTGCCTGGGACTT;MAPQ=60;MATEID=17238_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_6125001_6150001_71C;SPAN=33086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:33 DR:2 LR:-111.7 LO:111.7);ALT=G[chr1:6133792[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6257850	+	chr1	6259570	+	.	14	0	17642_1	24.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=17642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6257850(+)-1:6259570(-)__1_6247501_6272501D;SPAN=1720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:79 GQ:24.8 PL:[24.8, 0.0, 166.7] SR:0 DR:14 LR:-24.81 LO:30.91);ALT=G[chr1:6259570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	169201745	+	chr1	6259596	+	.	36	0	1779497_1	94.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=1779497_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6259596(-)-3:169201745(+)__3_169197001_169222001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:89 GQ:94.7 PL:[94.7, 0.0, 121.1] SR:0 DR:36 LR:-94.72 LO:94.9);ALT=]chr3:169201745]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	6399650	+	chr1	6409808	+	.	0	12	17994_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=17994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_6394501_6419501_301C;SPAN=10158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:12 DR:0 LR:-19.29 LO:25.9);ALT=C[chr1:6409808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6409927	+	chr1	6453316	+	.	14	10	18031_1	54.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=18031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_6394501_6419501_40C;SPAN=43389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:43 GQ:47.9 PL:[54.5, 0.0, 47.9] SR:10 DR:14 LR:-54.38 LO:54.38);ALT=C[chr1:6453316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6409928	+	chr1	6418885	+	.	12	5	18645_1	33.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=18645_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_6419001_6444001_153C;SPAN=8957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:0 GQ:3 PL:[33.0, 3.0, 0.0] SR:5 DR:12 LR:-33.01 LO:33.01);ALT=T[chr1:6418885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6845635	+	chr1	6880239	+	.	19	15	19365_1	66.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=19365_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_6835501_6860501_135C;SPAN=34604;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:12 GQ:6 PL:[66.0, 6.0, 0.0] SR:15 DR:19 LR:-66.02 LO:66.02);ALT=G[chr1:6880239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6845683	+	chr1	6885148	+	.	47	0	19397_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=19397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6845683(+)-1:6885148(-)__1_6884501_6909501D;SPAN=39465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=G[chr1:6885148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6845683	+	chr1	6931814	+	.	24	0	19367_1	69.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=19367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:6845683(+)-1:6931814(-)__1_6835501_6860501D;SPAN=86131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:3 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=G[chr1:6931814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	6880310	+	chr1	6885150	+	.	2	15	19398_1	44.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=19398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_6884501_6909501_125C;SPAN=4840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:45 GQ:44 PL:[44.0, 0.0, 63.8] SR:15 DR:2 LR:-43.93 LO:44.15);ALT=G[chr1:6885150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	7570071	+	chr1	7571527	+	TCCTGCACATGCTTA	18	13	21249_1	79.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TCCTGCACATGCTTA;MAPQ=60;MATEID=21249_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_1_7570501_7595501_54C;SPAN=1456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:25 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:13 DR:18 LR:-79.22 LO:79.22);ALT=A[chr1:7571527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	7831490	+	chr1	7837217	+	.	14	0	21975_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=21975_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:7831490(+)-1:7837217(-)__1_7815501_7840501D;SPAN=5727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:81 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:0 DR:14 LR:-24.27 LO:30.74);ALT=G[chr1:7837217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	7833573	+	chr1	7837218	+	.	0	12	21983_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=21983_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_7815501_7840501_318C;SPAN=3645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:12 DR:0 LR:-17.67 LO:25.46);ALT=T[chr1:7837218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	7837378	+	chr1	7839685	+	ATGTGGGCAATCGGGATTACTGTTCTGGTTATCTTCATCATCATCATCATC	2	13	21990_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGTGGGCAATCGGGATTACTGTTCTGGTTATCTTCATCATCATCATCATC;MAPQ=60;MATEID=21990_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_7815501_7840501_109C;SPAN=2307;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:79 GQ:21.5 PL:[21.5, 0.0, 170.0] SR:13 DR:2 LR:-21.51 LO:28.24);ALT=G[chr1:7839685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8021854	+	chr1	8025383	+	CTTGTAAACATATAACATAAAAATGGCTTCCAAAAGAGCTCTGGTCATCCTGGCTAAAGGAGCAGAGGAAATGGAGACGGTCATCCCTGTAGATGTCATGAGGCGAGCTGG	61	131	22705_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTTGTAAACATATAACATAAAAATGGCTTCCAAAAGAGCTCTGGTCATCCTGGCTAAAGGAGCAGAGGAAATGGAGACGGTCATCCCTGTAGATGTCATGAGGCGAGCTGG;MAPQ=60;MATEID=22705_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_8011501_8036501_97C;SPAN=3529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:99 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:131 DR:61 LR:-458.8 LO:458.8);ALT=G[chr1:8025383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8022935	+	chr1	8025383	+	.	20	107	22714_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=22714_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_1_8011501_8036501_97C;SPAN=2448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:100 GQ:33 PL:[363.0, 33.0, 0.0] SR:107 DR:20 LR:-363.1 LO:363.1);ALT=G[chr1:8025383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8025486	+	chr1	8030952	+	GACCATATGATGTGGTGGTTCTACCAGGAGGTAATCTGGGCGCACAGAATTTATCTG	2	104	22727_1	99.0	.	DISC_MAPQ=33;EVDNC=TSI_G;HOMSEQ=AGTCTGCTGCTGTGAAGGAGATACTGAAGGAGCAGGAAAACC;INSERTION=GACCATATGATGTGGTGGTTCTACCAGGAGGTAATCTGGGCGCACAGAATTTATCTG;MAPQ=60;MATEID=22727_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_8011501_8036501_240C;SECONDARY;SPAN=5466;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:94 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:104 DR:2 LR:-307.0 LO:307.0);ALT=G[chr1:8030952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8031025	+	chr1	8037710	+	.	0	17	22765_1	45.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=22765_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8036001_8061001_7C;SPAN=6685;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:17 DR:0 LR:-45.01 LO:45.06);ALT=T[chr1:8037710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8037800	+	chr1	8044952	+	.	7	17	22769_1	52.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=22769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8036001_8061001_364C;SPAN=7152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:88 GQ:52.1 PL:[52.1, 0.0, 161.0] SR:17 DR:7 LR:-52.08 LO:55.21);ALT=T[chr1:8044952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8923947	-	chr1	236647585	+	.	26	0	617062_1	71.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=617062_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:8923947(-)-1:236647585(-)__1_236645501_236670501D;SPAN=227723638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:53 GQ:55.1 PL:[71.6, 0.0, 55.1] SR:0 DR:26 LR:-71.55 LO:71.55);ALT=[chr1:236647585[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	8924153	+	chr1	8925344	+	.	32	12	25213_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=9;MATEID=25213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8918001_8943001_29C;SPAN=1191;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:78 GQ:64.7 PL:[124.1, 0.0, 64.7] SR:12 DR:32 LR:-125.1 LO:125.1);ALT=T[chr1:8925344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8926613	+	chr1	8928040	+	.	19	0	25226_1	40.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=25226_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:8926613(+)-1:8928040(-)__1_8918001_8943001D;SPAN=1427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:83 GQ:40.4 PL:[40.4, 0.0, 159.2] SR:0 DR:19 LR:-40.23 LO:44.33);ALT=G[chr1:8928040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8934978	+	chr1	8938639	+	.	122	58	25255_1	99.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=43;MATEID=25255_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_8918001_8943001_205C;SPAN=3661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:108 GQ:36 PL:[396.0, 36.0, 0.0] SR:58 DR:122 LR:-396.1 LO:396.1);ALT=T[chr1:8938639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	8938639	-	chr1	236646440	+	.	163	19	617066_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CTAGCCACTGGGTCTC;MAPQ=60;MATEID=617066_2;MATENM=12;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_1_236645501_236670501_12C;SPAN=227707801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:182 DP:79 GQ:49 PL:[538.0, 49.0, 0.0] SR:19 DR:163 LR:-538.0 LO:538.0);ALT=[chr1:236646440[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	9711885	+	chr1	9751525	+	.	8	0	27959_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=27959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:9711885(+)-1:9751525(-)__1_9702001_9727001D;SPAN=39640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:21 GQ:20.9 PL:[20.9, 0.0, 27.5] SR:0 DR:8 LR:-20.72 LO:20.82);ALT=C[chr1:9751525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9931335	+	chr1	9937962	+	GTTTGATCCCATCTTCCGCAGCATGAGCAGCACTCGGACCTTCTGCTGAATGTACATCTCCTCCGGACTCTTCCCGGGAGCTCCCTCGCGGTTCATCCCCCTGCCTGGCTCTGGGGACT	0	33	28660_1	83.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTGC;INSERTION=GTTTGATCCCATCTTCCGCAGCATGAGCAGCACTCGGACCTTCTGCTGAATGTACATCTCCTCCGGACTCTTCCCGGGAGCTCCCTCGCGGTTCATCCCCCTGCCTGGCTCTGGGGACT;MAPQ=60;MATEID=28660_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_9922501_9947501_174C;SPAN=6627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:93 GQ:83.9 PL:[83.9, 0.0, 140.0] SR:33 DR:0 LR:-83.74 LO:84.56);ALT=G[chr1:9937962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9932150	+	chr1	9937962	+	.	2	20	28664_1	44.0	.	DISC_MAPQ=49;EVDNC=TSI_L;HOMSEQ=CCTGC;MAPQ=60;MATEID=28664_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_9922501_9947501_174C;SPAN=5812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:93 GQ:44.3 PL:[44.3, 0.0, 179.6] SR:20 DR:2 LR:-44.13 LO:48.85);ALT=C[chr1:9937962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9932195	+	chr1	9970151	+	.	14	0	28665_1	38.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=28665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:9932195(+)-1:9970151(-)__1_9922501_9947501D;SPAN=37956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:27 GQ:25.7 PL:[38.9, 0.0, 25.7] SR:0 DR:14 LR:-39.02 LO:39.02);ALT=T[chr1:9970151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9938050	+	chr1	9970152	+	.	0	11	28706_1	29.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=28706_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_9947001_9972001_137C;SPAN=32102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:8 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:11 DR:0 LR:-29.71 LO:29.71);ALT=G[chr1:9970152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9990516	+	chr1	9991948	+	.	0	8	28847_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=28847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_9971501_9996501_174C;SPAN=1432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:8 DR:0 LR:-6.089 LO:15.75);ALT=C[chr1:9991948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9996687	+	chr1	10002682	+	.	0	18	28879_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=28879_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_9996001_10021001_129C;SPAN=5995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:83 GQ:37.1 PL:[37.1, 0.0, 162.5] SR:18 DR:0 LR:-36.93 LO:41.51);ALT=T[chr1:10002682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	9996731	+	chr1	10003335	+	.	8	0	28881_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=28881_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:9996731(+)-1:10003335(-)__1_9996001_10021001D;SPAN=6604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:81 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:0 DR:8 LR:-4.463 LO:15.47);ALT=A[chr1:10003335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	10473309	+	chr1	10477043	+	.	7	6	30790_1	13.0	.	DISC_MAPQ=39;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=30790_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_10461501_10486501_160C;SPAN=3734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:6 DR:7 LR:-13.28 LO:22.64);ALT=G[chr1:10477043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	10477604	+	chr1	10479470	+	.	9	0	30804_1	5.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=30804_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:10477604(+)-1:10479470(-)__1_10461501_10486501D;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:91 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.055 LO:17.41);ALT=T[chr1:10479470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	10529420	+	chr1	10532487	+	.	10	0	30934_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=30934_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:10529420(+)-1:10532487(-)__1_10510501_10535501D;SPAN=3067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:0 DR:10 LR:-12.69 LO:20.72);ALT=A[chr1:10532487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	10914199	+	chr4	130207312	+	.	2	3	31846_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=31846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_10902501_10927501_270C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:39 GQ:2.6 PL:[2.6, 0.0, 91.7] SR:3 DR:2 LR:-2.638 LO:7.803);ALT=A[chr4:130207312[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	11737007	+	chr1	11740410	+	TCTCCAGGAGTGGCTTGACGCAGTGCAGCGTGTCCTGGATATACTGATTCAGCTCCGGGTGGCAGGACAT	0	19	34253_1	40.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TCTCCAGGAGTGGCTTGACGCAGTGCAGCGTGTCCTGGATATACTGATTCAGCTCCGGGTGGCAGGACAT;MAPQ=60;MATEID=34253_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_11735501_11760501_32C;SPAN=3403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:83 GQ:40.4 PL:[40.4, 0.0, 159.2] SR:19 DR:0 LR:-40.23 LO:44.33);ALT=T[chr1:11740410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	11796295	+	chr1	11807496	+	ATTCTCCTAGGTCACTGGCTGCTGACAACCT	36	11	34432_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATTCTCCTAGGTCACTGGCTGCTGACAACCT;MAPQ=60;MATEID=34432_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_11784501_11809501_105C;SPAN=11201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:81 GQ:93.8 PL:[100.4, 0.0, 93.8] SR:11 DR:36 LR:-100.2 LO:100.2);ALT=G[chr1:11807496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	11796327	+	chr1	11808470	+	.	19	0	34433_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=34433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:11796327(+)-1:11808470(-)__1_11784501_11809501D;SPAN=12143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:90 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:0 DR:19 LR:-38.34 LO:43.57);ALT=G[chr1:11808470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	12008125	+	chr1	12009825	+	.	0	7	35181_1	3.0	.	EVDNC=ASSMB;HOMSEQ=TCCAGG;MAPQ=60;MATEID=35181_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_12005001_12030001_18C;SPAN=1700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:7 DR:0 LR:-3.059 LO:13.4);ALT=G[chr1:12009825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	12079644	+	chr1	12081700	+	.	21	0	35579_1	47.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=35579_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:12079644(+)-1:12081700(-)__1_12078501_12103501D;SPAN=2056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:82 GQ:47.3 PL:[47.3, 0.0, 149.6] SR:0 DR:21 LR:-47.11 LO:50.19);ALT=A[chr1:12081700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	12227230	+	chr1	12248849	+	.	0	7	36008_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCAGGTGG;MAPQ=60;MATEID=36008_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_12225501_12250501_190C;SPAN=21619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:76 GQ:2.6 PL:[2.6, 0.0, 180.8] SR:7 DR:0 LR:-2.517 LO:13.31);ALT=G[chr1:12248849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	13774313	-	chr1	13775496	+	.	10	0	40011_1	13.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=40011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:13774313(-)-1:13775496(-)__1_13769001_13794001D;SPAN=1183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:73 GQ:13.4 PL:[13.4, 0.0, 161.9] SR:0 DR:10 LR:-13.23 LO:20.85);ALT=[chr1:13775496[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	207446741	+	chr1	13796643	+	.	3	17	40471_1	66.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AGTAGCTGGGATTA;MAPQ=60;MATEID=40471_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_13793501_13818501_95C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:23 GQ:6 PL:[66.0, 6.0, 0.0] SR:17 DR:3 LR:-64.69 LO:64.69);ALT=]chr2:207446741]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	13796653	+	chr1	32921067	+	.	18	19	40474_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCTGCCTCCCGGGTTCACGCCATTCTCCTGCCTCAGCCTGCTGAGTAGCTGGGA;MAPQ=60;MATEID=40474_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_13793501_13818501_276C;SPAN=19124414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:18 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:19 DR:18 LR:-108.9 LO:108.9);ALT=A[chr1:32921067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	13881560	-	chr21	40685369	+	.	2	33	40265_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;MAPQ=18;MATEID=40265_2;MATENM=0;NM=7;NUMPARTS=2;SCTG=c_1_13867001_13892001_248C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:34 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:33 DR:2 LR:-102.3 LO:102.3);ALT=[chr21:40685369[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	13893343	-	chr1	13894621	+	.	12	0	40138_1	22.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=40138_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:13893343(-)-1:13894621(-)__1_13891501_13916501D;SPAN=1278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:64 GQ:22.4 PL:[22.4, 0.0, 131.3] SR:0 DR:12 LR:-22.27 LO:26.82);ALT=[chr1:13894621[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	15736778	+	chr1	15752367	+	.	10	13	45198_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GTA;MAPQ=60;MATEID=45198_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_15729001_15754001_149C;SPAN=15589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:82 GQ:37.4 PL:[37.4, 0.0, 159.5] SR:13 DR:10 LR:-37.2 LO:41.62);ALT=A[chr1:15752367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	15736778	+	chr1	15753644	+	TGATGCCGGGCGGGACGGCTTCATCGACCTGATGGAGCTAAAACTCATGATGGAGAAACTTGGGGCCCCTCAGACCCACCTGGGCCTGAAAAACATGATCAAGGAGGTGGATGAGGACTTTGACAGCAAGCTGAGCTTCCGGG	3	25	45199_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGATGCCGGGCGGGACGGCTTCATCGACCTGATGGAGCTAAAACTCATGATGGAGAAACTTGGGGCCCCTCAGACCCACCTGGGCCTGAAAAACATGATCAAGGAGGTGGATGAGGACTTTGACAGCAAGCTGAGCTTCCGGG;MAPQ=60;MATEID=45199_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_15729001_15754001_149C;SPAN=16866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:92 GQ:57.8 PL:[57.8, 0.0, 163.4] SR:25 DR:3 LR:-57.6 LO:60.51);ALT=A[chr1:15753644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	15752514	+	chr1	15753644	+	.	7	7	45234_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=45234_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCCTCC;SCTG=c_1_15729001_15754001_149C;SPAN=1130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:6.9 PL:[6.9, 0.0, 155.1] SR:7 DR:7 LR:-6.841 LO:16.53);ALT=G[chr1:15753644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	15753782	+	chr1	15755087	+	.	0	22	45566_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=45566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_15753501_15778501_340C;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:83 GQ:50.3 PL:[50.3, 0.0, 149.3] SR:22 DR:0 LR:-50.14 LO:52.96);ALT=T[chr1:15755087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	15908123	+	chr1	15972909	+	.	8	39	46375_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGGTGGCTCATGCCTGTAATCCCAGCA;MAPQ=60;MATEID=46375_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_15949501_15974501_328C;SPAN=64786;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:58 GQ:14 PL:[126.2, 0.0, 14.0] SR:39 DR:8 LR:-131.4 LO:131.4);ALT=A[chr1:15972909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	15972990	+	chr1	15908144	+	.	18	30	46376_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GGATCACCTGAGGTCAGGAGTTCGAGACCAGCCT;MAPQ=60;MATEID=46376_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_15949501_15974501_365C;SPAN=64846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:49 GQ:6.5 PL:[112.1, 0.0, 6.5] SR:30 DR:18 LR:-117.7 LO:117.7);ALT=]chr1:15972990]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	16154742	-	chr19	39926488	+	.	72	47	47148_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=CCGCTGCAGTCGGTGCAGGTCTTCGGACGCAAG;MAPQ=55;MATEID=47148_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_1_16145501_16170501_79C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:92 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:47 DR:72 LR:-283.9 LO:283.9);ALT=[chr19:39926488[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	16664256	-	chr1	16665360	+	.	8	0	48436_1	6.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=48436_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:16664256(-)-1:16665360(-)__1_16660001_16685001D;SPAN=1104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=[chr1:16665360[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	16693823	+	chr1	16719723	+	.	48	0	48680_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=48680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:16693823(+)-1:16719723(-)__1_16684501_16709501D;SPAN=25900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:49 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:48 LR:-145.2 LO:145.2);ALT=C[chr1:16719723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16767330	+	chr1	16774360	+	.	10	0	48606_1	8.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=48606_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:16767330(+)-1:16774360(-)__1_16758001_16783001D;SPAN=7030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:0 DR:10 LR:-8.627 LO:19.88);ALT=C[chr1:16774360[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16767349	+	chr1	16770125	+	.	14	11	48608_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=48608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_16758001_16783001_132C;SPAN=2776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:11 DR:14 LR:-32.87 LO:40.05);ALT=G[chr1:16770125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	16770228	+	chr1	16774361	+	.	0	9	48616_1	8.0	.	EVDNC=ASSMB;HOMSEQ=TCAGG;MAPQ=60;MATEID=48616_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_16758001_16783001_141C;SPAN=4133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:9 DR:0 LR:-8.306 LO:17.99);ALT=G[chr1:16774361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17051748	-	chr1	234912188	+	GCCCCATCCCGCCGGCTTCTGC	189	57	50768_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;INSERTION=GCCCCATCCCGCCGGCTTCTGC;MAPQ=60;MATEID=50768_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17027501_17052501_901C;SPAN=217860440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:229 DP:175 GQ:61.9 PL:[679.9, 61.9, 0.0] SR:57 DR:189 LR:-680.0 LO:680.0);ALT=[chr1:234912188[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	17345456	+	chr1	17349102	+	.	0	23	53581_1	63.0	.	EVDNC=ASSMB;HOMSEQ=CCTT;MAPQ=60;MATEID=53581_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17346001_17371001_181C;SPAN=3646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:47 GQ:50 PL:[63.2, 0.0, 50.0] SR:23 DR:0 LR:-63.26 LO:63.26);ALT=T[chr1:17349102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17355233	+	chr1	17359554	+	.	3	9	53611_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=53611_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_1_17346001_17371001_292C;SPAN=4321;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:80 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:9 DR:3 LR:-17.94 LO:25.53);ALT=T[chr1:17359554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17355233	+	chr1	17371256	+	TCTCTGCATGATCTTCGGAAGGTCAAAGTAGAGTCAACTTCATTCTTAATCTTGATTAAAGCATCCAATACCATGGGGCCACAT	3	33	53662_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TCTCTGCATGATCTTCGGAAGGTCAAAGTAGAGTCAACTTCATTCTTAATCTTGATTAAAGCATCCAATACCATGGGGCCACAT;MAPQ=60;MATEID=53662_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_17370501_17395501_273C;SPAN=16023;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:42 GQ:4.5 PL:[108.9, 4.5, 0.0] SR:33 DR:3 LR:-111.2 LO:111.2);ALT=T[chr1:17371256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17359690	+	chr1	17380463	+	.	16	0	53665_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=53665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:17359690(+)-1:17380463(-)__1_17370501_17395501D;SPAN=20773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:50 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.27 LO:40.1);ALT=A[chr1:17380463[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17371386	+	chr1	17380442	+	.	34	6	53672_1	95.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=53672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_17370501_17395501_125C;SPAN=9056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:74 GQ:82.4 PL:[95.6, 0.0, 82.4] SR:6 DR:34 LR:-95.52 LO:95.52);ALT=G[chr1:17380442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17634809	+	chr1	17657461	+	.	37	10	54878_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=54878_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_17640001_17665001_160C;SPAN=22652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:53 GQ:5.6 PL:[121.1, 0.0, 5.6] SR:10 DR:37 LR:-126.9 LO:126.9);ALT=G[chr1:17657461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17657646	+	chr1	17660436	+	.	0	14	54933_1	25.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=54933_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_17640001_17665001_59C;SPAN=2790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:78 GQ:25.1 PL:[25.1, 0.0, 163.7] SR:14 DR:0 LR:-25.08 LO:30.99);ALT=T[chr1:17660436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	17676184	+	chr1	17677654	+	.	47	20	54994_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CTGCACTCCAGCCTGGGTGACAGA;MAPQ=60;MATEID=54994_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_17664501_17689501_17C;SPAN=1470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:33 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:20 DR:47 LR:-184.8 LO:184.8);ALT=A[chr1:17677654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	20982273	+	chr1	20987374	+	AATGTCGGAGCTGGCAGCTACCAGCACACTGCCTCCGCCGTCAATAAAGGCACTGATGGTCTCCACGTTGATGTTGCCTCCAAAAT	2	36	64394_1	96.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AATGTCGGAGCTGGCAGCTACCAGCACACTGCCTCCGCCGTCAATAAAGGCACTGATGGTCTCCACGTTGATGTTGCCTCCAAAAT;MAPQ=60;MATEID=64394_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_20972001_20997001_167C;SPAN=5101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:82 GQ:96.8 PL:[96.8, 0.0, 100.1] SR:36 DR:2 LR:-96.62 LO:96.63);ALT=C[chr1:20987374[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	20982726	+	chr1	20987689	+	.	10	0	64396_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=64396_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:20982726(+)-1:20987689(-)__1_20972001_20997001D;SPAN=4963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:0 DR:10 LR:-8.627 LO:19.88);ALT=T[chr1:20987689[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	20998693	+	chr1	21009125	+	.	8	0	64695_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=64695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:20998693(+)-1:21009125(-)__1_20996501_21021501D;SPAN=10432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=A[chr1:21009125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21103245	+	chr1	21106305	+	.	0	37	64913_1	97.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=64913_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_151C;SPAN=3060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:90 GQ:97.7 PL:[97.7, 0.0, 120.8] SR:37 DR:0 LR:-97.75 LO:97.89);ALT=T[chr1:21106305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21106406	+	chr1	21113688	+	.	9	4	64932_1	18.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=64932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_189C;SPAN=7282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:4 DR:9 LR:-18.43 LO:23.96);ALT=T[chr1:21113688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21107034	+	chr1	21113005	+	.	33	6	64936_1	90.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=64936_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_27C;SPAN=5971;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:92 GQ:90.8 PL:[90.8, 0.0, 130.4] SR:6 DR:33 LR:-90.61 LO:91.04);ALT=C[chr1:21113005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21107035	+	chr1	21113686	+	.	34	8	64938_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=64938_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21094501_21119501_122C;SPAN=6651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:67 GQ:57.8 PL:[104.0, 0.0, 57.8] SR:8 DR:34 LR:-104.7 LO:104.7);ALT=T[chr1:21113686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	21180171	+	chr1	21181471	+	.	0	4	65085_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=65085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21168001_21193001_299C;SPAN=1300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:67 GQ:4.8 PL:[0.0, 4.8, 171.6] SR:4 DR:0 LR:4.948 LO:6.824);ALT=C[chr1:21181471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30035108	+	chr1	21724484	+	.	8	0	2767466_1	10.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2767466_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:21724484(-)-6:30035108(+)__6_30012501_30037501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=]chr6:30035108]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	21753941	-	chr1	21806984	+	.	10	0	67044_1	27.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=67044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:21753941(-)-1:21806984(-)__1_21805001_21830001D;SPAN=53043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:19 GQ:17.9 PL:[27.8, 0.0, 17.9] SR:0 DR:10 LR:-27.97 LO:27.97);ALT=[chr1:21806984[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	21822955	+	chr1	21828058	+	.	50	47	67085_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=67085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_21805001_21830001_245C;SPAN=5103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:47 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:47 DR:50 LR:-211.3 LO:211.3);ALT=G[chr1:21828058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	22016595	+	chr1	22021559	+	.	2	2	67840_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=67840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_22001001_22026001_252C;SPAN=4964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:2 DR:2 LR:4.677 LO:6.851);ALT=G[chr1:22021559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	22084278	+	chr1	22109317	+	.	0	8	68253_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=68253_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_22099001_22124001_80C;SPAN=25039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:62 GQ:9.8 PL:[9.8, 0.0, 138.5] SR:8 DR:0 LR:-9.611 LO:16.46);ALT=T[chr1:22109317[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	22271479	-	chr1	22272500	+	.	5	1	68570_1	1.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AAAAGAAAAAAGAAAA;MAPQ=50;MATEID=68570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_22270501_22295501_129C;SPAN=1021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:1 DR:5 LR:-1.062 LO:9.396);ALT=[chr1:22272500[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	22352136	+	chr1	22356770	+	.	19	5	68953_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAG;MAPQ=60;MATEID=68953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_22344001_22369001_279C;SPAN=4634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:79 GQ:44.6 PL:[44.6, 0.0, 146.9] SR:5 DR:19 LR:-44.62 LO:47.68);ALT=G[chr1:22356770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	22379323	+	chr4	22729560	-	.	33	0	1920745_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1920745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:22379323(+)-4:22729560(+)__4_22711501_22736501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:50 GQ:26 PL:[95.3, 0.0, 26.0] SR:0 DR:33 LR:-97.6 LO:97.6);ALT=C]chr4:22729560];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	22413359	+	chr1	22416434	+	.	0	8	69058_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=45;MATEID=69058_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_22393001_22418001_153C;SPAN=3075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:8 DR:0 LR:-3.921 LO:15.38);ALT=G[chr1:22416434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23420916	+	chr1	23495256	+	.	8	0	71555_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=71555_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:23420916(+)-1:23495256(-)__1_23397501_23422501D;SPAN=74340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=A[chr1:23495256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23435622	+	chr1	23495257	+	.	7	2	71918_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=71918_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_23471001_23496001_310C;SPAN=59635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:32 GQ:17.9 PL:[17.9, 0.0, 57.5] SR:2 DR:7 LR:-17.74 LO:19.02);ALT=T[chr1:23495257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23640197	+	chr1	23644971	+	.	7	7	72168_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTACCT;MAPQ=60;MATEID=72168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_23618001_23643001_128C;SPAN=4774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:7 DR:7 LR:-33.7 LO:33.85);ALT=T[chr1:23644971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23648157	+	chr1	23650049	+	.	4	4	72515_1	2.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=72515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_23642501_23667501_42C;SPAN=1892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:4 DR:4 LR:-2.788 LO:13.35);ALT=C[chr1:23650049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23650227	+	chr1	23660008	+	.	0	7	72519_1	3.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=72519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_23642501_23667501_228C;SPAN=9781;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:73 GQ:3.5 PL:[3.5, 0.0, 171.8] SR:7 DR:0 LR:-3.33 LO:13.44);ALT=T[chr1:23660008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23664356	+	chr1	23670702	+	.	9	0	72676_1	19.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=72676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:23664356(+)-1:23670702(-)__1_23667001_23692001D;SPAN=6346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:0 DR:9 LR:-19.68 LO:21.27);ALT=T[chr1:23670702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23665151	+	chr1	23670703	+	.	9	0	72678_1	19.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=72678_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:23665151(+)-1:23670703(-)__1_23667001_23692001D;SPAN=5552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:0 DR:9 LR:-19.41 LO:21.15);ALT=C[chr1:23670703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	23667531	+	chr1	23670702	+	.	13	0	72680_1	22.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=72680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:23667531(+)-1:23670702(-)__1_23667001_23692001D;SPAN=3171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:77 GQ:22.1 PL:[22.1, 0.0, 164.0] SR:0 DR:13 LR:-22.05 LO:28.39);ALT=G[chr1:23670702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	21915188	+	chr1	23670702	+	.	26	0	4539613_1	75.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4539613_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:23670702(-)-10:21915188(+)__10_21903001_21928001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:39 GQ:19.1 PL:[75.2, 0.0, 19.1] SR:0 DR:26 LR:-77.1 LO:77.1);ALT=]chr10:21915188]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	24019249	+	chr1	24021148	+	CTAGATACACTGTCAGATCCTTTGGCATCCGGAGAAATGAAAAGATTGCTGTCCACTGCACAGTTCGAGGGGCCAAGGCAGAAGAAATCTTGGAGAAGGGTCTAA	11	297	74075_1	99.0	.	DISC_MAPQ=11;EVDNC=TSI_G;HOMSEQ=AGGTG;INSERTION=CTAGATACACTGTCAGATCCTTTGGCATCCGGAGAAATGAAAAGATTGCTGTCCACTGCACAGTTCGAGGGGCCAAGGCAGAAGAAATCTTGGAGAAGGGTCTAA;MAPQ=60;MATEID=74075_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_24010001_24035001_104C;SPAN=1899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:308 DP:717 GQ:99 PL:[822.6, 0.0, 918.3] SR:297 DR:11 LR:-822.5 LO:822.8);ALT=G[chr1:24021148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	24117755	+	chr6	33334019	-	.	18	0	2783297_1	41.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=2783297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24117755(+)-6:33334019(+)__6_33320001_33345001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:66 GQ:41.6 PL:[41.6, 0.0, 117.5] SR:0 DR:18 LR:-41.54 LO:43.6);ALT=G]chr6:33334019];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	24144101	+	chr1	24151852	+	.	10	0	73979_1	8.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=73979_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24144101(+)-1:24151852(-)__1_24132501_24157501D;SPAN=7751;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:0 DR:10 LR:-8.627 LO:19.88);ALT=A[chr1:24151852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	24489414	+	chr7	48091486	+	.	2	10	3294628_1	29.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TTCCTTCCTTCCTTCCTTTTCTTT;MAPQ=60;MATEID=3294628_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_48069001_48094001_254C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:14 GQ:2.9 PL:[29.3, 0.0, 2.9] SR:10 DR:2 LR:-30.22 LO:30.22);ALT=T[chr7:48091486[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	24742438	+	chr1	24745791	+	.	8	0	75743_1	17.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=75743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24742438(+)-1:24745791(-)__1_24745001_24770001D;SPAN=3353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=C[chr1:24745791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	24969839	+	chrX	136067839	-	.	62	19	7535206_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7535206_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_23_136048501_136073501_21C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:26 GQ:21 PL:[231.0, 21.0, 0.0] SR:19 DR:62 LR:-231.1 LO:231.1);ALT=G]chrX:136067839];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	24969879	+	chr1	24972474	+	.	8	0	76457_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=76457_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24969879(+)-1:24972474(-)__1_24965501_24990501D;SPAN=2595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.443 LO:16.0);ALT=T[chr1:24972474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	24969882	+	chr1	24973155	+	.	56	0	76459_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=76459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24969882(+)-1:24973155(-)__1_24965501_24990501D;SPAN=3273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:84 GQ:40.1 PL:[162.2, 0.0, 40.1] SR:0 DR:56 LR:-166.1 LO:166.1);ALT=C[chr1:24973155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	24976587	+	chr1	24977897	+	.	8	0	76479_1	4.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=76479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:24976587(+)-1:24977897(-)__1_24965501_24990501D;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=A[chr1:24977897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25158703	+	chr1	25161510	+	.	60	51	77252_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTGATTTTTTATTTTT;MAPQ=60;MATEID=77252_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_25137001_25162001_156C;SPAN=2807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:32 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:51 DR:60 LR:-260.8 LO:260.8);ALT=T[chr1:25161510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25549922	+	chr1	25551492	+	.	3	7	78270_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=78270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25529001_25554001_279C;SPAN=1570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:7 DR:3 LR:-9.39 LO:18.21);ALT=C[chr1:25551492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25554782	+	chr1	25558931	+	.	10	0	78379_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=78379_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25554782(+)-1:25558931(-)__1_25553501_25578501D;SPAN=4149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:121 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.2281 LO:18.52);ALT=C[chr1:25558931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25555615	+	chr1	25558595	+	.	4	51	78381_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=78381_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25553501_25578501_317C;SPAN=2980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:106 GQ:99 PL:[149.6, 0.0, 106.7] SR:51 DR:4 LR:-149.9 LO:149.9);ALT=C[chr1:25558595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25555664	+	chr1	25558930	+	.	50	0	78382_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=78382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25555664(+)-1:25558930(-)__1_25553501_25578501D;SPAN=3266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:113 GQ:99 PL:[134.6, 0.0, 137.9] SR:0 DR:50 LR:-134.4 LO:134.4);ALT=C[chr1:25558930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25571794	+	chr1	25572935	+	.	11	3	78441_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=78441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25553501_25578501_363C;SPAN=1141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:3 DR:11 LR:-26.71 LO:31.54);ALT=T[chr1:25572935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25732108	+	chr1	25613679	+	.	9	3	78820_1	31.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=78820_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_25725001_25750001_270C;SPAN=118429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:29 GQ:31.7 PL:[31.7, 0.0, 38.3] SR:3 DR:9 LR:-31.76 LO:31.79);ALT=]chr1:25732108]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	25664908	+	chr1	25678116	+	.	12	0	78472_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=78472_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25664908(+)-1:25678116(-)__1_25676001_25701001D;SPAN=13208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:35 GQ:30.2 PL:[30.2, 0.0, 53.3] SR:0 DR:12 LR:-30.13 LO:30.52);ALT=C[chr1:25678116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25664911	+	chr1	25669451	+	.	39	0	78319_1	98.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=78319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:25664911(+)-1:25669451(-)__1_25651501_25676501D;SPAN=4540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:110 GQ:98.9 PL:[98.9, 0.0, 168.2] SR:0 DR:39 LR:-98.94 LO:99.92);ALT=C[chr1:25669451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25664947	+	chr1	25666965	+	.	60	41	78320_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=78320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_25651501_25676501_199C;SPAN=2018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:107 GQ:20.6 PL:[238.4, 0.0, 20.6] SR:41 DR:60 LR:-249.1 LO:249.1);ALT=C[chr1:25666965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25667070	+	chr1	25678117	+	TTTTTTACAGGCTGGTGGATTATCATAGATGCAGCTGTTATTTATCCCACCATGAAAGATTTCAACCACTCATACCATGCCTGTGGTGTTATAGCAACCATAGCCTTCCTAAT	0	96	78474_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTTTTACAGGCTGGTGGATTATCATAGATGCAGCTGTTATTTATCCCACCATGAAAGATTTCAACCACTCATACCATGCCTGTGGTGTTATAGCAACCATAGCCTTCCTAAT;MAPQ=60;MATEID=78474_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_25676001_25701001_153C;SPAN=11047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:36 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:96 DR:0 LR:-283.9 LO:283.9);ALT=A[chr1:25678117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25678186	+	chr1	25687150	+	GCTCGCATTTGGCTTTTCGTTGGTTTCATGTTGGCCTTTGGATCTCTGATTGCATCTATGTGGATTCTTTTTGGAGGTTATGTTGCTAAAGAAAAAGACATAGTATACCCTGGAATTGCTGTATTTTTCCAGAATGCCTTCATCTTTTTTG	2	19	78493_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GCTCGCATTTGGCTTTTCGTTGGTTTCATGTTGGCCTTTGGATCTCTGATTGCATCTATGTGGATTCTTTTTGGAGGTTATGTTGCTAAAGAAAAAGACATAGTATACCCTGGAATTGCTGTATTTTTCCAGAATGCCTTCATCTTTTTTG;MAPQ=60;MATEID=78493_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_25676001_25701001_4C;SPAN=8964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:75 GQ:45.8 PL:[45.8, 0.0, 134.9] SR:19 DR:2 LR:-45.7 LO:48.21);ALT=T[chr1:25687150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	25679465	+	chr1	25683282	+	.	3	6	78496_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=78496_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AAAA;SCTG=c_1_25676001_25701001_4C;SPAN=3817;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:65 GQ:2.3 PL:[2.3, 0.0, 154.1] SR:6 DR:3 LR:-2.196 LO:11.41);ALT=G[chr1:25683282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26146554	+	chr1	26149507	+	.	10	0	79609_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=79609_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26146554(+)-1:26149507(-)__1_26141501_26166501D;SPAN=2953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:0 DR:10 LR:-14.86 LO:21.25);ALT=A[chr1:26149507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26146564	+	chr1	26150133	+	.	14	0	79611_1	26.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=79611_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26146564(+)-1:26150133(-)__1_26141501_26166501D;SPAN=3569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:0 DR:14 LR:-26.17 LO:31.35);ALT=T[chr1:26150133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26149619	+	chr1	26152791	+	ACCATCCCAATCTGGCAAAACAAGCCACATGGGGCTGCTCGAAGTGTAGTAAGAAGAATTGGGACCAACCTACCCTTGAAGCCGTGTGCCCGGGCGTCCTTTG	0	28	79617_1	68.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACCATCCCAATCTGGCAAAACAAGCCACATGGGGCTGCTCGAAGTGTAGTAAGAAGAATTGGGACCAACCTACCCTTGAAGCCGTGTGCCCGGGCGTCCTTTG;MAPQ=60;MATEID=79617_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_26141501_26166501_170C;SPAN=3172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:90 GQ:68 PL:[68.0, 0.0, 150.5] SR:28 DR:0 LR:-68.05 LO:69.75);ALT=G[chr1:26152791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26150239	+	chr1	26152791	+	.	0	11	79620_1	14.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=79620_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_1_26141501_26166501_170C;SPAN=2552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:80 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:11 DR:0 LR:-14.64 LO:22.95);ALT=G[chr1:26152791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26228175	+	chr1	26230132	+	.	28	82	79994_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=79994_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_26215001_26240001_186C;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:105 DP:134 GQ:13.4 PL:[310.4, 0.0, 13.4] SR:82 DR:28 LR:-326.4 LO:326.4);ALT=T[chr1:26230132[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26228224	+	chr1	26232878	+	.	18	0	79996_1	7.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=79996_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26228224(+)-1:26232878(-)__1_26215001_26240001D;SPAN=4654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:194 GQ:7 PL:[7.0, 0.0, 462.5] SR:0 DR:18 LR:-6.859 LO:34.29);ALT=G[chr1:26232878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26228230	+	chr1	26231153	+	.	52	0	79997_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=79997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26228230(+)-1:26231153(-)__1_26215001_26240001D;SPAN=2923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:83 GQ:50.3 PL:[149.3, 0.0, 50.3] SR:0 DR:52 LR:-151.7 LO:151.7);ALT=G[chr1:26231153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26230334	+	chr1	26232878	+	.	37	0	80001_1	72.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=80001_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26230334(+)-1:26232878(-)__1_26215001_26240001D;SPAN=2544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:183 GQ:72.7 PL:[72.7, 0.0, 369.8] SR:0 DR:37 LR:-72.56 LO:84.05);ALT=A[chr1:26232878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26460160	+	chr1	26464769	+	.	31	0	80780_1	92.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=80780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:26460160(+)-1:26464769(-)__1_26435501_26460501D;SPAN=4609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:32 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:31 LR:-92.42 LO:92.42);ALT=G[chr1:26464769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26644562	+	chr1	26646657	+	.	96	39	81416_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TACAG;MAPQ=60;MATEID=81416_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_26631501_26656501_208C;SPAN=2095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:121 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:39 DR:96 LR:-356.5 LO:356.5);ALT=G[chr1:26646657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	26759500	+	chr1	26764657	+	.	2	6	81653_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=81653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_26754001_26779001_388C;SPAN=5157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:84 GQ:0.5 PL:[0.5, 0.0, 201.8] SR:6 DR:2 LR:-0.3493 LO:12.99);ALT=G[chr1:26764657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27248357	+	chr2	153246220	+	.	16	0	1046719_1	39.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1046719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27248357(+)-2:153246220(-)__2_153223001_153248001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.0 LO:39.93);ALT=G[chr2:153246220[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	27248361	+	chr1	27250577	+	.	22	0	83384_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=83384_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27248361(+)-1:27250577(-)__1_27244001_27269001D;SPAN=2216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:94 GQ:47.3 PL:[47.3, 0.0, 179.3] SR:0 DR:22 LR:-47.16 LO:51.57);ALT=G[chr1:27250577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27248443	+	chr1	27267945	+	.	26	0	83386_1	54.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=83386_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27248443(+)-1:27267945(-)__1_27244001_27269001D;SPAN=19502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:117 GQ:54.2 PL:[54.2, 0.0, 229.1] SR:0 DR:26 LR:-54.13 LO:60.28);ALT=C[chr1:27267945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27250657	+	chr1	27267946	+	.	0	48	83394_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=83394_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27244001_27269001_22C;SPAN=17289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:96 GQ:99 PL:[132.5, 0.0, 99.5] SR:48 DR:0 LR:-132.7 LO:132.7);ALT=G[chr1:27267946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27527952	+	chr7	132766769	+	.	28	0	3607591_1	64.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=3607591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27527952(+)-7:132766769(-)__7_132765501_132790501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:104 GQ:64.4 PL:[64.4, 0.0, 186.5] SR:0 DR:28 LR:-64.25 LO:67.63);ALT=T[chr7:132766769[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	27648885	+	chr1	27657211	+	.	8	6	84727_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTG;MAPQ=60;MATEID=84727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27636001_27661001_284C;SPAN=8326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:107 GQ:10.7 PL:[10.7, 0.0, 248.3] SR:6 DR:8 LR:-10.62 LO:23.9);ALT=G[chr1:27657211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27648890	+	chr1	27660448	+	.	11	0	84825_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=84825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27648890(+)-1:27660448(-)__1_27660501_27685501D;SPAN=11558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:16 GQ:5.6 PL:[32.0, 0.0, 5.6] SR:0 DR:11 LR:-32.89 LO:32.89);ALT=T[chr1:27660448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27651915	-	chr17	79478280	+	.	14	0	6517656_1	22.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6517656_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27651915(-)-17:79478280(-)__17_79478001_79503001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:88 GQ:22.4 PL:[22.4, 0.0, 190.7] SR:0 DR:14 LR:-22.37 LO:30.18);ALT=[chr17:79478280[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	27657296	+	chr1	27660449	+	AGGACAACATGGCCTTTGGAAAGCCTGCCAA	0	14	84753_1	27.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GTA;INSERTION=AGGACAACATGGCCTTTGGAAAGCCTGCCAA;MAPQ=60;MATEID=84753_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_27636001_27661001_277C;SPAN=3153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:71 GQ:27.2 PL:[27.2, 0.0, 142.7] SR:14 DR:0 LR:-26.98 LO:31.63);ALT=G[chr1:27660449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27668642	+	chr1	27671785	+	.	78	10	84847_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=84847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27660501_27685501_160C;SPAN=3143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:89 GQ:24 PL:[264.0, 24.0, 0.0] SR:10 DR:78 LR:-264.1 LO:264.1);ALT=G[chr1:27671785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27672016	+	chr1	27673909	+	.	6	12	84856_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=84856_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27660501_27685501_143C;SPAN=1893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:12 DR:6 LR:-19.34 LO:27.64);ALT=G[chr1:27673909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27755454	+	chr1	27816503	+	.	32	0	85404_1	91.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=85404_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27755454(+)-1:27816503(-)__1_27807501_27832501D;SPAN=61049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:53 GQ:35.3 PL:[91.4, 0.0, 35.3] SR:0 DR:32 LR:-92.5 LO:92.5);ALT=A[chr1:27816503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27796450	+	chr1	27816497	+	.	0	11	85405_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=85405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27807501_27832501_260C;SPAN=20047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:47 GQ:23.6 PL:[23.6, 0.0, 89.6] SR:11 DR:0 LR:-23.58 LO:25.79);ALT=G[chr1:27816497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27816587	-	chrX	47662621	+	.	29	0	7415900_1	83.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27816587(-)-23:47662621(-)__23_47652501_47677501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:44 GQ:21.2 PL:[83.9, 0.0, 21.2] SR:0 DR:29 LR:-85.73 LO:85.73);ALT=[chrX:47662621[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	27950441	+	chr1	27961574	+	CCTTAGGCCCCTACTCCTGGGTCAGTGGGGCTGCGGCATGATCCTTGGGAGGGGTCAGAG	31	21	85581_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=CCTTAGGCCCCTACTCCTGGGTCAGTGGGGCTGCGGCATGATCCTTGGGAGGGGTCAGAG;MAPQ=60;MATEID=85581_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_27954501_27979501_302C;SPAN=11133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:30 GQ:12 PL:[132.0, 12.0, 0.0] SR:21 DR:31 LR:-132.0 LO:132.0);ALT=C[chr1:27961574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27951665	+	chr1	27961574	+	.	9	8	85582_1	28.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=ACCTG;MAPQ=60;MATEID=85582_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_27954501_27979501_302C;SPAN=9909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:30 GQ:28.1 PL:[28.1, 0.0, 44.6] SR:8 DR:9 LR:-28.18 LO:28.39);ALT=G[chr1:27961574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48481808	+	chr1	27975966	+	.	31	0	1395853_1	86.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=1395853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27975966(-)-3:48481808(+)__3_48461001_48486001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:59 GQ:56.6 PL:[86.3, 0.0, 56.6] SR:0 DR:31 LR:-86.67 LO:86.67);ALT=]chr3:48481808]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	27995096	+	chr1	27998631	+	.	38	0	85776_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=85776_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:27995096(+)-1:27998631(-)__1_27979001_28004001D;SPAN=3535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:78 GQ:84.5 PL:[104.3, 0.0, 84.5] SR:0 DR:38 LR:-104.4 LO:104.4);ALT=G[chr1:27998631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	27995859	+	chr1	27998632	+	.	18	5	85779_1	46.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=85779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_27979001_28004001_130C;SPAN=2773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:72 GQ:46.7 PL:[46.7, 0.0, 125.9] SR:5 DR:18 LR:-46.51 LO:48.63);ALT=T[chr1:27998632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28099936	+	chr1	28116073	+	.	0	11	86113_1	26.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=86113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28101501_28126501_176C;SPAN=16137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:11 DR:0 LR:-26.29 LO:27.14);ALT=A[chr1:28116073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28233554	+	chr1	28240574	+	GTGAAATCTCAACATTCCCAATTCTGAACACTTCATCAACCAAAGTGGCAGAAAGCAGCTGAGATATAGTACAGGGCACAATGTGCTGGGCTCGGGCTCT	0	32	86593_1	81.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=GTGAAATCTCAACATTCCCAATTCTGAACACTTCATCAACCAAAGTGGCAGAAAGCAGCTGAGATATAGTACAGGGCACAATGTGCTGGGCTCGGGCTCT;MAPQ=60;MATEID=86593_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_28224001_28249001_311C;SPAN=7020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:88 GQ:81.8 PL:[81.8, 0.0, 131.3] SR:32 DR:0 LR:-81.79 LO:82.43);ALT=T[chr1:28240574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28233837	+	chr1	28240942	+	.	20	0	86596_1	43.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=86596_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28233837(+)-1:28240942(-)__1_28224001_28249001D;SPAN=7105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:84 GQ:43.4 PL:[43.4, 0.0, 158.9] SR:0 DR:20 LR:-43.26 LO:47.06);ALT=C[chr1:28240942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28384606	+	chr1	28415035	+	.	6	2	87047_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=87047_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AAA;SCTG=c_1_28395501_28420501_211C;SPAN=30429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:55 GQ:8.3 PL:[8.3, 0.0, 123.8] SR:2 DR:6 LR:-8.206 LO:14.35);ALT=C[chr1:28415035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28477601	+	chr1	28503110	+	.	8	0	87443_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=87443_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28477601(+)-1:28503110(-)__1_28493501_28518501D;SPAN=25509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.57 LO:18.13);ALT=A[chr1:28503110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28555536	+	chr1	28559427	+	.	32	11	87658_1	98.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=TTCACCT;MAPQ=60;MATEID=87658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28542501_28567501_63C;SPAN=3891;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:75 GQ:82.1 PL:[98.6, 0.0, 82.1] SR:11 DR:32 LR:-98.58 LO:98.58);ALT=T[chr1:28559427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28559446	-	chr14	35899082	+	.	41	0	5702808_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5702808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28559446(-)-14:35899082(-)__14_35892501_35917501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=[chr14:35899082[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	28562963	+	chr1	28564347	+	.	0	114	87689_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=87689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28542501_28567501_210C;SPAN=1384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:114 DP:177 GQ:99 PL:[328.4, 0.0, 100.7] SR:114 DR:0 LR:-335.0 LO:335.0);ALT=G[chr1:28564347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28696336	+	chr1	28733920	+	.	7	4	88243_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=88243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28714001_28739001_312C;SPAN=37584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:4 DR:7 LR:-18.87 LO:20.92);ALT=G[chr1:28733920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28832645	+	chr1	28835338	+	.	128	0	88659_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=88659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28832645(+)-1:28835338(-)__1_28812001_28837001D;SPAN=2693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:74 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:0 DR:128 LR:-379.6 LO:379.6);ALT=G[chr1:28835338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28897850	+	chr1	28904010	+	ACATATGAAGAAGTTGGAGATGATGCATTGGA	0	13	89033_1	23.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACATATGAAGAAGTTGGAGATGATGCATTGGA;MAPQ=60;MATEID=89033_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_28885501_28910501_349C;SPAN=6160;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:72 GQ:23.6 PL:[23.6, 0.0, 149.0] SR:13 DR:0 LR:-23.41 LO:28.82);ALT=G[chr1:28904010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28905193	+	chr1	28908102	+	CAACTCCATAGGTCCATAGTCACAAATGAGGACAGCTTTACATGTAACATGAATCTCCTCAGTATCACACACTGCCAGGAAACTTGGGGGCAACCAGGTCCCCTGCATTTCATCACTGTCATTACCCCGGAAGTCCTCGATCACCAGAAAAATCACCTTCTGTCATCTTAAGAGTCTTCAT	0	11	89070_1	11.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CAACTCCATAGGTCCATAGTCACAAATGAGGACAGCTTTACATGTAACATGAATCTCCTCAGTATCACACACTGCCAGGAAACTTGGGGGCAACCAGGTCCCCTGCATTTCATCACTGTCATTACCCCGGAAGTCCTCGATCACCAGAAAAATCACCTTCTGTCATCTTAAGAGTCTTCAT;MAPQ=60;MATEID=89070_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_1_28885501_28910501_387C;SPAN=2909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:11 DR:0 LR:-11.39 LO:22.24);ALT=C[chr1:28908102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28944544	+	chr1	28948422	+	.	0	14	88830_1	26.0	.	EVDNC=ASSMB;HOMSEQ=ATACCT;MAPQ=60;MATEID=88830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_28934501_28959501_22C;SPAN=3878;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:73 GQ:26.6 PL:[26.6, 0.0, 148.7] SR:14 DR:0 LR:-26.44 LO:31.44);ALT=T[chr1:28948422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	28948676	+	chr1	28969502	+	.	34	0	89185_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=89185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:28948676(+)-1:28969502(-)__1_28959001_28984001D;SPAN=20826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:0 DR:34 LR:-110.1 LO:110.1);ALT=A[chr1:28969502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29063659	+	chr1	29064769	+	AGACCAAAAGGTCAAGGAAACAA	0	34	89588_1	90.0	.	EVDNC=ASSMB;INSERTION=AGACCAAAAGGTCAAGGAAACAA;MAPQ=60;MATEID=89588_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_29057001_29082001_37C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:81 GQ:90.5 PL:[90.5, 0.0, 103.7] SR:34 DR:0 LR:-90.29 LO:90.36);ALT=G[chr1:29064769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29064850	+	chr1	29068915	+	.	0	8	89594_1	3.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=89594_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_29057001_29082001_294C;SPAN=4065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:8 DR:0 LR:-3.65 LO:15.33);ALT=C[chr1:29068915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29064851	+	chr1	29095441	+	.	0	8	89595_1	16.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=89595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_29057001_29082001_361C;SPAN=30590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:8 DR:0 LR:-16.65 LO:18.55);ALT=G[chr1:29095441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29476706	+	chr1	29481206	+	.	2	9	90770_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=90770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_29473501_29498501_43C;SPAN=4500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:9 DR:2 LR:-9.932 LO:18.32);ALT=T[chr1:29481206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29487030	+	chr1	29508158	+	.	0	11	91178_1	24.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=91178_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_29498001_29523001_228C;SPAN=21128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:44 GQ:24.5 PL:[24.5, 0.0, 80.6] SR:11 DR:0 LR:-24.39 LO:26.15);ALT=C[chr1:29508158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	29845254	+	chr2	142301926	+	.	8	18	91793_1	66.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TCTTCTTCTTCTTCTACTTCTTCTTCTCCTC;MAPQ=60;MATEID=91793_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_29841001_29866001_48C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:17 GQ:6 PL:[66.0, 6.0, 0.0] SR:18 DR:8 LR:-66.02 LO:66.02);ALT=C[chr2:142301926[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	30738623	+	chr1	30739932	+	.	48	32	93508_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCA;MAPQ=60;MATEID=93508_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_30723001_30748001_14C;SPAN=1309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:36 GQ:18 PL:[198.0, 18.0, 0.0] SR:32 DR:48 LR:-198.0 LO:198.0);ALT=A[chr1:30739932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31206766	+	chr1	31208017	+	.	10	11	94632_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=94632_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_31188501_31213501_83C;SPAN=1251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:98 GQ:36.2 PL:[36.2, 0.0, 201.2] SR:11 DR:10 LR:-36.17 LO:42.77);ALT=T[chr1:31208017[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31206812	+	chr1	31210448	+	.	14	0	94633_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=94633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31206812(+)-1:31210448(-)__1_31188501_31213501D;SPAN=3636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:80 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:0 DR:14 LR:-24.54 LO:30.82);ALT=G[chr1:31210448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31208114	+	chr1	31210449	+	.	2	5	94638_1	3.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=94638_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_31188501_31213501_295C;SPAN=2335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:73 GQ:3.5 PL:[3.5, 0.0, 171.8] SR:5 DR:2 LR:-3.33 LO:13.44);ALT=T[chr1:31210449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31210547	+	chr1	31211787	+	.	3	3	94648_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=94648_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_1_31188501_31213501_295C;SPAN=1240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:85 GQ:3 PL:[0.0, 3.0, 211.2] SR:3 DR:3 LR:3.223 LO:10.69);ALT=C[chr1:31211787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31214612	+	chr1	31230553	+	.	98	0	94531_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=94531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31214612(+)-1:31230553(-)__1_31213001_31238001D;SPAN=15941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:118 GQ:5.4 PL:[297.0, 5.4, 0.0] SR:0 DR:98 LR:-310.9 LO:310.9);ALT=C[chr1:31230553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31215397	+	chr1	31230506	+	.	102	28	94534_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=94534_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_31213001_31238001_235C;SPAN=15109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:127 GQ:14.4 PL:[336.6, 14.4, 0.0] SR:28 DR:102 LR:-345.9 LO:345.9);ALT=C[chr1:31230506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31532427	+	chr1	31538459	+	.	12	0	95607_1	15.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=95607_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31532427(+)-1:31538459(-)__1_31531501_31556501D;SPAN=6032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:89 GQ:15.5 PL:[15.5, 0.0, 200.3] SR:0 DR:12 LR:-15.5 LO:24.93);ALT=A[chr1:31538459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31568380	+	chr19	48282071	-	CGCCA	84	30	6842369_1	99.0	.	DISC_MAPQ=7;EVDNC=ASDIS;INSERTION=CGCCA;MAPQ=60;MATEID=6842369_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48265001_48290001_363C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:47 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:30 DR:84 LR:-310.3 LO:310.3);ALT=G]chr19:48282071];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	31624520	-	chr1	31625812	+	.	8	0	96206_1	7.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=96206_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31624520(-)-1:31625812(-)__1_31605001_31630001D;SPAN=1292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:0 DR:8 LR:-6.901 LO:15.9);ALT=[chr1:31625812[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	31764853	+	chr1	31766066	+	.	0	10	96505_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=96505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_31752001_31777001_118C;SPAN=1213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:10 DR:0 LR:-12.69 LO:20.72);ALT=A[chr1:31766066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31766225	+	chr1	31769543	+	.	17	0	96510_1	32.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=96510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31766225(+)-1:31769543(-)__1_31752001_31777001D;SPAN=3318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:87 GQ:32.6 PL:[32.6, 0.0, 177.8] SR:0 DR:17 LR:-32.55 LO:38.33);ALT=C[chr1:31769543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31769974	+	chr1	31791953	+	.	15	0	96526_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=96526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31769974(+)-1:31791953(-)__1_31752001_31777001D;SPAN=21979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:55 GQ:34.7 PL:[34.7, 0.0, 97.4] SR:0 DR:15 LR:-34.61 LO:36.33);ALT=C[chr1:31791953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31770069	+	chr1	31782902	+	.	8	0	96529_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=96529_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:31770069(+)-1:31782902(-)__1_31752001_31777001D;SPAN=12833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=T[chr1:31782902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31783013	+	chr1	31791954	+	.	2	17	96348_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=96348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_31776501_31801501_303C;SPAN=8941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:85 GQ:39.8 PL:[39.8, 0.0, 165.2] SR:17 DR:2 LR:-39.69 LO:44.11);ALT=T[chr1:31791954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31810122	+	chr1	31819487	+	ATGAAAAATGATAGAATAAAAGTATCCCTCTCCATGAAGGTTGTCAATCAAGGGACTGGGAAAGACCTTGATCCCAACAATGTTATCATTGA	0	20	96650_1	44.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGAAAAATGATAGAATAAAAGTATCCCTCTCCATGAAGGTTGTCAATCAAGGGACTGGGAAAGACCTTGATCCCAACAATGTTATCATTGA;MAPQ=60;MATEID=96650_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_31801001_31826001_322C;SPAN=9365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:82 GQ:44 PL:[44.0, 0.0, 152.9] SR:20 DR:0 LR:-43.8 LO:47.3);ALT=G[chr1:31819487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	31821822	+	chr1	31836877	+	.	4	6	96684_1	23.0	.	DISC_MAPQ=11;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=96684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_31801001_31826001_149C;SPAN=15055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:34 GQ:23.9 PL:[23.9, 0.0, 56.9] SR:6 DR:4 LR:-23.8 LO:24.62);ALT=G[chr1:31836877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32098916	+	chr1	32100821	+	.	0	11	97354_1	12.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=97354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32095001_32120001_172C;SPAN=1905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:11 DR:0 LR:-12.74 LO:22.52);ALT=C[chr1:32100821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32101089	+	chr1	32110440	+	.	23	0	97361_1	48.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=97361_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32101089(+)-1:32110440(-)__1_32095001_32120001D;SPAN=9351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:102 GQ:48.5 PL:[48.5, 0.0, 197.0] SR:0 DR:23 LR:-48.29 LO:53.49);ALT=G[chr1:32110440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32374588	+	chr1	32377295	+	.	8	0	98270_1	2.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=98270_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32374588(+)-1:32377295(-)__1_32364501_32389501D;SPAN=2707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=A[chr1:32377295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32479978	+	chr1	32495896	+	.	8	10	98656_1	38.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=98656_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_1_32462501_32487501_33C;SPAN=15918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:27 GQ:25.7 PL:[38.9, 0.0, 25.7] SR:10 DR:8 LR:-39.02 LO:39.02);ALT=G[chr1:32495896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32479978	+	chr1	32497123	+	AAATTGAGAAGATTCAGAAAGGAGACTCAAAAAAGGATGATGAGGAGAATTACTTGGATTTATTTTCTCATAAGAACATGAAACTGAAAGAGCGAGTGCTGATACCTGTCAAGCAGTATCCCA	6	13	98657_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAATTGAGAAGATTCAGAAAGGAGACTCAAAAAAGGATGATGAGGAGAATTACTTGGATTTATTTTCTCATAAGAACATGAAACTGAAAGAGCGAGTGCTGATACCTGTCAAGCAGTATCCCA;MAPQ=60;MATEID=98657_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_32462501_32487501_33C;SPAN=17145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:27 GQ:12.5 PL:[52.1, 0.0, 12.5] SR:13 DR:6 LR:-53.38 LO:53.38);ALT=G[chr1:32497123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32496023	+	chr1	32497123	+	.	4	7	98345_1	13.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=98345_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_32487001_32512001_204C;SPAN=1100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:7 DR:4 LR:-13.5 LO:20.92);ALT=G[chr1:32497123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32498936	+	chr1	32502510	+	.	8	3	98360_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=98360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32487001_32512001_86C;SPAN=3574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:3 DR:8 LR:-11.34 LO:20.42);ALT=G[chr1:32502510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32505175	+	chr1	32508127	+	.	7	4	98380_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=98380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32487001_32512001_319C;SPAN=2952;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:4 DR:7 LR:-4.242 LO:17.27);ALT=G[chr1:32508127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32667700	+	chr1	32669478	+	.	0	7	98971_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=98971_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32658501_32683501_249C;SPAN=1778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:69 GQ:4.4 PL:[4.4, 0.0, 162.8] SR:7 DR:0 LR:-4.413 LO:13.62);ALT=G[chr1:32669478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32688221	+	chr1	32690009	+	.	52	0	99289_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=99289_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32688221(+)-1:32690009(-)__1_32683001_32708001D;SPAN=1788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:102 GQ:99 PL:[144.2, 0.0, 101.3] SR:0 DR:52 LR:-144.4 LO:144.4);ALT=C[chr1:32690009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32688221	+	chr1	32691767	+	.	23	0	99290_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=99290_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32688221(+)-1:32691767(-)__1_32683001_32708001D;SPAN=3546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:89 GQ:51.8 PL:[51.8, 0.0, 164.0] SR:0 DR:23 LR:-51.81 LO:55.07);ALT=C[chr1:32691767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32688231	+	chr1	32689635	+	.	47	46	99292_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=99292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32683001_32708001_238C;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:86 GQ:23 PL:[184.7, 0.0, 23.0] SR:46 DR:47 LR:-191.8 LO:191.8);ALT=T[chr1:32689635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32689723	+	chr1	32691769	+	GGACACCAAGCATGTCCTCACTGGCTCAGCTGACAACAGCTGTCGTCTCTGGGACTGTGAAA	0	123	99300_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=GGACACCAAGCATGTCCTCACTGGCTCAGCTGACAACAGCTGTCGTCTCTGGGACTGTGAAA;MAPQ=60;MATEID=99300_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_32683001_32708001_66C;SPAN=2046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:98 GQ:33 PL:[363.0, 33.0, 0.0] SR:123 DR:0 LR:-363.1 LO:363.1);ALT=G[chr1:32691769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32690077	+	chr1	32691769	+	.	4	73	99301_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=46;MATEID=99301_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_32683001_32708001_66C;SPAN=1692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:74 DP:106 GQ:40.7 PL:[215.6, 0.0, 40.7] SR:73 DR:4 LR:-222.2 LO:222.2);ALT=G[chr1:32691769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32694811	+	chr1	32696524	+	.	0	10	99322_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CCAGGT;MAPQ=60;MATEID=99322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32683001_32708001_167C;SPAN=1713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:10 DR:0 LR:-14.59 LO:21.18);ALT=T[chr1:32696524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32757834	+	chr1	32782259	+	.	18	0	99521_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=99521_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32757834(+)-1:32782259(-)__1_32756501_32781501D;SPAN=24425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:36 GQ:36.5 PL:[49.7, 0.0, 36.5] SR:0 DR:18 LR:-49.75 LO:49.75);ALT=C[chr1:32782259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32757840	+	chr1	32768220	+	.	19	0	99522_1	38.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=99522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:32757840(+)-1:32768220(-)__1_32756501_32781501D;SPAN=10380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:88 GQ:38.9 PL:[38.9, 0.0, 174.2] SR:0 DR:19 LR:-38.88 LO:43.78);ALT=G[chr1:32768220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32768334	+	chr1	32782266	+	.	0	29	99568_1	82.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=99568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32756501_32781501_318C;SPAN=13932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:49 GQ:36.2 PL:[82.4, 0.0, 36.2] SR:29 DR:0 LR:-83.42 LO:83.42);ALT=T[chr1:32782266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	32782383	+	chr1	32790080	+	.	0	10	99435_1	13.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=99435_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_32781001_32806001_310C;SPAN=7697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:10 DR:0 LR:-12.96 LO:20.79);ALT=T[chr1:32790080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33099749	+	chr1	33116064	+	.	11	0	101375_1	18.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=101375_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:33099749(+)-1:33116064(-)__1_33099501_33124501D;SPAN=16315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:0 DR:11 LR:-18.43 LO:23.96);ALT=A[chr1:33116064[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33276660	+	chr1	33282788	+	.	14	12	100955_1	46.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=100955_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_33271001_33296001_43C;SPAN=6128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:85 GQ:46.4 PL:[46.4, 0.0, 158.6] SR:12 DR:14 LR:-46.29 LO:49.8);ALT=T[chr1:33282788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33283343	+	chr1	33291697	+	.	8	0	100980_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=100980_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:33283343(+)-1:33291697(-)__1_33271001_33296001D;SPAN=8354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:69 GQ:7.7 PL:[7.7, 0.0, 159.5] SR:0 DR:8 LR:-7.714 LO:16.06);ALT=G[chr1:33291697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33476415	+	chr2	32048487	+	.	11	0	101764_1	22.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=101764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:33476415(+)-2:32048487(-)__1_33467001_33492001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:0 DR:11 LR:-22.49 LO:25.34);ALT=C[chr2:32048487[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	33476436	+	chr1	33478825	+	.	8	0	101766_1	0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=101766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:33476436(+)-1:33478825(-)__1_33467001_33492001D;SPAN=2389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=T[chr1:33478825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	33885514	+	chr7	39749694	+	.	0	28	3264209_1	77.0	.	EVDNC=ASSMB;HOMSEQ=CCTC;MAPQ=60;MATEID=3264209_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_39739001_39764001_306C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:55 GQ:54.5 PL:[77.6, 0.0, 54.5] SR:28 DR:0 LR:-77.71 LO:77.71);ALT=C[chr7:39749694[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	35321630	+	chr1	35325267	+	.	24	0	106082_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=106082_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:35321630(+)-1:35325267(-)__1_35304501_35329501D;SPAN=3637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:76 GQ:58.7 PL:[58.7, 0.0, 124.7] SR:0 DR:24 LR:-58.63 LO:59.98);ALT=C[chr1:35325267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35447721	+	chr1	35450799	+	CATCATGAGCAGAATCAAGAACAAGTTACTGATCTCTTGCAGCATCGGTGGGCCCATGACCAGCAGCAACCCAGCCAGCAGTTCCAGAAAGCCCACAGCTATTTGGTAGTTCAGGGGATCTGGCTGGTAGCCAAATACCTTCAGCGGGAACACCTCAGCAAACTGCACGAACAGGGCATT	0	17	106407_1	35.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATCATGAGCAGAATCAAGAACAAGTTACTGATCTCTTGCAGCATCGGTGGGCCCATGACCAGCAGCAACCCAGCCAGCAGTTCCAGAAAGCCCACAGCTATTTGGTAGTTCAGGGGATCTGGCTGGTAGCCAAATACCTTCAGCGGGAACACCTCAGCAAACTGCACGAACAGGGCATT;MAPQ=60;MATEID=106407_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_35427001_35452001_272C;SPAN=3078;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:77 GQ:35.3 PL:[35.3, 0.0, 150.8] SR:17 DR:0 LR:-35.26 LO:39.36);ALT=C[chr1:35450799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35449601	+	chr1	35450813	+	.	33	0	106412_1	87.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=106412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:35449601(+)-1:35450813(-)__1_35427001_35452001D;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:80 GQ:87.2 PL:[87.2, 0.0, 107.0] SR:0 DR:33 LR:-87.26 LO:87.37);ALT=C[chr1:35450813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35650195	+	chr1	35652602	+	.	3	15	107006_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=107006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_35647501_35672501_54C;SPAN=2407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:15 DR:3 LR:-32.87 LO:40.05);ALT=C[chr1:35652602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35650243	+	chr1	35653573	+	.	8	0	107008_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=107008_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:35650243(+)-1:35653573(-)__1_35647501_35672501D;SPAN=3330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=T[chr1:35653573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35652725	+	chr1	35654603	+	CCCATGTTCATTGCTCCTCCGCCACCCATTCGCATGTCTCTTTCCCGTGGATCCATGTAGCCCATTCGGCTGTAACTTTCCTCTCTTTGGCGCCTCATTTGTTCTTCCATCTCACGTTGACGAATCATCATCTCTTCCTCTCTTCTACGTCGTTCCTCCTCTTG	0	45	107014_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CCCATGTTCATTGCTCCTCCGCCACCCATTCGCATGTCTCTTTCCCGTGGATCCATGTAGCCCATTCGGCTGTAACTTTCCTCTCTTTGGCGCCTCATTTGTTCTTCCATCTCACGTTGACGAATCATCATCTCTTCCTCTCTTCTACGTCGTTCCTCCTCTTG;MAPQ=60;MATEID=107014_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_35647501_35672501_22C;SPAN=1878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:88 GQ:88.4 PL:[124.7, 0.0, 88.4] SR:45 DR:0 LR:-125.0 LO:125.0);ALT=T[chr1:35654603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	35654983	+	chr1	35656098	+	.	17	25	107025_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=107025_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_35647501_35672501_341C;SPAN=1115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:87 GQ:99 PL:[101.9, 0.0, 108.5] SR:25 DR:17 LR:-101.9 LO:101.9);ALT=C[chr1:35656098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36035522	+	chr1	36039960	+	.	0	12	108101_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=108101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36015001_36040001_308C;SPAN=4438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:67 GQ:21.5 PL:[21.5, 0.0, 140.3] SR:12 DR:0 LR:-21.46 LO:26.55);ALT=T[chr1:36039960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36068977	+	chr1	36096875	+	CCTCCAGACATTTCCTAAGGAGTTCCACTGCCCTCTCACGTGAGATAGTCGGTGTGTAGTATCGGTCGAGGATACTGAGAGTCAGGAAGGCACCATAGCCGTGGGCTGCAAAAGGGGCCTTGGCCAAGGCTGCCAGGTAGTCCATGTAATACAGCGCTGGCCCTTCATGCTCATCATAGCCAGCCAGGAGGAGGTTCACATGATATGGGGT	0	36	108124_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCTCCAGACATTTCCTAAGGAGTTCCACTGCCCTCTCACGTGAGATAGTCGGTGTGTAGTATCGGTCGAGGATACTGAGAGTCAGGAAGGCACCATAGCCGTGGGCTGCAAAAGGGGCCTTGGCCAAGGCTGCCAGGTAGTCCATGTAATACAGCGCTGGCCCTTCATGCTCATCATAGCCAGCCAGGAGGAGGTTCACATGATATGGGGT;MAPQ=60;MATEID=108124_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_36064001_36089001_390C;SPAN=27898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:49 GQ:13.1 PL:[105.5, 0.0, 13.1] SR:36 DR:0 LR:-109.7 LO:109.7);ALT=T[chr1:36096875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36070883	+	chr1	36074847	+	.	2	20	108129_1	41.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=108129_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_36064001_36089001_390C;SPAN=3964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:89 GQ:41.9 PL:[41.9, 0.0, 173.9] SR:20 DR:2 LR:-41.91 LO:46.48);ALT=G[chr1:36074847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36075010	+	chr1	36096875	+	.	2	9	108342_1	20.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=108342_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_36088501_36113501_236C;SPAN=21865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:9 DR:2 LR:-20.87 LO:24.74);ALT=C[chr1:36096875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36096946	+	chr1	36101910	+	.	3	30	108374_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=108374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36088501_36113501_303C;SPAN=4964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:101 GQ:75.2 PL:[75.2, 0.0, 167.6] SR:30 DR:3 LR:-74.97 LO:77.0);ALT=C[chr1:36101910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36102034	+	chr1	36106943	+	.	66	62	108395_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=108395_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36088501_36113501_108C;SPAN=4909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:96 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:62 DR:66 LR:-283.9 LO:283.9);ALT=C[chr1:36106943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36181927	+	chr1	36184307	+	.	8	6	108627_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=108627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36162001_36187001_224C;SPAN=2380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:6 DR:8 LR:-8.898 LO:19.93);ALT=C[chr1:36184307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36605420	+	chr1	36614938	+	ATTTTGTCCAGCTGTTTATTCACATCTTCATCATTTTCATAGTCCTTACATAGCTGGGTGACCAGGGCACCATAGGTCAGGGTGAAGAGCTCAGAGCT	13	30	109670_1	91.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATTTTGTCCAGCTGTTTATTCACATCTTCATCATTTTCATAGTCCTTACATAGCTGGGTGACCAGGGCACCATAGGTCAGGGTGAAGAGCTCAGAGCT;MAPQ=60;MATEID=109670_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_36603001_36628001_206C;SPAN=9518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:89 GQ:91.4 PL:[91.4, 0.0, 124.4] SR:30 DR:13 LR:-91.42 LO:91.7);ALT=C[chr1:36614938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36605820	+	chr1	36615013	+	.	16	0	109672_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=109672_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36605820(+)-1:36615013(-)__1_36603001_36628001D;SPAN=9193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:115 GQ:21.8 PL:[21.8, 0.0, 256.1] SR:0 DR:16 LR:-21.66 LO:33.48);ALT=T[chr1:36615013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36690137	+	chr1	36724979	+	.	12	0	110356_1	27.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=110356_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36690137(+)-1:36724979(-)__1_36701001_36726001D;SPAN=34842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:44 GQ:27.8 PL:[27.8, 0.0, 77.3] SR:0 DR:12 LR:-27.69 LO:29.07);ALT=C[chr1:36724979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36690152	+	chr1	36748129	+	.	34	0	110059_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=110059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36690152(+)-1:36748129(-)__1_36725501_36750501D;SPAN=57977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:32 GQ:9 PL:[99.0, 9.0, 0.0] SR:0 DR:34 LR:-99.02 LO:99.02);ALT=T[chr1:36748129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36725087	+	chr1	36748132	+	.	0	19	110061_1	53.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=110061_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36725501_36750501_32C;SPAN=23045;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:34 GQ:27.2 PL:[53.6, 0.0, 27.2] SR:19 DR:0 LR:-53.9 LO:53.9);ALT=T[chr1:36748132[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36733250	+	chr1	36734642	-	AAA	28	60	110077_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAA;MAPQ=60;MATEID=110077_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_36725501_36750501_152C;SPAN=1392;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:67 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:60 DR:28 LR:-247.6 LO:247.6);ALT=A]chr1:36734642];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	36748301	+	chr1	36751967	+	.	3	13	110153_1	41.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=110153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36750001_36775001_318C;SPAN=3666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:42 GQ:41.6 PL:[41.6, 0.0, 58.1] SR:13 DR:3 LR:-41.44 LO:41.63);ALT=G[chr1:36751967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36859755	+	chr1	36863368	+	.	65	24	110817_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=110817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36848001_36873001_338C;SPAN=3613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:91 GQ:8.6 PL:[209.9, 0.0, 8.6] SR:24 DR:65 LR:-220.4 LO:220.4);ALT=C[chr1:36863368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36927824	+	chr1	36929867	+	.	11	0	110671_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=110671_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36927824(+)-1:36929867(-)__1_36921501_36946501D;SPAN=2043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:0 DR:11 LR:-13.82 LO:22.76);ALT=C[chr1:36929867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36943278	+	chr1	36945033	+	.	0	11	110711_1	15.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=110711_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_36921501_36946501_198C;SPAN=1755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:11 DR:0 LR:-15.45 LO:23.15);ALT=C[chr1:36945033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36943294	+	chr1	36948409	+	.	8	0	110729_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=110729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:36943294(+)-1:36948409(-)__1_36946001_36971001D;SPAN=5115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:30 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.28 LO:19.28);ALT=G[chr1:36948409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36945118	+	chr1	36948412	+	AGCTTTGTGATCTTGGACAAGTTACTTCACCTTTCCGAGCCGAGCCTCAGTTTCCCCAT	24	26	110731_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGCTTTGTGATCTTGGACAAGTTACTTCACCTTTCCGAGCCGAGCCTCAGTTTCCCCAT;MAPQ=60;MATEID=110731_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_36946001_36971001_303C;SPAN=3294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:31 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:26 DR:24 LR:-115.5 LO:115.5);ALT=C[chr1:36948412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	36947138	+	chr1	36948412	+	.	9	6	110737_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=110737_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_1_36946001_36971001_303C;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:6 DR:9 LR:-15.72 LO:23.22);ALT=T[chr1:36948412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	37423181	+	chr1	37425549	+	C	3	23	112226_1	64.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=0;MATEID=112226_2;MATENM=0;NM=1;NUMPARTS=2;REPSEQ=CCC;SCTG=c_1_37411501_37436501_308C;SECONDARY;SPAN=2368;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:81 GQ:64.1 PL:[64.1, 0.0, 130.1] SR:23 DR:3 LR:-63.88 LO:65.21);ALT=C[chr1:37425549[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	37975143	+	chr1	37979024	+	.	2	18	113441_1	52.0	.	DISC_MAPQ=30;EVDNC=ASDIS;MAPQ=60;MATEID=113441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_37950501_37975501_380C;SPAN=3881;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:39 GQ:42.2 PL:[52.1, 0.0, 42.2] SR:18 DR:2 LR:-52.2 LO:52.2);ALT=T[chr1:37979024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	37975184	+	chr1	37980276	+	.	23	0	113586_1	57.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=113586_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:37975184(+)-1:37980276(-)__1_37975001_38000001D;SPAN=5092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:69 GQ:57.2 PL:[57.2, 0.0, 110.0] SR:0 DR:23 LR:-57.23 LO:58.15);ALT=T[chr1:37980276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	37979140	+	chr1	37980257	+	.	36	15	113595_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=113595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_37975001_38000001_17C;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:71 GQ:43.7 PL:[126.2, 0.0, 43.7] SR:15 DR:36 LR:-128.0 LO:128.0);ALT=C[chr1:37980257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38058409	+	chr1	38061360	+	GCGCTCCTTTTGCCTATACATATTCAGGCGCCGGATGGTGGCCCGGTCCCTCATGTTTTGGCCTCCTGCTCCCTGCACTCGAT	0	26	113799_1	65.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GCGCTCCTTTTGCCTATACATATTCAGGCGCCGGATGGTGGCCCGGTCCCTCATGTTTTGGCCTCCTGCTCCCTGCACTCGAT;MAPQ=60;MATEID=113799_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_38048501_38073501_80C;SPAN=2951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:75 GQ:65.6 PL:[65.6, 0.0, 115.1] SR:26 DR:0 LR:-65.51 LO:66.29);ALT=T[chr1:38061360[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38059496	+	chr1	38061441	+	.	14	0	113802_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=113802_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:38059496(+)-1:38061441(-)__1_38048501_38073501D;SPAN=1945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:96 GQ:20.3 PL:[20.3, 0.0, 211.7] SR:0 DR:14 LR:-20.21 LO:29.6);ALT=T[chr1:38061441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11422016	+	chr1	38241383	+	.	10	24	6730983_1	90.0	.	DISC_MAPQ=49;EVDNC=ASDIS;MAPQ=60;MATEID=6730983_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_19_11417001_11442001_269C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:44 GQ:14.6 PL:[90.5, 0.0, 14.6] SR:24 DR:10 LR:-93.33 LO:93.33);ALT=]chr19:11422016]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	38323346	+	chr1	38325202	+	.	12	0	114559_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=114559_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:38323346(+)-1:38325202(-)__1_38318001_38343001D;SPAN=1856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:91 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:0 DR:12 LR:-14.96 LO:24.81);ALT=A[chr1:38325202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38465106	+	chr1	38471028	+	.	0	8	115070_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=115070_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_38440501_38465501_290C;SPAN=5922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:8 DR:0 LR:-15.3 LO:18.03);ALT=T[chr1:38471028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38478537	+	chr1	38484134	+	CCTGGCTTTCGAAAACATCTGGGCCTGCTGGAGAAAAAGAAAGATTACAAACTTCGTGCAGATGACTACCGTAAAAAACAAGAATACCTCAAAGCTCTTCGGAAGAAGGCTCTTGAAAAAAATCCAGATGAATTCTACTACAAAATGACTCGGGTTAAACTCC	2	12	114950_1	20.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CCTGGCTTTCGAAAACATCTGGGCCTGCTGGAGAAAAAGAAAGATTACAAACTTCGTGCAGATGACTACCGTAAAAAACAAGAATACCTCAAAGCTCTTCGGAAGAAGGCTCTTGAAAAAAATCCAGATGAATTCTACTACAAAATGACTCGGGTTAAACTCC;MAPQ=60;MATEID=114950_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_38465001_38490001_219C;SPAN=5597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:12 DR:2 LR:-20.7 LO:28.0);ALT=G[chr1:38484134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38478537	+	chr1	38483338	+	.	12	0	114949_1	17.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=114949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:38478537(+)-1:38483338(-)__1_38465001_38490001D;SPAN=4801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:84 GQ:17 PL:[17.0, 0.0, 185.3] SR:0 DR:12 LR:-16.85 LO:25.26);ALT=G[chr1:38483338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	38478537	+	chr1	38482029	+	.	5	6	114948_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=114948_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_38465001_38490001_219C;SPAN=3492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:6 DR:5 LR:2.36 LO:12.64);ALT=G[chr1:38482029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39330388	+	chr1	39332552	+	.	0	18	117113_1	41.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=117113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_39322501_39347501_49C;SPAN=2164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:66 GQ:41.6 PL:[41.6, 0.0, 117.5] SR:18 DR:0 LR:-41.54 LO:43.6);ALT=T[chr1:39332552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39332709	+	chr1	39338960	+	.	14	0	117123_1	26.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=117123_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:39332709(+)-1:39338960(-)__1_39322501_39347501D;SPAN=6251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:0 DR:14 LR:-26.71 LO:31.54);ALT=T[chr1:39338960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39492070	+	chr1	39494394	+	.	117	5	117884_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=117884_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_39494001_39519001_2C;SPAN=2324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:43 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:5 DR:117 LR:-346.6 LO:346.6);ALT=G[chr1:39494394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39492106	+	chr17	27348522	-	.	43	0	117765_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=117765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:39492106(+)-17:27348522(+)__1_39469501_39494501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:34 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=A]chr17:27348522];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	39492109	+	chr1	39500062	+	.	9	0	117766_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=117766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:39492109(+)-1:39500062(-)__1_39469501_39494501D;SPAN=7953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=T[chr1:39500062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	39696917	+	chr1	39715684	+	.	0	8	118840_1	14.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=118840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_39690001_39715001_393C;SPAN=18767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:8 DR:0 LR:-14.49 LO:17.76);ALT=T[chr1:39715684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40204647	+	chr1	40207034	+	.	12	0	120067_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=120067_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40204647(+)-1:40207034(-)__1_40204501_40229501D;SPAN=2387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:0 DR:12 LR:-19.29 LO:25.9);ALT=C[chr1:40207034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40204649	+	chr1	40208885	+	.	13	0	120069_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=120069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40204649(+)-1:40208885(-)__1_40204501_40229501D;SPAN=4236;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:74 GQ:23 PL:[23.0, 0.0, 155.0] SR:0 DR:13 LR:-22.86 LO:28.64);ALT=C[chr1:40208885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40205935	+	chr1	40209493	+	AAAAGCACCGAGGATTTGCTTTTGTTGAATTTGAGTTGGCAGAGGATGCTGCAGCAGCTATCGACAACATGAATGAATCTGAGCTTTTTGGACGTACAATTCGTGTCAATTTGGCCAAACCAATGAGAATTAAGGAAGGCTCTTCCAGGC	0	30	120074_1	77.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AAAAGCACCGAGGATTTGCTTTTGTTGAATTTGAGTTGGCAGAGGATGCTGCAGCAGCTATCGACAACATGAATGAATCTGAGCTTTTTGGACGTACAATTCGTGTCAATTTGGCCAAACCAATGAGAATTAAGGAAGGCTCTTCCAGGC;MAPQ=60;MATEID=120074_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_40204501_40229501_196C;SPAN=3558;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:78 GQ:77.9 PL:[77.9, 0.0, 110.9] SR:30 DR:0 LR:-77.9 LO:78.22);ALT=G[chr1:40209493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40506513	+	chr1	40525006	+	.	18	0	121103_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=121103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40506513(+)-1:40525006(-)__1_40523001_40548001D;SPAN=18493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:52 GQ:45.5 PL:[45.5, 0.0, 78.5] SR:0 DR:18 LR:-45.33 LO:45.88);ALT=G[chr1:40525006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40506524	+	chr1	40525736	+	.	33	0	121105_1	92.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=121105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40506524(+)-1:40525736(-)__1_40523001_40548001D;SPAN=19212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:59 GQ:50 PL:[92.9, 0.0, 50.0] SR:0 DR:33 LR:-93.63 LO:93.63);ALT=G[chr1:40525736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40525843	+	chr1	40527407	+	.	0	24	121116_1	57.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=121116_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_40523001_40548001_280C;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:81 GQ:57.5 PL:[57.5, 0.0, 136.7] SR:24 DR:0 LR:-57.28 LO:59.17);ALT=G[chr1:40527407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40527484	+	chr1	40529899	+	.	0	8	121117_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=121117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_40523001_40548001_225C;SPAN=2415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:8 DR:0 LR:-1.212 LO:14.96);ALT=A[chr1:40529899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40557846	+	chr1	40562786	+	CCATCAGGGTCTTCCCAATCTCTAAAGATAAGACGTAAATTCCAGGTATTTTCTTCTCCACCATTTTTTTAATAGCACCCATGCTTAAGGGATTGCAACAGCTGTCT	0	56	120959_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CCATCAGGGTCTTCCCAATCTCTAAAGATAAGACGTAAATTCCAGGTATTTTCTTCTCCACCATTTTTTTAATAGCACCCATGCTTAAGGGATTGCAACAGCTGTCT;MAPQ=60;MATEID=120959_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_40547501_40572501_72C;SPAN=4940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:87 GQ:49.1 PL:[161.3, 0.0, 49.1] SR:56 DR:0 LR:-164.5 LO:164.5);ALT=T[chr1:40562786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40558228	+	chr1	40562854	+	.	65	0	120961_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=120961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:40558228(+)-1:40562854(-)__1_40547501_40572501D;SPAN=4626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:98 GQ:49.4 PL:[188.0, 0.0, 49.4] SR:0 DR:65 LR:-192.5 LO:192.5);ALT=T[chr1:40562854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	40839896	+	chr1	40872406	+	.	2	3	122214_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=122214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_40817001_40842001_367C;SPAN=32510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:35 GQ:3.8 PL:[3.8, 0.0, 79.7] SR:3 DR:2 LR:-3.722 LO:8.002);ALT=G[chr1:40872406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	41157539	+	chr1	41204506	+	.	7	5	122913_1	12.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=122913_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_41184501_41209501_351C;SPAN=46967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:5 DR:7 LR:-12.86 LO:17.27);ALT=G[chr1:41204506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	41445503	+	chr1	41448947	+	.	8	1	123653_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=123653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_41429501_41454501_311C;SPAN=3444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:1 DR:8 LR:-10.97 LO:16.77);ALT=T[chr1:41448947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	42922316	+	chr6	136741384	-	.	15	0	127170_1	38.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=127170_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:42922316(+)-6:136741384(+)__1_42899501_42924501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:41 GQ:38.6 PL:[38.6, 0.0, 58.4] SR:0 DR:15 LR:-38.41 LO:38.69);ALT=C]chr6:136741384];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	42922318	+	chr1	42925264	+	.	38	0	127171_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=127171_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:42922318(+)-1:42925264(-)__1_42899501_42924501D;SPAN=2946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:42 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:38 LR:-122.1 LO:122.1);ALT=G[chr1:42925264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	42923021	+	chr1	42925271	+	.	6	31	127173_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=127173_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_42899501_42924501_156C;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:40 GQ:7.5 PL:[112.2, 7.5, 0.0] SR:31 DR:6 LR:-113.5 LO:113.5);ALT=G[chr1:42925271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	43124184	+	chr11	111901010	-	CATGCGGCCAACTT	65	6	5004785_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CATGCGGCCAACTT;MAPQ=60;MATEID=5004785_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_11_111891501_111916501_91C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:40 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:6 DR:65 LR:-208.0 LO:208.0);ALT=G]chr11:111901010];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	43124195	+	chr1	43130532	+	.	9	0	127703_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=127703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:43124195(+)-1:43130532(-)__1_43120001_43145001D;SPAN=6337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:0 DR:9 LR:-5.597 LO:17.5);ALT=G[chr1:43130532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	43133112	+	chr1	43142253	+	.	0	58	127727_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=127727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_43120001_43145001_127C;SPAN=9141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:109 GQ:99 PL:[161.9, 0.0, 102.5] SR:58 DR:0 LR:-162.6 LO:162.6);ALT=G[chr1:43142253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	43630477	+	chr1	43632496	+	.	0	14	129037_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=129037_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_43610001_43635001_80C;SPAN=2019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:85 GQ:23.3 PL:[23.3, 0.0, 181.7] SR:14 DR:0 LR:-23.19 LO:30.41);ALT=C[chr1:43632496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	43831334	+	chr1	43833585	+	.	32	0	129737_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=129737_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:43831334(+)-1:43833585(-)__1_43806001_43831001D;SPAN=2251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:0 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=T[chr1:43833585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	44173366	+	chr1	44201903	+	.	13	8	130669_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=130669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_44198001_44223001_289C;SPAN=28537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:46 GQ:50.3 PL:[50.3, 0.0, 60.2] SR:8 DR:13 LR:-50.26 LO:50.32);ALT=T[chr1:44201903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	44372365	+	chr1	44370282	+	.	9	0	131046_1	9.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=131046_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:44370282(-)-1:44372365(+)__1_44369501_44394501D;SPAN=2083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=]chr1:44372365]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	44372446	+	chr1	44371397	+	.	22	0	131052_1	56.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=131052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:44371397(-)-1:44372446(+)__1_44369501_44394501D;SPAN=1049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:60 GQ:56.3 PL:[56.3, 0.0, 89.3] SR:0 DR:22 LR:-56.37 LO:56.77);ALT=]chr1:44372446]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	44440811	+	chr1	44441972	+	.	19	0	131242_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=131242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:44440811(+)-1:44441972(-)__1_44418501_44443501D;SPAN=1161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:96 GQ:36.8 PL:[36.8, 0.0, 195.2] SR:0 DR:19 LR:-36.71 LO:42.96);ALT=A[chr1:44441972[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	44750579	+	chr1	44773981	+	.	0	9	132320_1	18.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=132320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_44761501_44786501_263C;SPAN=23402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:9 DR:0 LR:-18.6 LO:20.81);ALT=C[chr1:44773981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	44774075	+	chr1	44785300	+	CCAGCACTTGCTGCAGGCTTGGCTGACCATCCACCATGGCTTGAATAATCCCGGTGAG	6	11	132343_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCAGCACTTGCTGCAGGCTTGGCTGACCATCCACCATGGCTTGAATAATCCCGGTGAG;MAPQ=60;MATEID=132343_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_44761501_44786501_242C;SPAN=11225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:78 GQ:25.1 PL:[25.1, 0.0, 163.7] SR:11 DR:6 LR:-25.08 LO:30.99);ALT=T[chr1:44785300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	44871199	+	chr1	44877652	+	.	12	17	132406_1	54.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=132406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_44859501_44884501_206C;SPAN=6453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:91 GQ:54.8 PL:[54.8, 0.0, 163.7] SR:17 DR:12 LR:-54.57 LO:57.72);ALT=G[chr1:44877652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45235827	+	chr1	45236960	-	.	8	0	133601_1	4.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=133601_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45235827(+)-1:45236960(+)__1_45227001_45252001D;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:0 DR:8 LR:-4.192 LO:15.42);ALT=A]chr1:45236960];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	45241307	+	chr1	45242343	+	.	8	0	133617_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=133617_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45241307(+)-1:45242343(-)__1_45227001_45252001D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:151 GQ:14.2 PL:[0.0, 14.2, 392.7] SR:0 DR:8 LR:14.5 LO:13.22);ALT=A[chr1:45242343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45316677	+	chr1	45323376	+	.	0	11	133723_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=133723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_45300501_45325501_241C;SPAN=6699;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:11 DR:0 LR:-13.28 LO:22.64);ALT=T[chr1:45323376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45446850	+	chr1	45452165	+	.	17	2	134105_1	50.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=134105_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_45447501_45472501_284C;SPAN=5315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:45 GQ:50.6 PL:[50.6, 0.0, 57.2] SR:2 DR:17 LR:-50.53 LO:50.56);ALT=C[chr1:45452165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45977088	+	chr1	45980179	+	.	4	42	136020_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=53;MATEID=136020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_45962001_45987001_55C;SPAN=3091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:81 GQ:67.4 PL:[126.8, 0.0, 67.4] SR:42 DR:4 LR:-127.5 LO:127.5);ALT=T[chr1:45980179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45980668	+	chr1	45984609	+	ATGCTAGATGACAGAAGTGAGAATCCACAGAAGCACCAATCACTTGGCAGTTGAGTTTCTTAAATTCTTCTGCCCTATCACTGAAAGCAATGATCTCCGTGGGGCACACAAAGGTGAAGTCAAGAGGGTAAAAGAAGAACACAACATATTTT	2	163	136029_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GAGATGCCTTCATCAGCCTTTAAGACCCCATAATCCTGAGCAATGGTGCGCTTCGGGTCTGATACCAAAGGAATGTTCATGGGTCCCAGTCCTCCTTGTTTCTTAGGTGTATTGACCCATGCTAGATGACAGAAGTGAGAATCCACAGAAGCACCAATCACTTGGCAGTTGAGTTTCTTAAATTCTTCTGCCCTATCACTGAAAGCAATGATCTCCGTGGGGCACACAAAGGTGAAGTCAAGAGGGTAAAAGAAGAACACAACATATTTTCCT;INSERTION=ATGCTAGATGACAGAAGTGAGAATCCACAGAAGCACCAATCACTTGGCAGTTGAGTTTCTTAAATTCTTCTGCCCTATCACTGAAAGCAATGATCTCCGTGGGGCACACAAAGGTGAAGTCAAGAGGGTAAAAGAAGAACACAACATATTTT;MAPQ=60;MATEID=136029_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_45962001_45987001_248C;SECONDARY;SPAN=3941;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:163 DP:109 GQ:43.9 PL:[481.9, 43.9, 0.0] SR:163 DR:2 LR:-481.9 LO:481.9);ALT=C[chr1:45984609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45981481	+	chr1	45984609	+	.	5	125	136034_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=136034_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_45962001_45987001_248C;SPAN=3128;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:131 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:125 DR:5 LR:-386.2 LO:386.2);ALT=T[chr1:45984609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45981520	+	chr1	45987349	+	.	174	0	136055_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=136055_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45981520(+)-1:45987349(-)__1_45986501_46011501D;SPAN=5829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:45 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:0 DR:174 LR:-514.9 LO:514.9);ALT=A[chr1:45987349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	45984765	+	chr1	45987381	+	.	79	0	136057_1	99.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=136057_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:45984765(+)-1:45987381(-)__1_45986501_46011501D;SPAN=2616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:52 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=T[chr1:45987381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46016828	+	chr1	46027459	+	.	20	18	135741_1	93.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=135741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46011001_46036001_270C;SPAN=10631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:82 GQ:93.5 PL:[93.5, 0.0, 103.4] SR:18 DR:20 LR:-93.32 LO:93.36);ALT=G[chr1:46027459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46016829	+	chr1	46018106	+	.	15	3	135742_1	31.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=135742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46011001_46036001_208C;SPAN=1277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:68 GQ:31.1 PL:[31.1, 0.0, 133.4] SR:3 DR:15 LR:-31.09 LO:34.72);ALT=T[chr1:46018106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46016876	+	chr1	46032232	+	.	33	0	135744_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=135744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46016876(+)-1:46032232(-)__1_46011001_46036001D;SPAN=15356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=T[chr1:46032232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46018236	+	chr1	46027459	+	.	0	8	135748_1	3.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=135748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46011001_46036001_173C;SPAN=9223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:8 DR:0 LR:-3.109 LO:15.25);ALT=G[chr1:46027459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46027552	+	chr1	46032238	+	.	0	24	135771_1	53.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=135771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46011001_46036001_356C;SPAN=4686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:97 GQ:53 PL:[53.0, 0.0, 181.7] SR:24 DR:0 LR:-52.94 LO:56.94);ALT=T[chr1:46032238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46049805	+	chr1	46067923	+	.	38	0	136446_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=136446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46049805(+)-1:46067923(-)__1_46035501_46060501D;SPAN=18118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:44 GQ:8.4 PL:[122.1, 8.4, 0.0] SR:0 DR:38 LR:-122.5 LO:122.5);ALT=A[chr1:46067923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46068037	+	chr1	46072152	+	AGGTAAGAAGTATGGAGAGACAGCTAATGAGTGTGGAGAAGCCTTCTTTTTCTATGGGAAATCACTTCTGGAGTTGGCA	0	53	135840_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGGTAAGAAGTATGGAGAGACAGCTAATGAGTGTGGAGAAGCCTTCTTTTTCTATGGGAAATCACTTCTGGAGTTGGCA;MAPQ=60;MATEID=135840_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_46060001_46085001_136C;SPAN=4115;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:85 GQ:53 PL:[152.0, 0.0, 53.0] SR:53 DR:0 LR:-154.5 LO:154.5);ALT=T[chr1:46072152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46126949	+	chr1	46152129	+	.	18	0	135943_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=135943_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46126949(+)-1:46152129(-)__1_46109001_46134001D;SPAN=25180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:29 GQ:18.5 PL:[51.5, 0.0, 18.5] SR:0 DR:18 LR:-52.4 LO:52.4);ALT=T[chr1:46152129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46153952	+	chr8	98866023	-	.	9	0	3986936_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3986936_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46153952(+)-8:98866023(+)__8_98857501_98882501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:0 DR:9 LR:-19.41 LO:21.15);ALT=A]chr8:98866023];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	46153955	+	chr1	46156644	+	.	14	0	136246_1	29.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=136246_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46153955(+)-1:46156644(-)__1_46133501_46158501D;SPAN=2689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:64 GQ:29 PL:[29.0, 0.0, 124.7] SR:0 DR:14 LR:-28.88 LO:32.35);ALT=T[chr1:46156644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46153989	+	chr1	46158910	+	.	10	0	136499_1	23.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=136499_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:46153989(+)-1:46158910(-)__1_46158001_46183001D;SPAN=4921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=T[chr1:46158910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	46156782	+	chr1	46158874	+	.	0	15	136255_1	41.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=136255_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_46133501_46158501_143C;SPAN=2092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:31 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:15 DR:0 LR:-41.15 LO:41.15);ALT=G[chr1:46158874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	47046301	+	chr1	47048900	+	.	0	12	139294_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=139294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_47040001_47065001_226C;SPAN=2599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:77 GQ:18.8 PL:[18.8, 0.0, 167.3] SR:12 DR:0 LR:-18.75 LO:25.75);ALT=T[chr1:47048900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	47049004	+	chr1	47059785	+	.	0	12	139302_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CTA;MAPQ=60;MATEID=139302_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_47040001_47065001_120C;SPAN=10781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:77 GQ:18.8 PL:[18.8, 0.0, 167.3] SR:12 DR:0 LR:-18.75 LO:25.75);ALT=A[chr1:47059785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	47799788	+	chr1	47834139	+	.	0	13	141511_1	31.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=141511_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_47824001_47849001_137C;SPAN=34351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:44 GQ:31.1 PL:[31.1, 0.0, 74.0] SR:13 DR:0 LR:-30.99 LO:32.03);ALT=G[chr1:47834139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	45872386	+	chr1	47804186	+	.	60	42	2830453_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TCCCT;MAPQ=60;MATEID=2830453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_45864001_45889001_51C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:29 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:42 DR:60 LR:-211.3 LO:211.3);ALT=]chr6:45872386]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	123386971	+	chr1	48033106	+	.	7	13	141892_1	53.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=GAAATCCTGTCTCTACTAAAAATACAAAAA;MAPQ=60;MATEID=141892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_48020001_48045001_339C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:46 GQ:53.6 PL:[53.6, 0.0, 56.9] SR:13 DR:7 LR:-53.56 LO:53.57);ALT=]chr12:123386971]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	48691544	+	chr1	48692816	-	.	9	0	143365_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=143365_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:48691544(+)-1:48692816(+)__1_48681501_48706501D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=T]chr1:48692816];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	59004955	+	chr1	59012332	+	.	9	0	168400_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=168400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:59004955(+)-1:59012332(-)__1_58996001_59021001D;SPAN=7377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=G[chr1:59012332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	59096879	+	chr2	32048671	+	.	38	0	168730_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=168730_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:59096879(+)-2:32048671(-)__1_59094001_59119001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:64 GQ:45.5 PL:[108.2, 0.0, 45.5] SR:0 DR:38 LR:-109.4 LO:109.4);ALT=A[chr2:32048671[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	59956710	-	chr8	6536461	+	.	9	0	3726855_1	23.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=3726855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:59956710(-)-8:6536461(-)__8_6517001_6542001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:23 GQ:23.6 PL:[23.6, 0.0, 30.2] SR:0 DR:9 LR:-23.48 LO:23.56);ALT=[chr8:6536461[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	1324318	+	chr1	70319124	+	.	0	27	1885317_1	82.0	.	EVDNC=ASSMB;HOMSEQ=GCT;MAPQ=60;MATEID=1885317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1323001_1348001_38C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:27 DR:0 LR:-82.52 LO:82.52);ALT=]chr4:1324318]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	9946094	+	chr1	70385246	+	.	13	0	6725258_1	28.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=6725258_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:70385246(-)-19:9946094(+)__19_9922501_9947501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:55 GQ:28.1 PL:[28.1, 0.0, 104.0] SR:0 DR:13 LR:-28.01 LO:30.54);ALT=]chr19:9946094]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	70671508	+	chr1	70687295	+	.	27	0	195285_1	80.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=195285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:70671508(+)-1:70687295(-)__1_70658001_70683001D;SPAN=15787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:34 GQ:0.8 PL:[80.0, 0.0, 0.8] SR:0 DR:27 LR:-84.31 LO:84.31);ALT=T[chr1:70687295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70687522	+	chr1	70694105	+	.	0	17	195198_1	30.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=195198_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_70682501_70707501_226C;SPAN=6583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:96 GQ:30.2 PL:[30.2, 0.0, 201.8] SR:17 DR:0 LR:-30.11 LO:37.52);ALT=A[chr1:70694105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70698060	+	chr1	70700376	+	.	2	8	195225_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=195225_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_1_70682501_70707501_255C;SPAN=2316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:8 DR:2 LR:-7.764 LO:17.89);ALT=G[chr1:70700376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70698060	+	chr1	70703108	+	ATTGGCGCTGTTCCACTGGCTGCTTTGGGGGCTCCTACTCTTGATCCTGCCCTTGCTGCACTTGGGCTTCCTGGAGCAAACTTGAACTCTCAGTCTCTTGCTGCAGATCAGTTGCTGAAGCTTATGAGTACTGTTGATCCCAA	0	23	195226_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=ATTGGCGCTGTTCCACTGGCTGCTTTGGGGGCTCCTACTCTTGATCCTGCCCTTGCTGCACTTGGGCTTCCTGGAGCAAACTTGAACTCTCAGTCTCTTGCTGCAGATCAGTTGCTGAAGCTTATGAGTACTGTTGATCCCAA;MAPQ=60;MATEID=195226_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_70682501_70707501_255C;SPAN=5048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:72 GQ:56.6 PL:[56.6, 0.0, 116.0] SR:23 DR:0 LR:-56.42 LO:57.62);ALT=G[chr1:70703108[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70703235	+	chr1	70710365	+	ATAAGAAAGAAGAAAAAAGAAGGCATTCAAGATCAAGATCACGTTCTAGGAGGAGGAGGACTCCCTCATCTTCTAGACAC	5	63	195307_1	99.0	.	DISC_MAPQ=53;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATAAGAAAGAAGAAAAAAGAAGGCATTCAAGATCAAGATCACGTTCTAGGAGGAGGAGGACTCCCTCATCTTCTAGACAC;MAPQ=60;MATEID=195307_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_70707001_70732001_112C;SPAN=7130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:49 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:63 DR:5 LR:-188.1 LO:188.1);ALT=G[chr1:70710365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70703235	+	chr1	70705120	+	.	2	30	195241_1	81.0	.	DISC_MAPQ=35;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=195241_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_70682501_70707501_101C;SPAN=1885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:91 GQ:81.2 PL:[81.2, 0.0, 137.3] SR:30 DR:2 LR:-80.98 LO:81.84);ALT=G[chr1:70705120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70710498	+	chr1	70712499	+	.	3	16	195318_1	39.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=195318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_70707001_70732001_251C;SPAN=2001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:74 GQ:39.5 PL:[39.5, 0.0, 138.5] SR:16 DR:3 LR:-39.37 LO:42.55);ALT=G[chr1:70712499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	70712590	+	chr1	70715633	+	.	0	13	195324_1	23.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=195324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_70707001_70732001_292C;SPAN=3043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:74 GQ:23 PL:[23.0, 0.0, 155.0] SR:13 DR:0 LR:-22.86 LO:28.64);ALT=G[chr1:70715633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	71535050	+	chr1	71536508	+	.	3	3	197271_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCTGGA;MAPQ=60;MATEID=197271_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_71515501_71540501_134C;SPAN=1458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:3 DR:3 LR:5.711 LO:8.577);ALT=A[chr1:71536508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	71538233	+	chr1	71542477	+	.	0	7	197170_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=197170_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_71540001_71565001_190C;SPAN=4244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:27 GQ:15.8 PL:[15.8, 0.0, 48.8] SR:7 DR:0 LR:-15.79 LO:16.77);ALT=T[chr1:71542477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	71542560	+	chr1	71544140	+	.	0	30	197179_1	78.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=197179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_71540001_71565001_311C;SPAN=1580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:77 GQ:78.2 PL:[78.2, 0.0, 107.9] SR:30 DR:0 LR:-78.17 LO:78.44);ALT=A[chr1:71544140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	71544249	+	chr1	71546623	+	CCGACCACATCGATTACAGCTGGTTCTTCTAGCAAAGTTTACATTTCCACAT	0	32	197184_1	82.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCGACCACATCGATTACAGCTGGTTCTTCTAGCAAAGTTTACATTTCCACAT;MAPQ=60;MATEID=197184_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_71540001_71565001_274C;SPAN=2374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:85 GQ:82.7 PL:[82.7, 0.0, 122.3] SR:32 DR:0 LR:-82.6 LO:83.05);ALT=C[chr1:71546623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	71544391	+	chr1	71546623	+	.	44	9	197185_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=197185_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_1_71540001_71565001_274C;SPAN=2232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:73 GQ:29.9 PL:[145.4, 0.0, 29.9] SR:9 DR:44 LR:-149.4 LO:149.4);ALT=T[chr1:71546623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	72400997	+	chr1	72748000	+	.	3	4	199476_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTA;MAPQ=60;MATEID=199476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_72740501_72765501_50C;SPAN=347003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:30 GQ:5 PL:[5.0, 0.0, 67.7] SR:4 DR:3 LR:-5.076 LO:8.289);ALT=A[chr1:72748000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	72740291	-	chr10	5827814	+	.	11	0	4500058_1	29.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=4500058_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:72740291(-)-10:5827814(-)__10_5806501_5831501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:25 GQ:29.6 PL:[29.6, 0.0, 29.6] SR:0 DR:11 LR:-29.54 LO:29.54);ALT=[chr10:5827814[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	72766324	+	chr1	72811840	+	.	0	57	199343_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=199343_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_72789501_72814501_31C;SPAN=45516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:14 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:57 DR:0 LR:-168.3 LO:168.3);ALT=G[chr1:72811840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84517932	-	chrX	76411859	+	.	15	0	7454454_1	42.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7454454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:84517932(-)-23:76411859(-)__23_76391001_76416001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:27 GQ:22.4 PL:[42.2, 0.0, 22.4] SR:0 DR:15 LR:-42.49 LO:42.49);ALT=[chrX:76411859[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	84517939	+	chr1	84524630	+	.	41	15	224957_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGATTTGTTTTTCT;MAPQ=60;MATEID=224957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84500501_84525501_206C;SPAN=6691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:62 GQ:6.5 PL:[141.8, 0.0, 6.5] SR:15 DR:41 LR:-148.6 LO:148.6);ALT=T[chr1:84524630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84644921	+	chr1	84647881	+	.	0	10	224723_1	15.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=224723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84623001_84648001_294C;SPAN=2960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:10 DR:0 LR:-15.67 LO:21.47);ALT=G[chr1:84647881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84712005	+	chr1	84715875	+	GTGCACAAT	22	12	225130_1	78.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTGCACAAT;MAPQ=60;MATEID=225130_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84696501_84721501_273C;SPAN=3870;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:63 GQ:72.2 PL:[78.8, 0.0, 72.2] SR:12 DR:22 LR:-78.67 LO:78.67);ALT=T[chr1:84715875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84945193	+	chr1	84946637	+	.	0	12	225668_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=225668_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84941501_84966501_116C;SPAN=1444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:12 DR:0 LR:-17.67 LO:25.46);ALT=G[chr1:84946637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84962053	+	chr1	84963110	+	.	0	16	225710_1	30.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=225710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84941501_84966501_330C;SPAN=1057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:84 GQ:30.2 PL:[30.2, 0.0, 172.1] SR:16 DR:0 LR:-30.06 LO:35.88);ALT=G[chr1:84963110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	84964231	+	chr1	84971692	+	.	19	6	225723_1	59.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=225723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_84941501_84966501_42C;SPAN=7461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:51 GQ:59 PL:[59.0, 0.0, 62.3] SR:6 DR:19 LR:-58.81 LO:58.82);ALT=C[chr1:84971692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	109590094	+	chr1	84971740	+	.	53	0	225534_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=225534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:84971740(-)-23:109590094(+)__1_84966001_84991001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:72 GQ:17 PL:[155.6, 0.0, 17.0] SR:0 DR:53 LR:-161.6 LO:161.6);ALT=]chrX:109590094]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	85036405	+	chr1	85039919	+	.	21	22	225842_1	79.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GACCT;MAPQ=60;MATEID=225842_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_85039501_85064501_202C;SPAN=3514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:47 GQ:33.5 PL:[79.7, 0.0, 33.5] SR:22 DR:21 LR:-80.67 LO:80.67);ALT=T[chr1:85039919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	86392749	-	chr10	25707687	+	.	2	21	229513_1	58.0	.	DISC_MAPQ=5;EVDNC=ASDIS;MAPQ=47;MATEID=229513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_86387001_86412001_289C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:54 GQ:58.1 PL:[58.1, 0.0, 71.3] SR:21 DR:2 LR:-57.99 LO:58.09);ALT=[chr10:25707687[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	86680740	+	chr1	86683024	+	.	26	15	229825_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAACATTGTCTTTG;MAPQ=60;MATEID=229825_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_86681001_86706001_105C;SPAN=2284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:28 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:15 DR:26 LR:-95.72 LO:95.72);ALT=G[chr1:86683024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	87170654	+	chr1	87181404	+	.	33	15	231018_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=231018_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_87146501_87171501_143C;SPAN=10750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:29 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:15 DR:33 LR:-112.2 LO:112.2);ALT=G[chr1:87181404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	87337011	+	chr10	33386453	-	AGAAGGCCATGCAGAGGAAGAACCCTGGAGAGGAGCCCTGGGGTCTCCAGATGAGAGAGAAGATGAA	24	31	4568626_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;INSERTION=AGAAGGCCATGCAGAGGAAGAACCCTGGAGAGGAGCCCTGGGGTCTCCAGATGAGAGAGAAGATGAA;MAPQ=60;MATEID=4568626_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_10_33369001_33394001_162C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:31 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:31 DR:24 LR:-145.2 LO:145.2);ALT=T]chr10:33386453];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	87337011	+	chr10	36119127	-	.	13	22	4573145_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=4573145_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_36113001_36138001_13C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:31 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:22 DR:13 LR:-89.12 LO:89.12);ALT=T]chr10:36119127];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	87346457	+	chr1	87379731	+	.	26	0	231279_1	75.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=231279_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:87346457(+)-1:87379731(-)__1_87342501_87367501D;SPAN=33274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:17 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:0 DR:26 LR:-75.92 LO:75.92);ALT=G[chr1:87379731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	87365171	+	chr6	38932141	+	.	8	0	2805851_1	22.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2805851_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:87365171(+)-6:38932141(-)__6_38930501_38955501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:15 GQ:12.5 PL:[22.4, 0.0, 12.5] SR:0 DR:8 LR:-22.44 LO:22.44);ALT=G[chr6:38932141[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	87369132	+	chr1	87379708	+	.	74	16	231094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=231094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_87367001_87392001_123C;SPAN=10576;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:61 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:16 DR:74 LR:-237.7 LO:237.7);ALT=C[chr1:87379708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49371052	+	chr1	87512502	+	.	9	0	5491089_1	16.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5491089_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:87512502(-)-13:49371052(+)__13_49367501_49392501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-15.89 LO:19.85);ALT=]chr13:49371052]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	88336599	+	chr16	83666361	+	AAA	7	31	232810_1	99.0	.	DISC_MAPQ=8;EVDNC=ASDIS;INSERTION=AAA;MAPQ=13;MATEID=232810_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_88322501_88347501_134C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:33 GQ:9 PL:[99.0, 9.0, 0.0] SR:31 DR:7 LR:-99.02 LO:99.02);ALT=A[chr16:83666361[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	88972810	-	chr17	32063850	+	.	48	19	6371204_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6371204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_32046001_32071001_107C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:41 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:19 DR:48 LR:-158.4 LO:158.4);ALT=[chr17:32063850[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	88972825	+	chr17	32064663	-	C	20	21	6371205_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=6371205_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_32046001_32071001_448C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:46 GQ:2.4 PL:[115.5, 2.4, 0.0] SR:21 DR:20 LR:-120.3 LO:120.3);ALT=T]chr17:32064663];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	89150312	+	chr1	89206669	+	.	0	8	233795_1	19.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=233795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_89204501_89229501_2C;SPAN=56357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:8 DR:0 LR:-19.36 LO:19.88);ALT=G[chr1:89206669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89325971	+	chr1	89329663	+	.	4	3	234069_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=234069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_89302501_89327501_166C;SPAN=3692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:20 GQ:17.6 PL:[17.6, 0.0, 30.8] SR:3 DR:4 LR:-17.69 LO:17.88);ALT=T[chr1:89329663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89329800	+	chr1	89352940	+	.	0	8	233947_1	18.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=TCACCTA;MAPQ=60;MATEID=233947_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_1_89351501_89376501_200C;SPAN=23140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:8 DR:0 LR:-18.82 LO:19.57);ALT=A[chr1:89352940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89329838	+	chr1	89357165	+	.	9	0	233990_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=233990_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:89329838(+)-1:89357165(-)__1_89327001_89352001D;SPAN=27327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=A[chr1:89357165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89353051	+	chr1	89357166	+	.	14	4	233952_1	26.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=233952_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_89351501_89376501_200C;SPAN=4115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:4 DR:14 LR:-26.71 LO:31.54);ALT=C[chr1:89357166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89434498	+	chr1	89458268	+	ACACATTACTATCAAGTCCTTCAATCCGTTTTGCATTTGTGAATTTCAGTGACATTTT	4	16	234240_1	49.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ACACATTACTATCAAGTCCTTCAATCCGTTTTGCATTTGTGAATTTCAGTGACATTTT;MAPQ=60;MATEID=234240_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_89449501_89474501_221C;SPAN=23770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:26 GQ:12.8 PL:[49.1, 0.0, 12.8] SR:16 DR:4 LR:-50.15 LO:50.15);ALT=C[chr1:89458268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89435199	+	chr1	89458368	+	.	8	0	234242_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=234242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:89435199(+)-1:89458368(-)__1_89449501_89474501D;SPAN=23169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:25 GQ:19.7 PL:[19.7, 0.0, 39.5] SR:0 DR:8 LR:-19.64 LO:20.05);ALT=A[chr1:89458368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89570519	+	chr12	57081784	+	.	125	0	5205294_1	99.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=5205294_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:89570519(+)-12:57081784(-)__12_57060501_57085501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:72 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:0 DR:125 LR:-369.7 LO:369.7);ALT=T[chr12:57081784[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	89573976	+	chr1	89575359	+	.	0	5	234348_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=234348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_89572001_89597001_112C;SPAN=1383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:5 DR:0 LR:-3.23 LO:9.742);ALT=T[chr1:89575359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	89587667	+	chr1	89591545	+	.	4	2	234368_1	0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=234368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_89572001_89597001_11C;SPAN=3878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:59 GQ:2.7 PL:[0.0, 2.7, 148.5] SR:2 DR:4 LR:2.781 LO:7.052);ALT=C[chr1:89591545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	90460820	+	chr1	90470560	+	.	14	0	235642_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=235642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:90460820(+)-1:90470560(-)__1_90454001_90479001D;SPAN=9740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:64 GQ:29 PL:[29.0, 0.0, 124.7] SR:0 DR:14 LR:-28.88 LO:32.35);ALT=G[chr1:90470560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	90487905	+	chr1	90492911	+	.	6	2	235805_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=235805_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_90478501_90503501_144C;SPAN=5006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:61 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:2 DR:6 LR:-6.581 LO:14.02);ALT=G[chr1:90492911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	91267672	+	chr6	32468802	+	.	10	0	2777922_1	29.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=2777922_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:91267672(+)-6:32468802(-)__6_32462501_32487501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:10 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:10 LR:-29.71 LO:29.71);ALT=T[chr6:32468802[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	91561367	+	chr1	93514541	+	.	9	0	240896_1	22.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=240896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:91561367(+)-1:93514541(-)__1_93492001_93517001D;SPAN=1953174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:26 GQ:22.7 PL:[22.7, 0.0, 39.2] SR:0 DR:9 LR:-22.67 LO:22.94);ALT=G[chr1:93514541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	92764704	+	chr1	92767030	+	.	14	0	239508_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=239508_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:92764704(+)-1:92767030(-)__1_92757001_92782001D;SPAN=2326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:42 GQ:35 PL:[35.0, 0.0, 64.7] SR:0 DR:14 LR:-34.84 LO:35.4);ALT=G[chr1:92767030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	92767148	+	chr1	92769534	+	.	0	7	239511_1	9.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=239511_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_92757001_92782001_236C;SPAN=2386;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=G[chr1:92769534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93297682	+	chr1	93299099	+	.	50	0	240745_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=240745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93297682(+)-1:93299099(-)__1_93296001_93321001D;SPAN=1417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:128 GQ:99 PL:[130.4, 0.0, 179.9] SR:0 DR:50 LR:-130.4 LO:130.8);ALT=G[chr1:93299099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93297689	+	chr1	93300333	+	.	21	0	240750_1	47.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=240750_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93297689(+)-1:93300333(-)__1_93296001_93321001D;SPAN=2644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:83 GQ:47 PL:[47.0, 0.0, 152.6] SR:0 DR:21 LR:-46.83 LO:50.06);ALT=C[chr1:93300333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93300470	+	chr1	93301746	+	.	11	97	240761_1	99.0	.	DISC_MAPQ=15;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=240761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_93296001_93321001_254C;SPAN=1276;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:90 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:97 DR:11 LR:-320.2 LO:320.2);ALT=G[chr1:93301746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93301968	+	chr1	93303023	+	.	19	0	240774_1	21.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=240774_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93301968(+)-1:93303023(-)__1_93296001_93321001D;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:152 GQ:21.8 PL:[21.8, 0.0, 345.2] SR:0 DR:19 LR:-21.54 LO:38.8);ALT=A[chr1:93303023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93545088	+	chr1	93575785	+	.	6	8	241160_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=241160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_93565501_93590501_260C;SPAN=30697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:29 GQ:28.4 PL:[28.4, 0.0, 41.6] SR:8 DR:6 LR:-28.45 LO:28.6);ALT=G[chr1:93575785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93805158	+	chr1	93811280	+	.	59	0	241420_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=241420_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:93805158(+)-1:93811280(-)__1_93810501_93835501D;SPAN=6122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:19 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=T[chr1:93811280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	93806070	+	chr1	93811281	+	GAGGATCACCAACTTGAGAGCTTTGTTTG	16	9	241421_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;INSERTION=GAGGATCACCAACTTGAGAGCTTTGTTTG;MAPQ=60;MATEID=241421_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_93810501_93835501_145C;SPAN=5211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:19 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:9 DR:16 LR:-56.11 LO:56.11);ALT=G[chr1:93811281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	94288375	+	chr1	94291257	+	.	69	27	242166_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CCA;MAPQ=60;MATEID=242166_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_94276001_94301001_16C;SPAN=2882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:22 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:27 DR:69 LR:-254.2 LO:254.2);ALT=A[chr1:94291257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	94343442	+	chr1	94344635	+	.	35	0	242407_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=242407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:94343442(+)-1:94344635(-)__1_94325001_94350001D;SPAN=1193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:57 GQ:37.4 PL:[100.1, 0.0, 37.4] SR:0 DR:35 LR:-101.6 LO:101.6);ALT=G[chr1:94344635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	94884144	+	chr1	94930329	+	TAAGAAAAGTGGAAAACCACCATTACAGAACAATG	5	5	243066_1	12.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TAAGAAAAGTGGAAAACCACCATTACAGAACAATG;MAPQ=60;MATEID=243066_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_94913001_94938001_22C;SPAN=46185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:26 GQ:12.8 PL:[12.8, 0.0, 49.1] SR:5 DR:5 LR:-12.76 LO:14.02);ALT=G[chr1:94930329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	95699864	+	chr1	95712309	+	.	12	0	244265_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=244265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:95699864(+)-1:95712309(-)__1_95697001_95722001D;SPAN=12445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:56 GQ:24.5 PL:[24.5, 0.0, 110.3] SR:0 DR:12 LR:-24.44 LO:27.6);ALT=C[chr1:95712309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	102821887	-	chr12	106603652	+	.	0	45	5324286_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AATGCAAA;MAPQ=60;MATEID=5324286_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_106599501_106624501_214C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:13 GQ:12 PL:[132.0, 12.0, 0.0] SR:45 DR:0 LR:-132.0 LO:132.0);ALT=[chr12:106603652[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	102892281	+	chr1	102970232	-	.	9	0	254082_1	21.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=254082_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:102892281(+)-1:102970232(+)__1_102949001_102974001D;SPAN=77951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:30 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.58 LO:22.25);ALT=T]chr1:102970232];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	109202586	+	chr1	109203806	+	.	6	5	261900_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=261900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_109196501_109221501_172C;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:5 DR:6 LR:-13.4 LO:17.42);ALT=T[chr1:109203806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109633531	+	chr1	109635510	+	.	18	0	262687_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=262687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109633531(+)-1:109635510(-)__1_109613001_109638001D;SPAN=1979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:48 GQ:46.4 PL:[46.4, 0.0, 69.5] SR:0 DR:18 LR:-46.41 LO:46.68);ALT=G[chr1:109635510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109756677	+	chr1	109770970	+	.	10	0	263007_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=263007_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109756677(+)-1:109770970(-)__1_109760001_109785001D;SPAN=14293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:27 GQ:25.7 PL:[25.7, 0.0, 38.9] SR:0 DR:10 LR:-25.7 LO:25.86);ALT=G[chr1:109770970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109756753	+	chr1	109766600	+	.	0	13	263009_1	35.0	.	EVDNC=ASSMB;HOMSEQ=GTA;MAPQ=60;MATEID=263009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_109760001_109785001_115C;SPAN=9847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:28 GQ:32 PL:[35.3, 0.0, 32.0] SR:13 DR:0 LR:-35.33 LO:35.33);ALT=A[chr1:109766600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109766670	+	chr1	109770972	+	.	0	11	263035_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=263035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_109760001_109785001_167C;SPAN=4302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:11 DR:0 LR:-21.68 LO:25.03);ALT=G[chr1:109770972[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109944714	+	chr1	109953633	+	CAATGTTTGTTGCATTCAGCTTCTCCTCCATTACTTGTTTGAGGATGATGAGTGAAGACTTGATGGCTTCTTTCAAAGTCATAGA	0	30	263221_1	82.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTTG;INSERTION=CAATGTTTGTTGCATTCAGCTTCTCCTCCATTACTTGTTTGAGGATGATGAGTGAAGACTTGATGGCTTCTTTCAAAGTCATAGA;MAPQ=60;MATEID=263221_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_109931501_109956501_178C;SPAN=8919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:63 GQ:68.9 PL:[82.1, 0.0, 68.9] SR:30 DR:0 LR:-82.0 LO:82.0);ALT=T[chr1:109953633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109944714	+	chr1	109952550	+	.	3	23	263220_1	70.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=263220_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_1_109931501_109956501_178C;SPAN=7836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:58 GQ:70.1 PL:[70.1, 0.0, 70.1] SR:23 DR:3 LR:-70.11 LO:70.11);ALT=T[chr1:109952550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109957987	+	chr1	109964482	+	.	12	44	263426_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=263426_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_109956001_109981001_288C;SPAN=6495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:76 GQ:22.4 PL:[161.0, 0.0, 22.4] SR:44 DR:12 LR:-166.9 LO:166.9);ALT=T[chr1:109964482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109958043	+	chr1	109968976	+	.	44	0	263428_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=263428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109958043(+)-1:109968976(-)__1_109956001_109981001D;SPAN=10933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:60 GQ:16.7 PL:[128.9, 0.0, 16.7] SR:0 DR:44 LR:-134.0 LO:134.0);ALT=C[chr1:109968976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	109964601	+	chr1	109968979	+	.	30	0	263441_1	82.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=263441_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:109964601(+)-1:109968979(-)__1_109956001_109981001D;SPAN=4378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:60 GQ:62.9 PL:[82.7, 0.0, 62.9] SR:0 DR:30 LR:-82.92 LO:82.92);ALT=A[chr1:109968979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110091366	+	chr1	110116357	+	.	12	0	263625_1	30.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=263625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110091366(+)-1:110116357(-)__1_110103001_110128001D;SPAN=24991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:0 DR:12 LR:-30.4 LO:30.71);ALT=A[chr1:110116357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110116660	+	chr1	110121826	+	.	2	4	263646_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=263646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_110103001_110128001_103C;SPAN=5166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:59 GQ:2.7 PL:[0.0, 2.7, 148.5] SR:4 DR:2 LR:2.781 LO:7.052);ALT=G[chr1:110121826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	155531853	+	chr1	110191229	+	.	25	0	1738105_1	73.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=1738105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110191229(-)-3:155531853(+)__3_155526001_155551001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:35 GQ:10.4 PL:[73.1, 0.0, 10.4] SR:0 DR:25 LR:-75.56 LO:75.56);ALT=]chr3:155531853]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	110210806	+	chr6	111368654	-	.	12	0	2984549_1	25.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2984549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110210806(+)-6:111368654(+)__6_111352501_111377501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=G]chr6:111368654];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	110230551	+	chr6	111368672	-	.	82	0	2984550_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2984550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110230551(+)-6:111368672(+)__6_111352501_111377501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:47 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=A]chr6:111368672];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	110230551	+	chr1	110231846	+	.	10	0	263617_1	29.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=263617_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110230551(+)-1:110231846(-)__1_110225501_110250501D;SPAN=1295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:3 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:10 LR:-29.71 LO:29.71);ALT=A[chr1:110231846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110944206	+	chr1	110946540	+	.	0	64	265034_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=265034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_110936001_110961001_204C;SPAN=2334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:64 DR:0 LR:-208.0 LO:208.0);ALT=C[chr1:110946540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110944251	+	chr1	110950206	+	.	40	0	265035_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=265035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:110944251(+)-1:110950206(-)__1_110936001_110961001D;SPAN=5955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:74 GQ:65.9 PL:[112.1, 0.0, 65.9] SR:0 DR:40 LR:-112.6 LO:112.6);ALT=C[chr1:110950206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110946658	+	chr1	110950208	+	AATGAAGAATCCCTCCATTGTTGGAGTCCTGTGCACAGATTCACAAGGACTTAATCTGGGTT	61	52	265041_1	99.0	.	DISC_MAPQ=39;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATGAAGAATCCCTCCATTGTTGGAGTCCTGTGCACAGATTCACAAGGACTTAATCTGGGTT;MAPQ=60;MATEID=265041_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_110936001_110961001_85C;SPAN=3550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:79 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:52 DR:61 LR:-290.5 LO:290.5);ALT=C[chr1:110950208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	110949001	+	chr1	110950208	+	.	6	13	265047_1	22.0	.	DISC_MAPQ=29;EVDNC=TSI_L;MAPQ=60;MATEID=265047_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACA;SCTG=c_1_110936001_110961001_85C;SPAN=1207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:13 DR:6 LR:-22.32 LO:28.48);ALT=T[chr1:110950208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111415871	+	chr1	111434012	+	.	37	10	265768_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=265768_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_111426001_111451001_77C;SPAN=18141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:23 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:10 DR:37 LR:-112.2 LO:112.2);ALT=G[chr1:111434012[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111415901	+	chr1	111441744	+	.	17	0	265769_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=265769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111415901(+)-1:111441744(-)__1_111426001_111451001D;SPAN=25843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:35 GQ:36.8 PL:[46.7, 0.0, 36.8] SR:0 DR:17 LR:-46.68 LO:46.68);ALT=C[chr1:111441744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111415908	+	chr1	111434965	+	.	72	0	265771_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=265771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111415908(+)-1:111434965(-)__1_111426001_111451001D;SPAN=19057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:41 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:0 DR:72 LR:-211.3 LO:211.3);ALT=A[chr1:111434965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111435155	+	chr1	111437580	+	TTCTTCATCCTGCTGCTGATTATCCTCCTTGCTGAGGTGACCTTGGCCATCCTGCTCTTTGTATATGAACAGA	3	18	265788_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTCTTCATCCTGCTGCTGATTATCCTCCTTGCTGAGGTGACCTTGGCCATCCTGCTCTTTGTATATGAACAGA;MAPQ=60;MATEID=265788_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_111426001_111451001_29C;SPAN=2425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:78 GQ:48.2 PL:[48.2, 0.0, 140.6] SR:18 DR:3 LR:-48.19 LO:50.73);ALT=G[chr1:111437580[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111437677	+	chr1	111439275	+	.	3	8	265794_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=265794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_111426001_111451001_233C;SPAN=1598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:8 DR:3 LR:-10.42 LO:16.64);ALT=T[chr1:111439275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111990201	+	chr1	111991238	+	.	0	7	266584_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CACCTG;MAPQ=60;MATEID=266584_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_111989501_112014501_216C;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:55 GQ:8.3 PL:[8.3, 0.0, 123.8] SR:7 DR:0 LR:-8.206 LO:14.35);ALT=G[chr1:111991238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111992203	+	chr16	75743669	-	CCCC	30	54	266596_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CCCC;MAPQ=60;MATEID=266596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_111989501_112014501_283C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:28 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:54 DR:30 LR:-181.5 LO:181.5);ALT=G]chr16:75743669];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	111992219	+	chr1	111996831	+	.	83	0	266598_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=266598_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111992219(+)-1:111996831(-)__1_111989501_112014501D;SPAN=4612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:71 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:0 DR:83 LR:-244.3 LO:244.3);ALT=C[chr1:111996831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111992243	+	chr1	111998705	+	.	16	0	266599_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=266599_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:111992243(+)-1:111998705(-)__1_111989501_112014501D;SPAN=6462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:52 GQ:38.9 PL:[38.9, 0.0, 85.1] SR:0 DR:16 LR:-38.73 LO:39.77);ALT=T[chr1:111998705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	111996979	+	chr1	111998706	+	.	0	75	266604_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=266604_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_111989501_112014501_219C;SPAN=1727;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:65 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:75 DR:0 LR:-221.2 LO:221.2);ALT=G[chr1:111998706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112002259	+	chr1	112003535	+	.	10	0	266614_1	16.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=266614_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:112002259(+)-1:112003535(-)__1_111989501_112014501D;SPAN=1276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.48 LO:21.7);ALT=G[chr1:112003535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112016653	+	chr1	112019419	+	GGATGACAGCATGGGAAGCAATGGCTCCACATGTAAACCCGACACT	24	15	266511_1	72.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GGATGACAGCATGGGAAGCAATGGCTCCACATGTAAACCCGACACT;MAPQ=60;MATEID=266511_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_112014001_112039001_212C;SPAN=2766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:75 GQ:72.2 PL:[72.2, 0.0, 108.5] SR:15 DR:24 LR:-72.11 LO:72.54);ALT=G[chr1:112019419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112016653	+	chr1	112018638	+	.	2	4	266510_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=266510_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_112014001_112039001_212C;SPAN=1985;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:4 DR:2 LR:6.574 LO:6.671);ALT=G[chr1:112018638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112016693	+	chr1	112019952	+	.	30	0	266513_1	84.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=266513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:112016693(+)-1:112019952(-)__1_112014001_112039001D;SPAN=3259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:53 GQ:41.9 PL:[84.8, 0.0, 41.9] SR:0 DR:30 LR:-85.37 LO:85.37);ALT=A[chr1:112019952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112162556	+	chr1	112233955	+	.	12	9	266912_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=266912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_112210001_112235001_166C;SPAN=71399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:28 GQ:25.4 PL:[41.9, 0.0, 25.4] SR:9 DR:12 LR:-42.13 LO:42.13);ALT=G[chr1:112233955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112691792	+	chr1	112704704	+	.	68	26	267593_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=267593_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_1_112675501_112700501_71C;SPAN=12912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:7 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:26 DR:68 LR:-241.0 LO:241.0);ALT=G[chr1:112704704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	112835105	+	chr1	112837666	+	.	19	15	267916_1	95.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=AAAAGAGGACACAAACAA;MAPQ=60;MATEID=267916_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_112822501_112847501_136C;SPAN=2561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:26 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:15 DR:19 LR:-95.72 LO:95.72);ALT=A[chr1:112837666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113162537	+	chr1	113197084	+	.	9	0	268504_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=268504_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:113162537(+)-1:113197084(-)__1_113190001_113215001D;SPAN=34547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:21 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.02 LO:24.03);ALT=C[chr1:113197084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113162542	+	chr1	113192038	+	.	9	0	268505_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=268505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:113162542(+)-1:113192038(-)__1_113190001_113215001D;SPAN=29496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:0 DR:9 LR:-23.21 LO:23.34);ALT=G[chr1:113192038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113246430	+	chr1	113247722	+	.	6	7	268626_1	25.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=268626_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_113239001_113264001_110C;SPAN=1292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:65 GQ:25.4 PL:[25.4, 0.0, 131.0] SR:7 DR:6 LR:-25.3 LO:29.46);ALT=T[chr1:113247722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113246472	+	chr1	113249698	+	.	25	0	268627_1	69.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=268627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:113246472(+)-1:113249698(-)__1_113239001_113264001D;SPAN=3226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:47 GQ:43.4 PL:[69.8, 0.0, 43.4] SR:0 DR:25 LR:-70.1 LO:70.1);ALT=G[chr1:113249698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	113317478	+	chr17	4959232	-	.	8	0	6295889_1	17.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6295889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:113317478(+)-17:4959232(+)__17_4949001_4974001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=C]chr17:4959232];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	119401193	+	chr2	141852922	-	TTTTTTTTTTTTTTATTTTTTTTTTTT	18	28	1020923_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TTTTTTTTTTTTTTATTTTTTTTTTTT;MAPQ=60;MATEID=1020923_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_141830501_141855501_322C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:32 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:28 DR:18 LR:-108.9 LO:108.9);ALT=A]chr2:141852922];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr15	44038799	+	chr1	146649791	+	.	36	0	5938554_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5938554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146649791(-)-15:44038799(+)__15_44026501_44051501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:61 GQ:43.1 PL:[102.5, 0.0, 43.1] SR:0 DR:36 LR:-103.5 LO:103.5);ALT=]chr15:44038799]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	146676498	+	chr21	30445877	+	.	74	0	307153_1	99.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=307153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146676498(+)-21:30445877(-)__1_146657001_146682001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:65 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:0 DR:74 LR:-217.9 LO:217.9);ALT=G[chr21:30445877[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	146701616	+	chr1	146818880	-	.	25	0	307685_1	63.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=307685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146701616(+)-1:146818880(+)__1_146804001_146829001D;SPAN=117264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:70 GQ:63.5 PL:[63.5, 0.0, 106.4] SR:0 DR:25 LR:-63.56 LO:64.15);ALT=T]chr1:146818880];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	146702258	-	chr1	146818239	+	.	31	0	307686_1	89.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=307686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146702258(-)-1:146818239(-)__1_146804001_146829001D;SPAN=115981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:48 GQ:26.6 PL:[89.3, 0.0, 26.6] SR:0 DR:31 LR:-91.16 LO:91.16);ALT=[chr1:146818239[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	146714439	+	chr1	146726520	+	.	12	0	307047_1	11.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=307047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146714439(+)-1:146726520(-)__1_146706001_146731001D;SPAN=12081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:106 GQ:11 PL:[11.0, 0.0, 245.3] SR:0 DR:12 LR:-10.89 LO:23.95);ALT=C[chr1:146726520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	146714481	+	chr1	146724276	+	.	12	8	307049_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=307049_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_146706001_146731001_226C;SPAN=9795;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:128 GQ:18.2 PL:[18.2, 0.0, 292.1] SR:8 DR:12 LR:-18.14 LO:32.68);ALT=G[chr1:146724276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	146724390	+	chr1	146726521	+	.	0	11	307086_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=307086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_146706001_146731001_97C;SPAN=2131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:109 GQ:6.8 PL:[6.8, 0.0, 257.6] SR:11 DR:0 LR:-6.78 LO:21.38);ALT=G[chr1:146726521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	146779548	-	chr9	1422886	+	.	17	0	307525_1	42.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=307525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:146779548(-)-9:1422886(-)__1_146779501_146804501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:0 DR:17 LR:-42.84 LO:43.35);ALT=[chr9:1422886[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	150193064	+	chr1	150198939	+	CTCTTCTTCCTCTTCTTCCCCTTCTTCAACATAGTCATCATCATCTTCTTCAT	0	11	321523_1	13.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTCTTCTTCCTCTTCTTCCCCTTCTTCAACATAGTCATCATCATCTTCTTCAT;MAPQ=60;MATEID=321523_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_150185001_150210001_248C;SPAN=5875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:11 DR:0 LR:-13.28 LO:22.64);ALT=C[chr1:150198939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150193064	+	chr1	150195512	+	.	3	6	321522_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=321522_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTTCTT;SCTG=c_1_150185001_150210001_248C;SPAN=2448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:6 PL:[0.0, 6.0, 174.2] SR:6 DR:3 LR:6.44 LO:7.904);ALT=C[chr1:150195512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150199128	+	chr1	150201405	+	.	7	18	321556_1	45.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=321556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150185001_150210001_263C;SPAN=2277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:113 GQ:45.5 PL:[45.5, 0.0, 227.0] SR:18 DR:7 LR:-45.31 LO:52.32);ALT=C[chr1:150201405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150201571	+	chr1	150202906	+	.	0	10	321569_1	8.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=321569_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150185001_150210001_223C;SPAN=1335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:10 DR:0 LR:-8.627 LO:19.88);ALT=C[chr1:150202906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150204266	+	chr1	150208077	+	.	0	13	321583_1	17.0	.	EVDNC=ASSMB;HOMSEQ=TCACCT;MAPQ=60;MATEID=321583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150185001_150210001_260C;SPAN=3811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:95 GQ:17.3 PL:[17.3, 0.0, 212.0] SR:13 DR:0 LR:-17.18 LO:27.1);ALT=T[chr1:150208077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150246573	+	chr1	150248929	+	ATGACTTTAGTGCAGATTTCACCATTGATTACTCCATATTTGAGTCAGAGGACAGGCT	0	13	321656_1	13.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGACTTTAGTGCAGATTTCACCATTGATTACTCCATATTTGAGTCAGAGGACAGGCT;MAPQ=60;MATEID=321656_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_150234001_150259001_230C;SPAN=2356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:108 GQ:13.7 PL:[13.7, 0.0, 248.0] SR:13 DR:0 LR:-13.65 LO:26.32);ALT=G[chr1:150248929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150249040	+	chr1	150252054	+	.	0	9	321671_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=321671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150234001_150259001_379C;SPAN=3014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:108 GQ:0.5 PL:[0.5, 0.0, 261.2] SR:9 DR:0 LR:-0.4492 LO:16.7);ALT=T[chr1:150252054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150266371	+	chr1	150280474	+	.	52	0	321972_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=321972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150266371(+)-1:150280474(-)__1_150258501_150283501D;SPAN=14103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:150 GQ:99 PL:[131.0, 0.0, 233.3] SR:0 DR:52 LR:-131.0 LO:132.6);ALT=A[chr1:150280474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150266869	+	chr1	150280478	+	.	35	51	321977_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ACAG;MAPQ=60;MATEID=321977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150258501_150283501_326C;SPAN=13609;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:134 GQ:86 PL:[237.8, 0.0, 86.0] SR:51 DR:35 LR:-241.5 LO:241.5);ALT=G[chr1:150280478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150600098	+	chr1	150601888	+	.	10	0	323892_1	5.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=323892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150600098(+)-1:150601888(-)__1_150577001_150602001D;SPAN=1790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.918 LO:19.39);ALT=T[chr1:150601888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	83159363	+	chr1	150601553	+	.	9	0	323513_1	9.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=323513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150601553(-)-14:83159363(+)__1_150601501_150626501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=]chr14:83159363]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	150667373	+	chr1	150669527	+	.	10	0	323956_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=323956_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150667373(+)-1:150669527(-)__1_150650501_150675501D;SPAN=2154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=A[chr1:150669527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150702492	+	chr15	83667946	+	.	11	0	6005106_1	32.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=6005106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150702492(+)-15:83667946(-)__15_83643001_83668001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:16 GQ:5.6 PL:[32.0, 0.0, 5.6] SR:0 DR:11 LR:-32.89 LO:32.89);ALT=T[chr15:83667946[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	150705623	+	chr1	150720253	+	.	3	9	324219_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=324219_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150699501_150724501_413C;SPAN=14630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:9 DR:3 LR:-3.158 LO:17.1);ALT=T[chr1:150720253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150722648	+	chr1	150724256	+	.	8	5	324302_1	11.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=324302_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150699501_150724501_349C;SPAN=1608;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:115 GQ:11.9 PL:[11.9, 0.0, 266.0] SR:5 DR:8 LR:-11.76 LO:25.94);ALT=C[chr1:150724256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150724484	+	chr1	150727476	+	.	12	11	324306_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=324306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_150699501_150724501_42C;SPAN=2992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:65 GQ:51.8 PL:[51.8, 0.0, 104.6] SR:11 DR:12 LR:-51.71 LO:52.74);ALT=C[chr1:150727476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150727627	+	chr1	150737114	+	ATGTCTCCCAGGTGGTTCATGCCCAGATCGTATGAGTGCATTCCCATTGAATGCTCCAGGTTGTGAAGCATCACAAACTTTAGATTCTTTTCCCAGATGAGACGTCGTACTGCTTCTTCATT	6	95	324086_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ATGTCTCCCAGGTGGTTCATGCCCAGATCGTATGAGTGCATTCCCATTGAATGCTCCAGGTTGTGAAGCATCACAAACTTTAGATTCTTTTCCCAGATGAGACGTCGTACTGCTTCTTCATT;MAPQ=60;MATEID=324086_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_150724001_150749001_119C;SPAN=9487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:99 DP:144 GQ:60.2 PL:[287.9, 0.0, 60.2] SR:95 DR:6 LR:-296.0 LO:296.0);ALT=C[chr1:150737114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150730458	+	chr1	150737114	+	.	0	71	324107_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=324107_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_1_150724001_150749001_119C;SPAN=6656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:141 GQ:99 PL:[196.4, 0.0, 143.6] SR:71 DR:0 LR:-196.6 LO:196.6);ALT=T[chr1:150737114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150730506	+	chr1	150738173	+	.	66	0	324108_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=324108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150730506(+)-1:150738173(-)__1_150724001_150749001D;SPAN=7667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:91 GQ:25.1 PL:[193.4, 0.0, 25.1] SR:0 DR:66 LR:-200.4 LO:200.4);ALT=A[chr1:150738173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150898995	+	chr1	150900177	+	.	13	0	325134_1	10.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=325134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150898995(+)-1:150900177(-)__1_150895501_150920501D;SPAN=1182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:121 GQ:10.4 PL:[10.4, 0.0, 281.0] SR:0 DR:13 LR:-10.13 LO:25.64);ALT=T[chr1:150900177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150941030	+	chr1	150947092	+	.	8	0	325998_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=325998_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150941030(+)-1:150947092(-)__1_150944501_150969501D;SPAN=6062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:21.5 PL:[21.5, 0.0, 21.5] SR:0 DR:8 LR:-21.53 LO:21.53);ALT=G[chr1:150947092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	150941574	+	chr1	150947093	+	.	20	0	325999_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=325999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:150941574(+)-1:150947093(-)__1_150944501_150969501D;SPAN=5519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:19 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:20 LR:-59.41 LO:59.41);ALT=G[chr1:150947093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151028472	+	chr1	151031954	+	.	44	11	325374_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=325374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151018001_151043001_167C;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:106 GQ:99 PL:[133.1, 0.0, 123.2] SR:11 DR:44 LR:-133.0 LO:133.0);ALT=G[chr1:151031954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151033030	+	chr1	151039693	+	.	9	7	325388_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=325388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151018001_151043001_51C;SPAN=6663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:116 GQ:14.9 PL:[14.9, 0.0, 265.7] SR:7 DR:9 LR:-14.79 LO:28.36);ALT=G[chr1:151039693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151129235	+	chr1	151139407	+	.	22	0	325840_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=325840_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151129235(+)-1:151139407(-)__1_151116001_151141001D;SPAN=10172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:89 GQ:48.5 PL:[48.5, 0.0, 167.3] SR:0 DR:22 LR:-48.51 LO:52.18);ALT=G[chr1:151139407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151129242	+	chr1	151131191	+	.	10	0	325841_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=325841_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151129242(+)-1:151131191(-)__1_151116001_151141001D;SPAN=1949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:0 DR:10 LR:-6.73 LO:19.53);ALT=G[chr1:151131191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151158428	+	chr1	151162480	+	.	0	12	326158_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=326158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151140501_151165501_223C;SPAN=4052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:122 GQ:6.8 PL:[6.8, 0.0, 287.3] SR:12 DR:0 LR:-6.559 LO:23.18);ALT=T[chr1:151162480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151227315	+	chr1	151236388	+	.	12	0	326515_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=326515_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151227315(+)-1:151236388(-)__1_151214001_151239001D;SPAN=9073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:137 GQ:2.6 PL:[2.6, 0.0, 329.3] SR:0 DR:12 LR:-2.495 LO:22.54);ALT=G[chr1:151236388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151227320	+	chr1	151234635	+	.	13	0	326517_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=326517_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151227320(+)-1:151234635(-)__1_151214001_151239001D;SPAN=7315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:117 GQ:11.3 PL:[11.3, 0.0, 272.0] SR:0 DR:13 LR:-11.21 LO:25.84);ALT=G[chr1:151234635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151227321	+	chr10	95719620	-	.	76	0	4663360_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4663360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151227321(+)-10:95719620(+)__10_95697001_95722001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:31 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:0 DR:76 LR:-224.5 LO:224.5);ALT=G]chr10:95719620];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	151867716	+	chr1	151881832	+	.	9	0	329228_1	17.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=329228_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151867716(+)-1:151881832(-)__1_151851001_151876001D;SPAN=14116;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=C[chr1:151881832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151955800	+	chr1	151958579	+	TTCA	0	106	329502_1	99.0	.	EVDNC=ASSMB;INSERTION=TTCA;MAPQ=60;MATEID=329502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151949001_151974001_112C;SPAN=2779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:350 GQ:99 PL:[255.1, 0.0, 595.1] SR:106 DR:0 LR:-255.1 LO:262.6);ALT=T[chr1:151958579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151955849	+	chr1	151966225	+	.	91	0	329503_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=329503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:151955849(+)-1:151966225(-)__1_151949001_151974001D;SPAN=10376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:91 DP:191 GQ:99 PL:[248.9, 0.0, 212.6] SR:0 DR:91 LR:-248.8 LO:248.8);ALT=T[chr1:151966225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	151958729	+	chr1	151966227	+	.	142	17	329512_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=329512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151949001_151974001_205C;SPAN=7498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:151 DP:241 GQ:99 PL:[433.4, 0.0, 149.5] SR:17 DR:142 LR:-440.6 LO:440.6);ALT=T[chr1:151966227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	152005335	+	chr1	152009385	+	.	40	0	329888_1	95.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=329888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:152005335(+)-1:152009385(-)__1_151998001_152023001D;SPAN=4050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:136 GQ:95.3 PL:[95.3, 0.0, 233.9] SR:0 DR:40 LR:-95.2 LO:98.46);ALT=A[chr1:152009385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	152006277	+	chr1	152009388	+	.	120	24	329893_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=329893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_151998001_152023001_209C;SPAN=3111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:141 DP:150 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:24 DR:120 LR:-445.6 LO:445.6);ALT=C[chr1:152009388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153330413	+	chr1	153333117	+	.	10	0	333844_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=333844_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153330413(+)-1:153333117(-)__1_153321001_153346001D;SPAN=2704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:218 GQ:25.9 PL:[0.0, 25.9, 580.9] SR:0 DR:10 LR:26.05 LO:15.89);ALT=C[chr1:153333117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153330909	+	chr1	153333118	+	.	91	147	333846_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=333846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_153321001_153346001_137C;SPAN=2209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:218 DP:315 GQ:99 PL:[634.4, 0.0, 129.4] SR:147 DR:91 LR:-653.0 LO:653.0);ALT=G[chr1:153333118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153346492	+	chr1	153348024	+	.	20	0	333729_1	35.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=333729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153346492(+)-1:153348024(-)__1_153345501_153370501D;SPAN=1532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:112 GQ:35.9 PL:[35.9, 0.0, 233.9] SR:0 DR:20 LR:-35.68 LO:44.22);ALT=G[chr1:153348024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153516400	+	chr1	153518229	+	CCCAAGAAGCTGGGCAGCTCCCGGGTCAGCAGCTCCTTTAGTTCTGACTTGTTGAGCTTGAACTTGTCACCCTCTTTGCCCGAGTACTTGTGGAAGGTGGACACCATCACATCCAGGGCCTTCTCCAGAGGGCACGCCATGACAGCAGTCAGGAT	50	99	334414_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCCAAGAAGCTGGGCAGCTCCCGGGTCAGCAGCTCCTTTAGTTCTGACTTGTTGAGCTTGAACTTGTCACCCTCTTTGCCCGAGTACTTGTGGAAGGTGGACACCATCACATCCAGGGCCTTCTCCAGAGGGCACGCCATGACAGCAGTCAGGAT;MAPQ=60;MATEID=334414_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_153492501_153517501_92C;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:123 DP:340 GQ:99 PL:[313.9, 0.0, 512.0] SR:99 DR:50 LR:-313.9 LO:316.5);ALT=C[chr1:153518229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153632043	+	chr1	153633674	+	.	0	13	334885_1	15.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=334885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_153615001_153640001_367C;SPAN=1631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:100 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:13 DR:0 LR:-15.82 LO:26.79);ALT=G[chr1:153633674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153640603	+	chr1	153643392	+	.	17	0	334926_1	28.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=334926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153640603(+)-1:153643392(-)__1_153639501_153664501D;SPAN=2789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:103 GQ:28.4 PL:[28.4, 0.0, 219.8] SR:0 DR:17 LR:-28.21 LO:36.95);ALT=T[chr1:153643392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153641034	+	chr1	153642645	+	TCAGGCCCTTTGTACCACATATCCCATTTGACTTCTATTT	4	55	334930_1	99.0	.	DISC_MAPQ=52;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TCAGGCCCTTTGTACCACATATCCCATTTGACTTCTATTT;MAPQ=60;MATEID=334930_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_153639501_153664501_375C;SPAN=1611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:117 GQ:99 PL:[156.5, 0.0, 126.8] SR:55 DR:4 LR:-156.6 LO:156.6);ALT=C[chr1:153642645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153641105	+	chr1	153643392	+	.	58	0	334932_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=334932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153641105(+)-1:153643392(-)__1_153639501_153664501D;SPAN=2287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:111 GQ:99 PL:[161.6, 0.0, 105.5] SR:0 DR:58 LR:-161.9 LO:161.9);ALT=C[chr1:153643392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	153947313	+	chr1	153949169	+	TTTGAACTCATTTCTCTTAGATGAGCTGCATGTGATTTTCTCTACATATCCTGTGGGACCACACTCAGGGGTAGTTTT	7	31	336321_1	82.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTTGAACTCATTTCTCTTAGATGAGCTGCATGTGATTTTCTCTACATATCCTGTGGGACCACACTCAGGGGTAGTTTT;MAPQ=60;MATEID=336321_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_153933501_153958501_370C;SPAN=1856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:109 GQ:82.7 PL:[82.7, 0.0, 181.7] SR:31 DR:7 LR:-82.7 LO:84.75);ALT=T[chr1:153949169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56374762	+	chr1	153958676	+	.	32	0	5202764_1	92.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5202764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:153958676(-)-12:56374762(+)__12_56374501_56399501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:47 GQ:20.3 PL:[92.9, 0.0, 20.3] SR:0 DR:32 LR:-95.43 LO:95.43);ALT=]chr12:56374762]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	154130172	+	chr1	154143122	+	.	15	0	337156_1	20.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=337156_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154130172(+)-1:154143122(-)__1_154129501_154154501D;SPAN=12950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:107 GQ:20.6 PL:[20.6, 0.0, 238.4] SR:0 DR:15 LR:-20.53 LO:31.44);ALT=C[chr1:154143122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154145693	+	chr1	154148590	+	.	8	0	337205_1	0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=337205_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154145693(+)-1:154148590(-)__1_154129501_154154501D;SPAN=2897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:115 GQ:4.5 PL:[0.0, 4.5, 287.1] SR:0 DR:8 LR:4.748 LO:14.2);ALT=C[chr1:154148590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154148590	-	chr19	42012395	+	.	13	0	6820991_1	20.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6820991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154148590(-)-19:42012395(-)__19_41993001_42018001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:84 GQ:20.3 PL:[20.3, 0.0, 182.0] SR:0 DR:13 LR:-20.16 LO:27.85);ALT=[chr19:42012395[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	154148745	+	chr1	154155474	+	.	94	0	337633_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=337633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154148745(+)-1:154155474(-)__1_154154001_154179001D;SPAN=6729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:97 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:0 DR:94 LR:-287.2 LO:287.2);ALT=G[chr1:154155474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154187051	+	chr1	154192817	+	.	0	36	337353_1	78.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=337353_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154178501_154203501_251C;SPAN=5766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:149 GQ:78.5 PL:[78.5, 0.0, 283.1] SR:36 DR:0 LR:-78.47 LO:84.97);ALT=C[chr1:154192817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154187052	+	chr1	154192311	+	.	0	7	337354_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=337354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154178501_154203501_195C;SPAN=5259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:124 GQ:10.2 PL:[0.0, 10.2, 320.1] SR:7 DR:0 LR:10.49 LO:11.77);ALT=T[chr1:154192311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154197690	+	chr1	154201091	+	CCACTGCAGAACAAATTAGACTTGCACAGATGATTTCGGACCATAATGATGCTGACTTTGAGGAGAAGGTGAAACAA	3	11	337401_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CCACTGCAGAACAAATTAGACTTGCACAGATGATTTCGGACCATAATGATGCTGACTTTGAGGAGAAGGTGAAACAA;MAPQ=60;MATEID=337401_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_154178501_154203501_320C;SPAN=3401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:11 DR:3 LR:-15.01 LO:26.61);ALT=G[chr1:154201091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154221913	+	chr1	154223516	+	.	2	4	337508_1	0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=337508_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154203001_154228001_29C;SPAN=1603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:101 GQ:10.5 PL:[0.0, 10.5, 264.0] SR:4 DR:2 LR:10.86 LO:8.114);ALT=G[chr1:154223516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154378190	+	chr1	154401671	+	.	4	5	338325_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=338325_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154399001_154424001_187C;SPAN=23481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:52 GQ:9.2 PL:[9.2, 0.0, 114.8] SR:5 DR:4 LR:-9.019 LO:14.54);ALT=G[chr1:154401671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154498415	-	chr1	154499443	+	.	10	0	338695_1	8.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=338695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:154498415(-)-1:154499443(-)__1_154497001_154522001D;SPAN=1028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:0 DR:10 LR:-8.085 LO:19.77);ALT=[chr1:154499443[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	154575106	+	chr1	154580467	+	.	0	14	339196_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CCTGC;MAPQ=60;MATEID=339196_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_154570501_154595501_6C;SPAN=5361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:117 GQ:14.6 PL:[14.6, 0.0, 268.7] SR:14 DR:0 LR:-14.52 LO:28.31);ALT=C[chr1:154580467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154897743	+	chr1	154898829	+	.	3	4	340402_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=340402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154889001_154914001_264C;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:122 GQ:16.2 PL:[0.0, 16.2, 326.7] SR:4 DR:3 LR:16.55 LO:7.697);ALT=T[chr1:154898829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154898960	+	chr1	154901500	+	.	3	7	340406_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=340406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_154889001_154914001_89C;SPAN=2540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:7 DR:3 LR:6.374 LO:14.01);ALT=C[chr1:154901500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154901655	+	chr1	154909067	+	AGCATACTGTTCCTTGAGTGGACCAGAGAGCCGGAGGACAGCACAGACATCAGCTCCAAGT	25	28	340424_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTGC;INSERTION=AGCATACTGTTCCTTGAGTGGACCAGAGAGCCGGAGGACAGCACAGACATCAGCTCCAAGT;MAPQ=60;MATEID=340424_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_154889001_154914001_395C;SPAN=7412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:123 GQ:99 PL:[105.5, 0.0, 191.3] SR:28 DR:25 LR:-105.3 LO:106.7);ALT=G[chr1:154909067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	154904895	+	chr1	154909067	+	.	12	16	340435_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTGC;MAPQ=60;MATEID=340435_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_154889001_154914001_395C;SPAN=4172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:120 GQ:30.2 PL:[30.2, 0.0, 261.2] SR:16 DR:12 LR:-30.21 LO:40.92);ALT=C[chr1:154909067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155023944	+	chr1	155025145	+	.	0	12	340785_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AGGTG;MAPQ=60;MATEID=340785_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155011501_155036501_407C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:109 GQ:10.1 PL:[10.1, 0.0, 254.3] SR:12 DR:0 LR:-10.08 LO:23.8);ALT=G[chr1:155025145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155025253	+	chr1	155026384	+	ACCAGTCTGCCTGAGCCCCTGAGGATCAAGTTGGAGCTGGACGGTGACAGTCATATCCTGGAGCTGCTACAGAAT	0	29	340790_1	63.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ACCAGTCTGCCTGAGCCCCTGAGGATCAAGTTGGAGCTGGACGGTGACAGTCATATCCTGGAGCTGCTACAGAAT;MAPQ=60;MATEID=340790_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_155011501_155036501_329C;SPAN=1131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:121 GQ:63.2 PL:[63.2, 0.0, 228.2] SR:29 DR:0 LR:-62.95 LO:68.33);ALT=G[chr1:155026384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155108507	+	chr1	155110034	+	.	17	0	341199_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=341199_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155108507(+)-1:155110034(-)__1_155085001_155110001D;SPAN=1527;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:87 GQ:32.6 PL:[32.6, 0.0, 177.8] SR:0 DR:17 LR:-32.55 LO:38.33);ALT=G[chr1:155110034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155108852	+	chr1	155110037	+	.	2	15	341202_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=341202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155085001_155110001_212C;SPAN=1185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:90 GQ:31.7 PL:[31.7, 0.0, 186.8] SR:15 DR:2 LR:-31.73 LO:38.05);ALT=A[chr1:155110037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155108858	+	chr1	155110453	+	.	11	0	341203_1	19.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=341203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155108858(+)-1:155110453(-)__1_155085001_155110001D;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:64 GQ:19.1 PL:[19.1, 0.0, 134.6] SR:0 DR:11 LR:-18.97 LO:24.12);ALT=G[chr1:155110453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155145213	-	chr2	45223753	+	.	29	0	341394_1	67.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=341394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155145213(-)-2:45223753(-)__1_155134001_155159001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:105 GQ:67.4 PL:[67.4, 0.0, 186.2] SR:0 DR:29 LR:-67.28 LO:70.43);ALT=[chr2:45223753[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	155145423	+	chr1	155151247	+	.	17	0	341396_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=341396_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155145423(+)-1:155151247(-)__1_155134001_155159001D;SPAN=5824;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:108 GQ:26.9 PL:[26.9, 0.0, 234.8] SR:0 DR:17 LR:-26.86 LO:36.56);ALT=G[chr1:155151247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155145951	+	chr1	155151248	+	.	49	13	341400_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=341400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155134001_155159001_20C;SPAN=5297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:82 GQ:47.3 PL:[149.6, 0.0, 47.3] SR:13 DR:49 LR:-152.2 LO:152.2);ALT=C[chr1:155151248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155230453	+	chr1	155231877	+	.	12	7	341797_1	49.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=341797_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155232001_155257001_255C;SPAN=1424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:0 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:7 DR:12 LR:-49.51 LO:49.51);ALT=G[chr1:155231877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155278788	+	chr1	155282043	+	.	17	0	341886_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=341886_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155278788(+)-1:155282043(-)__1_155281001_155306001D;SPAN=3255;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:58 GQ:40.4 PL:[40.4, 0.0, 99.8] SR:0 DR:17 LR:-40.4 LO:41.81);ALT=A[chr1:155282043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155279998	+	chr1	155282044	+	.	6	10	341887_1	36.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=0;MATEID=341887_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155281001_155306001_17C;SECONDARY;SPAN=2046;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:10 DR:6 LR:-36.83 LO:38.71);ALT=T[chr1:155282044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155658965	+	chr1	155679563	+	.	11	2	343833_1	24.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=343833_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_1_155648501_155673501_166C;SPAN=20598;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:2 DR:11 LR:-24.71 LO:27.71);ALT=G[chr1:155679563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155658973	+	chr1	155686794	+	.	35	0	343834_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=343834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155658973(+)-1:155686794(-)__1_155648501_155673501D;SPAN=27821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:54 GQ:28.4 PL:[101.0, 0.0, 28.4] SR:0 DR:35 LR:-103.0 LO:103.0);ALT=A[chr1:155686794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155658982	+	chr1	155691305	+	.	12	0	343835_1	25.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=343835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155658982(+)-1:155691305(-)__1_155648501_155673501D;SPAN=32323;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=A[chr1:155691305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155686920	+	chr1	155691307	+	.	0	17	343710_1	26.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=343710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155673001_155698001_356C;SPAN=4387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:112 GQ:26 PL:[26.0, 0.0, 243.8] SR:17 DR:0 LR:-25.77 LO:36.27);ALT=G[chr1:155691307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155823604	+	chr1	155826937	+	.	26	0	344526_1	56.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=344526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155823604(+)-1:155826937(-)__1_155820001_155845001D;SPAN=3333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:111 GQ:56 PL:[56.0, 0.0, 211.1] SR:0 DR:26 LR:-55.75 LO:60.96);ALT=G[chr1:155826937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155898178	-	chr1	155899748	+	.	10	0	344765_1	4.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=344765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155898178(-)-1:155899748(-)__1_155893501_155918501D;SPAN=1570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:0 DR:10 LR:-4.292 LO:19.12);ALT=[chr1:155899748[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	155939093	+	chr1	155948156	+	.	0	10	345407_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=345407_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155918001_155943001_256C;SPAN=9063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:66 GQ:15.2 PL:[15.2, 0.0, 143.9] SR:10 DR:0 LR:-15.13 LO:21.33);ALT=T[chr1:155948156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155979441	+	chr1	155981601	+	.	6	8	345703_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=345703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155967001_155992001_24C;SPAN=2160;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:121 GQ:13.7 PL:[13.7, 0.0, 277.7] SR:8 DR:6 LR:-13.43 LO:28.09);ALT=G[chr1:155981601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155981679	+	chr1	155984752	+	.	3	15	345720_1	24.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=345720_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_155967001_155992001_266C;SPAN=3073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:118 GQ:24.2 PL:[24.2, 0.0, 261.8] SR:15 DR:3 LR:-24.15 LO:35.85);ALT=C[chr1:155984752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155981679	+	chr1	155988061	+	ACAACGGGCCCATCCTCCTGGGCCAGGTAAGTAATTGTTGCCGAGGTGAAGTTGAAATAACCAGCCTTGAGAGGGCGCAGGACCACAGTGTGGGAGACATTGCTAGCA	0	87	345721_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ACAACGGGCCCATCCTCCTGGGCCAGGTAAGTAATTGTTGCCGAGGTGAAGTTGAAATAACCAGCCTTGAGAGGGCGCAGGACCACAGTGTGGGAGACATTGCTAGCA;MAPQ=60;MATEID=345721_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_155967001_155992001_266C;SPAN=6382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:145 GQ:99 PL:[248.0, 0.0, 102.8] SR:87 DR:0 LR:-251.1 LO:251.1);ALT=C[chr1:155988061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155984907	+	chr1	155990678	+	.	33	0	345740_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=345740_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155984907(+)-1:155990678(-)__1_155967001_155992001D;SPAN=5771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:149 GQ:68.6 PL:[68.6, 0.0, 293.0] SR:0 DR:33 LR:-68.57 LO:76.45);ALT=G[chr1:155990678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155988161	+	chr1	155989804	+	.	0	104	345758_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=345758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_155967001_155992001_344C;SPAN=1643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:104 DP:175 GQ:99 PL:[296.0, 0.0, 127.7] SR:104 DR:0 LR:-299.5 LO:299.5);ALT=T[chr1:155989804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	155988214	+	chr1	155990676	+	.	93	0	345760_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=345760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:155988214(+)-1:155990676(-)__1_155967001_155992001D;SPAN=2462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:93 DP:145 GQ:83 PL:[267.8, 0.0, 83.0] SR:0 DR:93 LR:-273.0 LO:273.0);ALT=C[chr1:155990676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156024751	+	chr1	156027767	+	.	17	0	345464_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=345464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156024751(+)-1:156027767(-)__1_156016001_156041001D;SPAN=3016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:138 GQ:18.8 PL:[18.8, 0.0, 315.8] SR:0 DR:17 LR:-18.73 LO:34.6);ALT=G[chr1:156027767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156025217	+	chr1	156028104	+	AGGGCCGTGTAGCCATCACCCGAGTGGCCAACCTTCTGCTGTGTATGTATGCCAAGGAGACCGTGGGCTTTGGAATGCTCAAGGCCA	3	158	345469_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AGGGCCGTGTAGCCATCACCCGAGTGGCCAACCTTCTGCTGTGTATGTATGCCAAGGAGACCGTGGGCTTTGGAATGCTCAAGGCCA;MAPQ=60;MATEID=345469_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_156016001_156041001_265C;SPAN=2887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:160 DP:158 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:158 DR:3 LR:-475.3 LO:475.3);ALT=G[chr1:156028104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156085065	+	chr1	156100407	+	.	0	7	345778_1	7.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=345778_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156089501_156114501_161C;SPAN=15342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:58 GQ:7.4 PL:[7.4, 0.0, 132.8] SR:7 DR:0 LR:-7.393 LO:14.18);ALT=G[chr1:156100407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156100564	+	chr1	156104192	+	.	8	8	345821_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=345821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156089501_156114501_135C;SPAN=3628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:117 GQ:11.3 PL:[11.3, 0.0, 272.0] SR:8 DR:8 LR:-11.21 LO:25.84);ALT=G[chr1:156104192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156146525	-	chr1	156148110	+	.	8	0	346271_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=346271_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156146525(-)-1:156148110(-)__1_156138501_156163501D;SPAN=1585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:119 GQ:5.7 PL:[0.0, 5.7, 300.3] SR:0 DR:8 LR:5.832 LO:14.07);ALT=[chr1:156148110[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	156182881	+	chr1	156203417	+	.	11	0	346572_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=346572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156182881(+)-1:156203417(-)__1_156187501_156212501D;SPAN=20536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:53 GQ:22.1 PL:[22.1, 0.0, 104.6] SR:0 DR:11 LR:-21.95 LO:25.13);ALT=T[chr1:156203417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156182967	+	chr1	156202108	+	.	0	36	346212_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=346212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156163001_156188001_434C;SPAN=19141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:66 GQ:58.1 PL:[101.0, 0.0, 58.1] SR:36 DR:0 LR:-101.5 LO:101.5);ALT=G[chr1:156202108[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156202217	+	chr1	156203418	+	.	0	19	346629_1	26.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=346629_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_156187501_156212501_336C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:135 GQ:26.3 PL:[26.3, 0.0, 300.2] SR:19 DR:0 LR:-26.14 LO:39.86);ALT=G[chr1:156203418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156203520	+	chr1	156206078	+	.	3	6	346640_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=346640_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_156187501_156212501_80C;SPAN=2558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:124 GQ:6.9 PL:[0.0, 6.9, 313.5] SR:6 DR:3 LR:7.187 LO:13.93);ALT=G[chr1:156206078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156206275	+	chr1	156209336	+	.	6	2	346655_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=346655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156187501_156212501_45C;SPAN=3061;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:120 GQ:9.3 PL:[0.0, 9.3, 310.2] SR:2 DR:6 LR:9.404 LO:11.87);ALT=G[chr1:156209336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156248826	+	chr1	156252397	+	.	0	7	346528_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=346528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156236501_156261501_322C;SPAN=3571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:124 GQ:10.2 PL:[0.0, 10.2, 320.1] SR:7 DR:0 LR:10.49 LO:11.77);ALT=C[chr1:156252397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156252821	+	chr1	156254970	+	.	8	0	346547_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=346547_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156252821(+)-1:156254970(-)__1_156236501_156261501D;SPAN=2149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=C[chr1:156254970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156279096	+	chr1	156280349	+	.	0	10	346435_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=346435_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156261001_156286001_11C;SPAN=1253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:103 GQ:5.3 PL:[5.3, 0.0, 242.9] SR:10 DR:0 LR:-5.105 LO:19.26);ALT=T[chr1:156280349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156287040	+	chr1	156288659	+	GAGATGCCCTTTTCAGTGATGACCACATCGGGCTTCAGTTGGATAATGTCCTCACAGAGCTGCTGGATGTACTCTTCCTCCATCTGGAGAATTCGGGTGAAGTCCTCCTCTCGTGTAATCTCAATGTCAGT	2	10	346783_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GAGATGCCCTTTTCAGTGATGACCACATCGGGCTTCAGTTGGATAATGTCCTCACAGAGCTGCTGGATGTACTCTTCCTCCATCTGGAGAATTCGGGTGAAGTCCTCCTCTCGTGTAATCTCAATGTCAGT;MAPQ=60;MATEID=346783_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_156285501_156310501_198C;SPAN=1619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:107 GQ:4.1 PL:[4.1, 0.0, 254.9] SR:10 DR:2 LR:-4.021 LO:19.08);ALT=T[chr1:156288659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156287341	+	chr1	156288659	+	.	3	6	346785_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=346785_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_156285501_156310501_198C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:6 DR:3 LR:-1.804 LO:16.9);ALT=G[chr1:156288659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156294881	+	chr1	156307944	+	AAGAATAATTACTGATGTGGTCCCATCTCCAACCTCTTCATCCTGGGTCCGGCTAATTTCGATCATGGACTTGGCCGCTGGATGCTGGACTTGAATCTCTCGAAGAATGGCATTGCCATCATTGGTCATCACAATGCCTCCCATTGGGTCCAAAAGCATCTTCATCATGGACTTGGGTCCCAAACATGTTCGGATGATATCTGCAATAGTCTTGGCAGCATTGATGTTTCCAGATTGAACTTTTCTTCCGGATTCACGCTTTGTGTTCTGG	0	32	346826_1	70.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AAGAATAATTACTGATGTGGTCCCATCTCCAACCTCTTCATCCTGGGTCCGGCTAATTTCGATCATGGACTTGGCCGCTGGATGCTGGACTTGAATCTCTCGAAGAATGGCATTGCCATCATTGGTCATCACAATGCCTCCCATTGGGTCCAAAAGCATCTTCATCATGGACTTGGGTCCCAAACATGTTCGGATGATATCTGCAATAGTCTTGGCAGCATTGATGTTTCCAGATTGAACTTTTCTTCCGGATTCACGCTTTGTGTTCTGG;MAPQ=60;MATEID=346826_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_1_156285501_156310501_160C;SPAN=13063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:129 GQ:70.7 PL:[70.7, 0.0, 242.3] SR:32 DR:0 LR:-70.68 LO:75.96);ALT=C[chr1:156307944[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156303489	+	chr1	156307943	+	.	24	0	346871_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=346871_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156303489(+)-1:156307943(-)__1_156285501_156310501D;SPAN=4454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:115 GQ:48.2 PL:[48.2, 0.0, 229.7] SR:0 DR:24 LR:-48.07 LO:54.89);ALT=G[chr1:156307943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156304760	+	chr1	156307943	+	.	57	0	346887_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=346887_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156304760(+)-1:156307943(-)__1_156285501_156310501D;SPAN=3183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:134 GQ:99 PL:[152.0, 0.0, 171.8] SR:0 DR:57 LR:-151.9 LO:151.9);ALT=G[chr1:156307943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156305679	+	chr1	156307944	+	.	22	13	346890_1	48.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=346890_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_1_156285501_156310501_160C;SPAN=2265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:137 GQ:48.8 PL:[48.8, 0.0, 283.1] SR:13 DR:22 LR:-48.71 LO:58.26);ALT=C[chr1:156307944[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156526723	+	chr1	156528936	+	.	110	73	347636_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGAAATTGAGTAGCTCAGC;MAPQ=60;MATEID=347636_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_1_156506001_156531001_299C;SPAN=2213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:48 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:73 DR:110 LR:-432.4 LO:432.4);ALT=C[chr1:156528936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156568334	+	chr1	156571199	+	.	13	0	347930_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=347930_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156568334(+)-1:156571199(-)__1_156555001_156580001D;SPAN=2865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:140 GQ:5 PL:[5.0, 0.0, 335.0] SR:0 DR:13 LR:-4.984 LO:24.77);ALT=G[chr1:156571199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156568939	+	chr1	156571200	+	.	10	0	347933_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=347933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156568939(+)-1:156571200(-)__1_156555001_156580001D;SPAN=2261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:116 GQ:1.7 PL:[1.7, 0.0, 278.9] SR:0 DR:10 LR:-1.583 LO:18.71);ALT=C[chr1:156571200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	156705398	+	chr14	61033233	+	.	12	0	348886_1	32.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=348886_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:156705398(+)-14:61033233(-)__1_156702001_156727001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:25 GQ:26.3 PL:[32.9, 0.0, 26.3] SR:0 DR:12 LR:-32.86 LO:32.86);ALT=A[chr14:61033233[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	156708559	+	chr1	156710804	+	.	73	2	348902_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=348902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_156702001_156727001_150C;SPAN=2245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:122 GQ:86 PL:[208.1, 0.0, 86.0] SR:2 DR:73 LR:-210.6 LO:210.6);ALT=G[chr1:156710804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	157030415	+	chr9	33076580	+	.	9	0	4172766_1	12.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=4172766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:157030415(+)-9:33076580(-)__9_33075001_33100001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:63 GQ:12.8 PL:[12.8, 0.0, 138.2] SR:0 DR:9 LR:-12.64 LO:18.94);ALT=G[chr9:33076580[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	157279009	+	chr10	130774980	-	.	4	29	4719234_1	89.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=4719234_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_130756501_130781501_220C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:24 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:29 DR:4 LR:-89.12 LO:89.12);ALT=T]chr10:130774980];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	157348495	+	chr1	157457782	-	.	31	0	350898_1	89.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=350898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:157348495(+)-1:157457782(+)__1_157437001_157462001D;SPAN=109287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:27 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=T]chr1:157457782];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	158801348	+	chr1	158811922	+	.	22	22	354864_1	94.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=354864_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_158784501_158809501_109C;SPAN=10574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:43 GQ:8.3 PL:[94.1, 0.0, 8.3] SR:22 DR:22 LR:-97.88 LO:97.88);ALT=G[chr1:158811922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	158815827	+	chr1	158817514	+	.	8	0	354754_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=354754_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:158815827(+)-1:158817514(-)__1_158809001_158834001D;SPAN=1687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=C[chr1:158817514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	158961355	+	chr1	158966212	+	CATGGT	129	74	355055_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=CATGGT;MAPQ=60;MATEID=355055_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_158956001_158981001_36C;SPAN=4857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:166 DP:55 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:74 DR:129 LR:-491.8 LO:491.8);ALT=G[chr1:158966212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	158979850	+	chr1	158984448	+	.	10	0	355474_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=355474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:158979850(+)-1:158984448(-)__1_158980501_159005501D;SPAN=4598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.48 LO:21.7);ALT=G[chr1:158984448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	158990319	+	chr1	159002311	+	.	5	4	355526_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=355526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_158980501_159005501_342C;SPAN=11992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:109 GQ:9.6 PL:[0.0, 9.6, 283.8] SR:4 DR:5 LR:9.725 LO:10.02);ALT=G[chr1:159002311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159023516	+	chr1	159024606	+	.	3	4	355315_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAAGGT;MAPQ=60;MATEID=355315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_159005001_159030001_163C;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:100 GQ:7.2 PL:[0.0, 7.2, 257.4] SR:4 DR:3 LR:7.287 LO:10.25);ALT=T[chr1:159024606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159272222	+	chr1	159273715	+	.	8	0	356130_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=356130_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159272222(+)-1:159273715(-)__1_159250001_159275001D;SPAN=1493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=T[chr1:159273715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159428659	+	chr1	159494970	-	.	8	0	356742_1	10.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=356742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159428659(+)-1:159494970(+)__1_159421501_159446501D;SPAN=66311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:0 DR:8 LR:-10.69 LO:16.71);ALT=C]chr1:159494970];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr1	159888618	+	chr1	159895238	+	.	8	0	358325_1	0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=358325_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159888618(+)-1:159895238(-)__1_159887001_159912001D;SPAN=6620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:396 GQ:80.6 PL:[0.0, 80.6, 1122.0] SR:0 DR:8 LR:80.88 LO:9.856);ALT=C[chr1:159895238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159889673	+	chr1	159895237	+	.	92	0	358330_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=358330_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159889673(+)-1:159895237(-)__1_159887001_159912001D;SPAN=5564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:304 GQ:99 PL:[221.5, 0.0, 515.3] SR:0 DR:92 LR:-221.3 LO:227.8);ALT=C[chr1:159895237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	159890358	+	chr1	159895237	+	.	112	0	358338_1	99.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=358338_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:159890358(+)-1:159895237(-)__1_159887001_159912001D;SPAN=4879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:295 GQ:99 PL:[289.9, 0.0, 425.3] SR:0 DR:112 LR:-289.8 LO:291.2);ALT=C[chr1:159895237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	160175312	+	chr1	160181332	+	.	17	8	359131_1	47.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=359131_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_160181001_160206001_24C;SPAN=6020;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:68 GQ:47.6 PL:[47.6, 0.0, 116.9] SR:8 DR:17 LR:-47.6 LO:49.23);ALT=G[chr1:160181332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	160253450	+	chr1	160254861	+	.	8	0	359126_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=359126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:160253450(+)-1:160254861(-)__1_160230001_160255001D;SPAN=1411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:108 GQ:2.7 PL:[0.0, 2.7, 267.3] SR:0 DR:8 LR:2.852 LO:14.42);ALT=G[chr1:160254861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	160314616	+	chr1	160318789	+	.	2	7	359661_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=359661_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_160303501_160328501_274C;SPAN=4173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:99 GQ:2.9 PL:[2.9, 0.0, 237.2] SR:7 DR:2 LR:-2.887 LO:17.06);ALT=T[chr1:160318789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	160654981	+	chr1	160681470	+	.	15	6	361269_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=361269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_160646501_160671501_384C;SPAN=26489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:6 DR:15 LR:-39.0 LO:39.93);ALT=T[chr1:160681470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	21958921	+	chr1	160864770	+	.	36	0	361704_1	99.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=361704_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:160864770(-)-23:21958921(+)__1_160842501_160867501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:70 GQ:70.1 PL:[99.8, 0.0, 70.1] SR:0 DR:36 LR:-100.2 LO:100.2);ALT=]chrX:21958921]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	160970917	+	chr1	160990799	+	GATTATTCTCAGGAATTCTGACTTCAGGTTCAGAAGAGTGCACTGTAACACTGCCCAATGCCAGGGAG	17	23	362433_1	73.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GATTATTCTCAGGAATTCTGACTTCAGGTTCAGAAGAGTGCACTGTAACACTGCCCAATGCCAGGGAG;MAPQ=60;MATEID=362433_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_160989501_161014501_13C;SPAN=19882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:45 GQ:34.1 PL:[73.7, 0.0, 34.1] SR:23 DR:17 LR:-74.35 LO:74.35);ALT=G[chr1:160990799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161013186	+	chr1	161015705	+	.	8	0	362549_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=362549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161013186(+)-1:161015705(-)__1_160989501_161014501D;SPAN=2519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=A[chr1:161015705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161070651	+	chr1	161071838	+	.	3	40	362598_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=362598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161063001_161088001_288C;SPAN=1187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:129 GQ:99 PL:[103.7, 0.0, 209.3] SR:40 DR:3 LR:-103.7 LO:105.7);ALT=T[chr1:161071838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161070700	+	chr1	161087762	+	.	15	0	362600_1	17.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=362600_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161070700(+)-1:161087762(-)__1_161063001_161088001D;SPAN=17062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:118 GQ:17.6 PL:[17.6, 0.0, 268.4] SR:0 DR:15 LR:-17.55 LO:30.75);ALT=C[chr1:161087762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161072167	+	chr1	161087738	+	.	142	20	362607_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCACCT;MAPQ=60;MATEID=362607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161063001_161088001_274C;SPAN=15571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:113 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:20 DR:142 LR:-448.9 LO:448.9);ALT=T[chr1:161087738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161094374	+	chr1	161102339	+	.	19	0	362368_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=362368_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161094374(+)-1:161102339(-)__1_161087501_161112501D;SPAN=7965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:120 GQ:30.2 PL:[30.2, 0.0, 261.2] SR:0 DR:19 LR:-30.21 LO:40.92);ALT=A[chr1:161102339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161123910	+	chr1	161126739	+	.	46	60	362922_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=362922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161112001_161137001_325C;SPAN=2829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:84 DP:132 GQ:76.7 PL:[241.7, 0.0, 76.7] SR:60 DR:46 LR:-246.1 LO:246.1);ALT=G[chr1:161126739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161123929	+	chr1	161127042	+	.	40	0	362924_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=362924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161123929(+)-1:161127042(-)__1_161112001_161137001D;SPAN=3113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:137 GQ:95 PL:[95.0, 0.0, 236.9] SR:0 DR:40 LR:-94.92 LO:98.31);ALT=G[chr1:161127042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161123944	+	chr1	161127405	+	.	27	0	362926_1	52.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=362926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161123944(+)-1:161127405(-)__1_161112001_161137001D;SPAN=3461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:137 GQ:52.1 PL:[52.1, 0.0, 279.8] SR:0 DR:27 LR:-52.01 LO:61.0);ALT=T[chr1:161127405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161172305	+	chr1	161176195	+	.	35	0	362703_1	86.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=362703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161172305(+)-1:161176195(-)__1_161161001_161186001D;SPAN=3890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:109 GQ:86 PL:[86.0, 0.0, 178.4] SR:0 DR:35 LR:-86.01 LO:87.78);ALT=C[chr1:161176195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161173333	+	chr1	161176196	+	.	0	42	362708_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=362708_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_1_161161001_161186001_231C;SPAN=2863;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:114 GQ:99 PL:[107.9, 0.0, 167.3] SR:42 DR:0 LR:-107.8 LO:108.5);ALT=G[chr1:161176196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161185160	+	chr1	161187773	+	.	38	2	362759_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=362759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_161161001_161186001_355C;SPAN=2613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:2 DR:38 LR:-120.9 LO:120.9);ALT=G[chr1:161187773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161284254	+	chr1	161298185	+	.	14	0	363668_1	15.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=363668_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161284254(+)-1:161298185(-)__1_161283501_161308501D;SPAN=13931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:115 GQ:15.2 PL:[15.2, 0.0, 262.7] SR:0 DR:14 LR:-15.06 LO:28.42);ALT=T[chr1:161298185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	161298185	-	chr17	1761687	+	.	18	0	6284008_1	43.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=6284008_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:161298185(-)-17:1761687(-)__17_1739501_1764501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:60 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:0 DR:18 LR:-43.16 LO:44.49);ALT=[chr17:1761687[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	161748111	+	chr1	161751702	+	.	0	10	366040_1	20.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=366040_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_161724501_161749501_302C;SPAN=3591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:10 DR:0 LR:-20.82 LO:23.18);ALT=G[chr1:161751702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	190999445	+	chr1	164240436	+	.	28	45	1134641_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1134641_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_190977501_191002501_91C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:27 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:45 DR:28 LR:-181.5 LO:181.5);ALT=]chr2:190999445]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	164240562	+	chr2	190999443	+	TTAAAACACATTTCC	28	34	1134642_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TTAAAACACATTTCC;MAPQ=60;MATEID=1134642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_190977501_191002501_209C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:27 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:34 DR:28 LR:-148.5 LO:148.5);ALT=A[chr2:190999443[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	165600530	+	chr1	165619075	+	.	52	14	379424_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=379424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165595501_165620501_23C;SPAN=18545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:161 GQ:99 PL:[138.2, 0.0, 250.4] SR:14 DR:52 LR:-137.9 LO:139.8);ALT=G[chr1:165619075[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600565	+	chr1	165623513	+	.	12	0	379506_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=379506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:165600565(+)-1:165623513(-)__1_165620001_165645001D;SPAN=22948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:0 DR:12 LR:-23.36 LO:27.2);ALT=C[chr1:165623513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600578	+	chr1	165621212	+	.	41	0	379508_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=379508_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:165600578(+)-1:165621212(-)__1_165620001_165645001D;SPAN=20634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:61 GQ:26.6 PL:[119.0, 0.0, 26.6] SR:0 DR:41 LR:-121.8 LO:121.8);ALT=G[chr1:165621212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165600581	+	chr1	165620247	+	.	90	0	379509_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=379509_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:165600581(+)-1:165620247(-)__1_165620001_165645001D;SPAN=19666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:88 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:0 DR:90 LR:-267.4 LO:267.4);ALT=C[chr1:165620247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165619201	+	chr1	165620249	+	.	8	109	379500_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=379500_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165595501_165620501_107C;SPAN=1048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:114 DP:175 GQ:94.7 PL:[329.0, 0.0, 94.7] SR:109 DR:8 LR:-336.0 LO:336.0);ALT=G[chr1:165620249[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165623588	+	chr1	165624603	+	.	0	59	379530_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=379530_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165620001_165645001_268C;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:143 GQ:99 PL:[156.2, 0.0, 189.2] SR:59 DR:0 LR:-156.0 LO:156.2);ALT=G[chr1:165624603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165664635	+	chr1	165667614	+	.	0	8	380093_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=380093_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165644501_165669501_390C;SPAN=2979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:8 DR:0 LR:-0.9411 LO:14.92);ALT=C[chr1:165667614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165697362	+	chr1	165712404	+	.	4	8	379706_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGT;MAPQ=60;MATEID=379706_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165693501_165718501_16C;SPAN=15042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:114 GQ:5.6 PL:[5.6, 0.0, 269.6] SR:8 DR:4 LR:-5.426 LO:21.15);ALT=T[chr1:165712404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165712548	+	chr1	165721339	+	.	3	9	379805_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=379805_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165718001_165743001_298C;SPAN=8791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:46 GQ:27.2 PL:[27.2, 0.0, 83.3] SR:9 DR:3 LR:-27.15 LO:28.79);ALT=T[chr1:165721339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165723513	+	chr1	165737918	+	ATTTTCTTTTTCTGTTGTCGACCAGCTGACTCTGTTATTGTTTCCTTCTTCTTTTCCAATTTTTTACTCTGTTTTTCCACTTCTGCCTTCAGTCTCTTGTACTTGTCTGTCCTGTAAACCAGGACCCAGGTTATG	5	43	379828_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=ATTTTCTTTTTCTGTTGTCGACCAGCTGACTCTGTTATTGTTTCCTTCTTCTTTTCCAATTTTTTACTCTGTTTTTCCACTTCTGCCTTCAGTCTCTTGTACTTGTCTGTCCTGTAAACCAGGACCCAGGTTATG;MAPQ=60;MATEID=379828_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_1_165718001_165743001_187C;SPAN=14405;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:117 GQ:99 PL:[113.6, 0.0, 169.7] SR:43 DR:5 LR:-113.5 LO:114.2);ALT=T[chr1:165737918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	165797169	+	chr1	165859439	+	.	14	5	381077_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=381077_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_165840501_165865501_142C;SPAN=62270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:52 GQ:35.6 PL:[35.6, 0.0, 88.4] SR:5 DR:14 LR:-35.43 LO:36.77);ALT=G[chr1:165859439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	166246845	+	chr22	29664367	-	.	10	0	7258364_1	19.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=7258364_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:166246845(+)-22:29664367(+)__22_29645001_29670001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=T]chr22:29664367];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	167511538	+	chr1	167515336	+	.	6	12	385859_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=385859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167506501_167531501_6C;SPAN=3798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:87 GQ:32.6 PL:[32.6, 0.0, 177.8] SR:12 DR:6 LR:-32.55 LO:38.33);ALT=C[chr1:167515336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167515524	+	chr1	167517237	+	.	3	9	385878_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=385878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167506501_167531501_323C;SPAN=1713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:9 DR:3 LR:-10.84 LO:22.13);ALT=T[chr1:167517237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167517360	+	chr1	167522624	+	.	2	7	385891_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=385891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167506501_167531501_154C;SPAN=5264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:103 GQ:4.5 PL:[0.0, 4.5, 257.4] SR:7 DR:2 LR:4.798 LO:12.35);ALT=T[chr1:167522624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167582929	-	chr9	97246437	+	.	14	0	4342036_1	32.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=4342036_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167582929(-)-9:97246437(-)__9_97240501_97265501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:52 GQ:32.3 PL:[32.3, 0.0, 91.7] SR:0 DR:14 LR:-32.13 LO:33.82);ALT=[chr9:97246437[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	167599628	+	chr1	167654655	+	.	12	0	386822_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=386822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167599628(+)-1:167654655(-)__1_167580001_167605001D;SPAN=55027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:63 GQ:22.7 PL:[22.7, 0.0, 128.3] SR:0 DR:12 LR:-22.54 LO:26.91);ALT=G[chr1:167654655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167599667	+	chr1	167653135	+	.	31	24	386823_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=386823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167580001_167605001_296C;SPAN=53468;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:74 GQ:52.7 PL:[125.3, 0.0, 52.7] SR:24 DR:31 LR:-126.7 LO:126.7);ALT=G[chr1:167653135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167653238	+	chr1	167654656	+	.	0	24	386270_1	62.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=386270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167629001_167654001_331C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:61 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:24 DR:0 LR:-62.7 LO:62.89);ALT=G[chr1:167654656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167691479	+	chr1	167734820	+	.	0	11	386579_1	21.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=386579_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167678001_167703001_52C;SPAN=43341;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:55 GQ:21.5 PL:[21.5, 0.0, 110.6] SR:11 DR:0 LR:-21.41 LO:24.93);ALT=T[chr1:167734820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167887599	+	chr1	167889217	+	.	0	19	387258_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=387258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_167874001_167899001_382C;SPAN=1618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:101 GQ:35.6 PL:[35.6, 0.0, 207.2] SR:19 DR:0 LR:-35.36 LO:42.49);ALT=T[chr1:167889217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167889920	+	chr1	167905144	+	.	8	0	387271_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=387271_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167889920(+)-1:167905144(-)__1_167874001_167899001D;SPAN=15224;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=A[chr1:167905144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	167893833	+	chr1	167905138	+	.	10	0	387285_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=387285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:167893833(+)-1:167905138(-)__1_167874001_167899001D;SPAN=11305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:0 DR:10 LR:-22.44 LO:23.91);ALT=T[chr1:167905138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168024574	+	chr1	168025733	+	.	106	53	387728_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGGCTTAAGTTTTT;MAPQ=60;MATEID=387728_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_168021001_168046001_352C;SPAN=1159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:82 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:53 DR:106 LR:-379.6 LO:379.6);ALT=T[chr1:168025733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168148419	+	chr1	168153140	+	.	19	24	388240_1	74.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=388240_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_168143501_168168501_83C;SPAN=4721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:116 GQ:74.3 PL:[74.3, 0.0, 206.3] SR:24 DR:19 LR:-74.21 LO:77.7);ALT=A[chr1:168153140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	168186185	-	chr17	74319260	+	.	9	0	388874_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=388874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:168186185(-)-17:74319260(-)__1_168168001_168193001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:63 GQ:12.8 PL:[12.8, 0.0, 138.2] SR:0 DR:9 LR:-12.64 LO:18.94);ALT=[chr17:74319260[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	168186489	+	chr3	53175885	+	TT	83	83	388883_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TT;MAPQ=60;MATEID=388883_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_168168001_168193001_141C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:62 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:83 DR:83 LR:-366.4 LO:366.4);ALT=T[chr3:53175885[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	168195382	+	chr1	168200750	+	.	9	2	388334_1	8.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=388334_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_168192501_168217501_241C;SPAN=5368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:103 GQ:8.6 PL:[8.6, 0.0, 239.6] SR:2 DR:9 LR:-8.406 LO:21.66);ALT=T[chr1:168200750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169076164	+	chr1	169080617	+	TTAAGATCA	8	9	391099_1	32.0	.	DISC_MAPQ=52;EVDNC=ASDIS;INSERTION=TTAAGATCA;MAPQ=60;MATEID=391099_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_169074501_169099501_147C;SPAN=4453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:89 GQ:32 PL:[32.0, 0.0, 183.8] SR:9 DR:8 LR:-32.01 LO:38.15);ALT=T[chr1:169080617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169094277	+	chr1	169096461	+	.	3	3	391160_1	0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=391160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_169074501_169099501_35C;SPAN=2184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:99 GQ:10.2 PL:[0.0, 10.2, 260.7] SR:3 DR:3 LR:10.32 LO:8.158);ALT=G[chr1:169096461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169292522	+	chr1	169293631	+	.	0	20	391669_1	34.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=391669_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_169270501_169295501_385C;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:117 GQ:34.4 PL:[34.4, 0.0, 248.9] SR:20 DR:0 LR:-34.32 LO:43.8);ALT=C[chr1:169293631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169292569	+	chr1	169336945	+	.	15	0	391767_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=391767_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169292569(+)-1:169336945(-)__1_169319501_169344501D;SPAN=44376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:71 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:0 DR:15 LR:-30.28 LO:34.4);ALT=A[chr1:169336945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169293754	+	chr1	169336955	+	.	14	0	391768_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=391768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169293754(+)-1:169336955(-)__1_169319501_169344501D;SPAN=43201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:0 DR:14 LR:-26.71 LO:31.54);ALT=G[chr1:169336955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169660974	+	chr1	169670655	+	.	8	0	392996_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=392996_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169660974(+)-1:169670655(-)__1_169662501_169687501D;SPAN=9681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=T[chr1:169670655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169670829	+	chr1	169672396	+	.	9	6	393026_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=393026_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_169662501_169687501_216C;SPAN=1567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:90 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:6 DR:9 LR:-11.93 LO:22.35);ALT=T[chr1:169672396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169677945	+	chr1	169679577	+	.	0	38	393051_1	92.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=393051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_169662501_169687501_184C;SPAN=1632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:120 GQ:92.9 PL:[92.9, 0.0, 198.5] SR:38 DR:0 LR:-92.93 LO:95.02);ALT=C[chr1:169679577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169677993	+	chr1	169680636	+	.	40	0	393052_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=393052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:169677993(+)-1:169680636(-)__1_169662501_169687501D;SPAN=2643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:112 GQ:99 PL:[101.9, 0.0, 167.9] SR:0 DR:40 LR:-101.7 LO:102.6);ALT=A[chr1:169680636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	169962744	+	chr11	61875134	+	AAGAGGTCTTTCAAGCATCACG	4	103	394216_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;INSERTION=AAGAGGTCTTTCAAGCATCACG;MAPQ=60;MATEID=394216_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AGAG;SCTG=c_1_169956501_169981501_190C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:19 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:103 DR:4 LR:-307.0 LO:307.0);ALT=C[chr11:61875134[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	61875192	+	chr1	169962829	+	AAG	9	70	394228_1	99.0	.	DISC_MAPQ=43;EVDNC=TSI_L;INSERTION=AAG;MAPQ=60;MATEID=394228_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CC;SCTG=c_1_169956501_169981501_190C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:46 GQ:21 PL:[231.0, 21.0, 0.0] SR:70 DR:9 LR:-231.1 LO:231.1);ALT=]chr11:61875192]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	170024579	+	chr1	170043576	+	.	6	4	394115_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=394115_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_170005501_170030501_223C;SPAN=18997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:50 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:4 DR:6 LR:-9.561 LO:14.67);ALT=T[chr1:170043576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	171454875	+	chr1	171481170	+	.	0	47	398519_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=398519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_171475501_171500501_216C;SPAN=26295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:76 GQ:48.8 PL:[134.6, 0.0, 48.8] SR:47 DR:0 LR:-136.7 LO:136.7);ALT=G[chr1:171481170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	171482311	+	chr1	171483675	+	.	0	23	398546_1	43.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=398546_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_171475501_171500501_155C;SPAN=1364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:120 GQ:43.4 PL:[43.4, 0.0, 248.0] SR:23 DR:0 LR:-43.41 LO:51.65);ALT=A[chr1:171483675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	171485032	+	chr1	171486729	+	.	12	0	398554_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=398554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:171485032(+)-1:171486729(-)__1_171475501_171500501D;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:102 GQ:12.2 PL:[12.2, 0.0, 233.3] SR:0 DR:12 LR:-11.98 LO:24.17);ALT=T[chr1:171486729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	171492661	+	chr1	171493957	+	.	6	5	398580_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=398580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_171475501_171500501_41C;SPAN=1296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:5 DR:6 LR:-7.272 LO:19.63);ALT=G[chr1:171493957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4849218	+	chr1	171639680	+	.	14	0	6294104_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6294104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:171639680(-)-17:4849218(+)__17_4826501_4851501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:14 DP:262 GQ:24.4 PL:[0.0, 24.4, 683.2] SR:0 DR:14 LR:24.77 LO:23.19);ALT=]chr17:4849218]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	171639792	+	chr17	4849923	+	.	5	28	399192_1	83.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TCTTGTCAGTCTTGGTGACAGTGACATTGAAGGTGGGGGC;MAPQ=60;MATEID=399192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_171622501_171647501_66C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:95 GQ:83.3 PL:[83.3, 0.0, 146.0] SR:28 DR:5 LR:-83.2 LO:84.17);ALT=C[chr17:4849923[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	171639989	+	chr17	4851664	+	.	20	0	6294522_1	0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6294522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:171639989(+)-17:4851664(-)__17_4851001_4876001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:20 DP:464 GQ:59.4 PL:[0.0, 59.4, 1244.0] SR:0 DR:20 LR:59.69 LO:31.23);ALT=T[chr17:4851664[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	171697222	+	chr1	171707489	+	AGAAAAAAGTCCTCTTCTTCATCTGAATCATCTTCCAAAAGATTTCT	0	11	399231_1	11.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGAAAAAAGTCCTCTTCTTCATCTGAATCATCTTCCAAAAGATTTCT;MAPQ=60;MATEID=399231_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_171696001_171721001_23C;SPAN=10267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:11 DR:0 LR:-10.84 LO:22.13);ALT=T[chr1:171707489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	171707605	+	chr1	171711048	+	.	13	11	399269_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=399269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_171696001_171721001_75C;SPAN=3443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:108 GQ:30.2 PL:[30.2, 0.0, 231.5] SR:11 DR:13 LR:-30.16 LO:39.2);ALT=T[chr1:171711048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	172411979	+	chr1	172413126	+	.	21	0	401419_1	44.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=401419_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:172411979(+)-1:172413126(-)__1_172406501_172431501D;SPAN=1147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:91 GQ:44.9 PL:[44.9, 0.0, 173.6] SR:0 DR:21 LR:-44.67 LO:49.08);ALT=A[chr1:172413126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	173446631	+	chr1	173450465	+	.	100	60	404769_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=404769_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_173435501_173460501_334C;SPAN=3834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:118 GQ:36 PL:[396.0, 36.0, 0.0] SR:60 DR:100 LR:-396.1 LO:396.1);ALT=C[chr1:173450465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	173446631	+	chr1	173454498	+	ATGGGGCATTCTCTTCTCCCACCCTCGGGACTTTACCCCAGTGTGCACCACAGAGCTTGGCAGAGCTGCAAAGCTGGCACCAGAATTTGCCAAGAGGAATGTTAAGTTGATTGCCCTTTCAATAGACAGTGTTGAGGACCATCTTGCCTGGAGCA	6	89	404770_1	99.0	.	DISC_MAPQ=51;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGGGGCATTCTCTTCTCCCACCCTCGGGACTTTACCCCAGTGTGCACCACAGAGCTTGGCAGAGCTGCAAAGCTGGCACCAGAATTTGCCAAGAGGAATGTTAAGTTGATTGCCCTTTCAATAGACAGTGTTGAGGACCATCTTGCCTGGAGCA;MAPQ=60;MATEID=404770_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_173435501_173460501_334C;SPAN=7867;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:100 GQ:27 PL:[297.0, 27.0, 0.0] SR:89 DR:6 LR:-297.1 LO:297.1);ALT=C[chr1:173454498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	173450622	+	chr1	173454498	+	.	2	25	404786_1	53.0	.	DISC_MAPQ=49;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=404786_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_1_173435501_173460501_334C;SPAN=3876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:132 GQ:53.6 PL:[53.6, 0.0, 264.8] SR:25 DR:2 LR:-53.37 LO:61.49);ALT=G[chr1:173454498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	173455541	+	chr1	173456872	+	.	9	24	404798_1	69.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=57;MATEID=404798_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_173435501_173460501_40C;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:120 GQ:69.8 PL:[69.8, 0.0, 221.6] SR:24 DR:9 LR:-69.82 LO:74.22);ALT=G[chr1:173456872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	174128798	+	chr1	174188261	+	.	7	5	407682_1	19.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=407682_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_174170501_174195501_215C;SPAN=59463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:5 DR:7 LR:-19.73 LO:22.76);ALT=G[chr1:174188261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	89181129	+	chr1	174471740	+	.	16	25	3444653_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=ATATATGTGTGTATATA;MAPQ=60;MATEID=3444653_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_7_89180001_89205001_14C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:47 GQ:10.4 PL:[102.8, 0.0, 10.4] SR:25 DR:16 LR:-107.1 LO:107.1);ALT=]chr7:89181129]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	174471803	+	chr7	89181110	+	.	22	35	3444656_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=CATATATATGTGTGT;MAPQ=55;MATEID=3444656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_89180001_89205001_375C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:46 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:35 DR:22 LR:-135.3 LO:135.3);ALT=T[chr7:89181110[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	174969320	+	chr2	184472885	-	.	18	0	1120394_1	43.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1120394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:174969320(+)-2:184472885(+)__2_184460501_184485501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:59 GQ:43.4 PL:[43.4, 0.0, 99.5] SR:0 DR:18 LR:-43.43 LO:44.65);ALT=G]chr2:184472885];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	174969358	+	chr1	174973747	+	.	52	0	410248_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=410248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:174969358(+)-1:174973747(-)__1_174954501_174979501D;SPAN=4389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:110 GQ:99 PL:[141.8, 0.0, 125.3] SR:0 DR:52 LR:-141.9 LO:141.9);ALT=A[chr1:174973747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	174983989	+	chr1	174987553	+	.	0	15	410293_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=410293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_174979001_175004001_282C;SPAN=3564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:120 GQ:17 PL:[17.0, 0.0, 274.4] SR:15 DR:0 LR:-17.0 LO:30.63);ALT=T[chr1:174987553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	174984037	+	chr1	174992499	+	.	11	0	410294_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=410294_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:174984037(+)-1:174992499(-)__1_174979001_175004001D;SPAN=8462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:129 GQ:1.4 PL:[1.4, 0.0, 311.6] SR:0 DR:11 LR:-1.362 LO:20.53);ALT=T[chr1:174992499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	174987726	+	chr1	174992490	+	.	16	0	410313_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=410313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:174987726(+)-1:174992490(-)__1_174979001_175004001D;SPAN=4764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:140 GQ:14.9 PL:[14.9, 0.0, 325.1] SR:0 DR:16 LR:-14.89 LO:32.01);ALT=A[chr1:174992490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	175200569	+	chr1	175201937	-	.	50	55	411167_1	99.0	.	DISC_MAPQ=28;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=411167_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_175199501_175224501_362C;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:64 GQ:24 PL:[264.0, 24.0, 0.0] SR:55 DR:50 LR:-264.1 LO:264.1);ALT=A]chr1:175201937];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	155949600	+	chr1	175401048	+	.	4	18	411746_1	52.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TCTCTCTCTCTCTCTCTCTCTCTC;MAPQ=60;MATEID=411746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_175395501_175420501_332C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:18 DR:4 LR:-52.2 LO:52.37);ALT=]chr2:155949600]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	182274475	+	chr17	74319261	+	AAAAAAAAAAAA	38	25	435733_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=AAAAAAAAAAAA;MAPQ=60;MATEID=435733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_182255501_182280501_315C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:52 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:25 DR:38 LR:-155.1 LO:155.1);ALT=A[chr17:74319261[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	182342851	-	chr1	182344042	+	.	14	0	435218_1	21.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=435218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:182342851(-)-1:182344042(-)__1_182329001_182354001D;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:0 DR:14 LR:-21.29 LO:29.89);ALT=[chr1:182344042[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	182356429	+	chr1	182357707	+	.	2	25	435482_1	55.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=435482_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_182353501_182378501_97C;SPAN=1278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:126 GQ:55.1 PL:[55.1, 0.0, 249.8] SR:25 DR:2 LR:-54.99 LO:62.11);ALT=T[chr1:182357707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	182356456	+	chr1	182360864	+	.	9	0	435483_1	0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=435483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:182356456(+)-1:182360864(-)__1_182353501_182378501D;SPAN=4408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:143 GQ:8.7 PL:[0.0, 8.7, 363.0] SR:0 DR:9 LR:9.033 LO:15.57);ALT=T[chr1:182360864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	182357889	+	chr1	182360814	+	.	84	13	435488_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=435488_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_182353501_182378501_373C;SPAN=2925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:122 GQ:23.3 PL:[270.8, 0.0, 23.3] SR:13 DR:84 LR:-282.5 LO:282.5);ALT=G[chr1:182360814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	182808576	+	chr1	182811697	+	.	10	0	437220_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=437220_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:182808576(+)-1:182811697(-)__1_182794501_182819501D;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=C[chr1:182811697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183556114	+	chr1	183559290	+	.	0	11	439713_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=439713_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_183554001_183579001_366C;SPAN=3176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:111 GQ:6.5 PL:[6.5, 0.0, 260.6] SR:11 DR:0 LR:-6.238 LO:21.28);ALT=T[chr1:183559290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183596731	+	chr1	183599595	+	.	5	15	439932_1	32.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=439932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_183578501_183603501_273C;SPAN=2864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:123 GQ:32.9 PL:[32.9, 0.0, 263.9] SR:15 DR:5 LR:-32.7 LO:43.32);ALT=T[chr1:183599595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183599774	+	chr1	183602216	+	.	3	51	439942_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=439942_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_183578501_183603501_113C;SPAN=2442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:134 GQ:99 PL:[142.1, 0.0, 181.7] SR:51 DR:3 LR:-142.0 LO:142.2);ALT=T[chr1:183602216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183599774	+	chr1	183604651	+	TCACTGCCTGACTCTTGGTGTTGATAGGGGGGTTCTTCAGAGCTGCCTGTAGGGCAGCTGTCATGTTTCC	24	79	439943_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=T;INSERTION=TCACTGCCTGACTCTTGGTGTTGATAGGGGGGTTCTTCAGAGCTGCCTGTAGGGCAGCTGTCATGTTTCC;MAPQ=60;MATEID=439943_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_183578501_183603501_113C;SPAN=4877;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:74 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:79 DR:24 LR:-260.8 LO:260.8);ALT=T[chr1:183604651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	183602343	+	chr1	183604752	+	.	62	0	439783_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=439783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:183602343(+)-1:183604752(-)__1_183603001_183628001D;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:89 GQ:35.3 PL:[180.5, 0.0, 35.3] SR:0 DR:62 LR:-186.1 LO:186.1);ALT=A[chr1:183604752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	184020950	+	chr1	184023485	+	.	8	0	441048_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=441048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:184020950(+)-1:184023485(-)__1_184019501_184044501D;SPAN=2535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:0 DR:8 LR:0.4135 LO:14.74);ALT=G[chr1:184023485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	184020961	+	chr1	184023861	+	.	12	0	441049_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=441049_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:184020961(+)-1:184023861(-)__1_184019501_184044501D;SPAN=2900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:114 GQ:8.9 PL:[8.9, 0.0, 266.3] SR:0 DR:12 LR:-8.727 LO:23.55);ALT=T[chr1:184023861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	184868475	+	chr1	184943525	+	.	8	0	443866_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=443866_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:184868475(+)-1:184943525(-)__1_184852501_184877501D;SPAN=75050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=A[chr1:184943525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	185014781	+	chr1	185056683	+	.	5	7	444079_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=444079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_184999501_185024501_350C;SPAN=41902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:7 DR:5 LR:-16.65 LO:18.55);ALT=G[chr1:185056683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	103156483	+	chr1	188827982	+	.	8	0	2120874_1	9.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=2120874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:188827982(-)-4:103156483(+)__4_103145001_103170001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:0 DR:8 LR:-9.34 LO:16.4);ALT=]chr4:103156483]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	201115977	+	chr1	201120889	+	.	0	10	492189_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=492189_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_201096001_201121001_372C;SPAN=4912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:126 GQ:0.9 PL:[0.0, 0.9, 306.9] SR:10 DR:0 LR:1.127 LO:18.34);ALT=C[chr1:201120889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201181092	+	chr1	201179775	+	.	31	0	492236_1	69.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=492236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201179775(-)-1:201181092(+)__1_201169501_201194501D;SPAN=1317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:122 GQ:69.5 PL:[69.5, 0.0, 224.6] SR:0 DR:31 LR:-69.28 LO:73.96);ALT=]chr1:201181092]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	201458112	+	chr1	201459304	+	.	0	14	493159_1	16.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=493159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_201439001_201464001_309C;SPAN=1192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:109 GQ:16.7 PL:[16.7, 0.0, 247.7] SR:14 DR:0 LR:-16.68 LO:28.77);ALT=T[chr1:201459304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201459472	+	chr1	201465320	+	.	0	24	493182_1	65.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=493182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_201463501_201488501_397C;SPAN=5848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:51 GQ:55.7 PL:[65.6, 0.0, 55.7] SR:24 DR:0 LR:-65.43 LO:65.43);ALT=A[chr1:201465320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201459515	+	chr1	201476196	+	.	33	0	493183_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=493183_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201459515(+)-1:201476196(-)__1_201463501_201488501D;SPAN=16681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:43 GQ:5 PL:[97.4, 0.0, 5.0] SR:0 DR:33 LR:-101.9 LO:101.9);ALT=G[chr1:201476196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201465461	+	chr1	201476197	+	.	11	0	493193_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=493193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201465461(+)-1:201476197(-)__1_201463501_201488501D;SPAN=10736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:109 GQ:6.8 PL:[6.8, 0.0, 257.6] SR:0 DR:11 LR:-6.78 LO:21.38);ALT=A[chr1:201476197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201612566	+	chr1	201611191	+	.	15	0	493651_1	32.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=493651_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201611191(-)-1:201612566(+)__1_201610501_201635501D;SPAN=1375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:0 DR:15 LR:-32.72 LO:35.42);ALT=]chr1:201612566]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	201924726	+	chr1	201932741	+	.	17	0	495027_1	40.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=495027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201924726(+)-1:201932741(-)__1_201929001_201954001D;SPAN=8015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:59 GQ:40.1 PL:[40.1, 0.0, 102.8] SR:0 DR:17 LR:-40.13 LO:41.66);ALT=C[chr1:201932741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201924726	+	chr1	201926636	+	.	21	0	494765_1	31.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=494765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:201924726(+)-1:201926636(-)__1_201904501_201929501D;SPAN=1910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:142 GQ:31.1 PL:[31.1, 0.0, 311.6] SR:0 DR:21 LR:-30.85 LO:44.54);ALT=C[chr1:201926636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	201926705	+	chr1	201932742	+	.	3	31	495029_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=495029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_201929001_201954001_126C;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:60 GQ:49.7 PL:[95.9, 0.0, 49.7] SR:31 DR:3 LR:-96.77 LO:96.77);ALT=A[chr1:201932742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202127476	+	chr1	202129669	+	.	20	0	495546_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=495546_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:202127476(+)-1:202129669(-)__1_202125001_202150001D;SPAN=2193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:125 GQ:32.3 PL:[32.3, 0.0, 269.9] SR:0 DR:20 LR:-32.15 LO:43.17);ALT=G[chr1:202129669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202301090	+	chr1	202302137	+	.	2	5	496649_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=496649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_202296501_202321501_316C;SPAN=1047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:5 DR:2 LR:1.547 LO:12.74);ALT=T[chr1:202302137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202304908	+	chr1	202311021	+	.	8	0	496662_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=496662_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:202304908(+)-1:202311021(-)__1_202296501_202321501D;SPAN=6113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:128 GQ:8.1 PL:[0.0, 8.1, 326.7] SR:0 DR:8 LR:8.27 LO:13.81);ALT=A[chr1:202311021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202828254	+	chr1	202830592	+	.	8	0	498505_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=498505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:202828254(+)-1:202830592(-)__1_202811001_202836001D;SPAN=2338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=T[chr1:202830592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	202828524	-	chr1	202829565	+	.	8	0	498506_1	1.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=498506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:202828524(-)-1:202829565(-)__1_202811001_202836001D;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:0 DR:8 LR:-0.9411 LO:14.92);ALT=[chr1:202829565[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	202844794	+	chr6	90582117	-	.	8	13	2938285_1	60.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=GGTGAAACCCCGTCTCTACTAAAAATACAAAAAATTAGCCGGGCACAGTGGC;MAPQ=60;MATEID=2938285_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_90576501_90601501_116C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:32 GQ:14.6 PL:[60.8, 0.0, 14.6] SR:13 DR:8 LR:-62.01 LO:62.01);ALT=C]chr6:90582117];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	202920292	+	chr1	202927313	+	.	56	8	498953_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=498953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_202909001_202934001_304C;SPAN=7021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:109 GQ:99 PL:[165.2, 0.0, 99.2] SR:8 DR:56 LR:-166.1 LO:166.1);ALT=A[chr1:202927313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	203274876	+	chr1	203276227	+	.	0	23	500108_1	46.0	.	EVDNC=ASSMB;HOMSEQ=CACAG;MAPQ=60;MATEID=500108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_203252001_203277001_11C;SPAN=1351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:110 GQ:46.1 PL:[46.1, 0.0, 221.0] SR:23 DR:0 LR:-46.12 LO:52.63);ALT=G[chr1:203276227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	203830843	+	chr19	5576940	-	.	86	0	6708348_1	99.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=6708348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:203830843(+)-19:5576940(+)__19_5561501_5586501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:47 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:0 DR:86 LR:-254.2 LO:254.2);ALT=T]chr19:5576940];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	203830843	+	chr9	6748969	-	.	35	0	4132425_1	99.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4132425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:203830843(+)-9:6748969(+)__9_6737501_6762501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:27 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:35 LR:-102.3 LO:102.3);ALT=T]chr9:6748969];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	204485667	+	chr1	204494608	+	.	13	0	505061_1	13.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=505061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:204485667(+)-1:204494608(-)__1_204477001_204502001D;SPAN=8941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:111 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:0 DR:13 LR:-12.84 LO:26.15);ALT=G[chr1:204494608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	204485739	+	chr1	204495482	+	.	12	0	505063_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=505063_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:204485739(+)-1:204495482(-)__1_204477001_204502001D;SPAN=9743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:111 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:0 DR:12 LR:-9.539 LO:23.7);ALT=G[chr1:204495482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	204516006	+	chr1	204518239	+	.	0	7	505216_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=505216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_204501501_204526501_199C;SPAN=2233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:88 GQ:0.6 PL:[0.0, 0.6, 214.5] SR:7 DR:0 LR:0.7344 LO:12.84);ALT=G[chr1:204518239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220156742	+	chr1	220160482	+	GAGAATACCAATCAGCAAGATTTTCTTCTTTTTTTGCCTCAAGACCCA	0	9	556135_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=GAGAATACCAATCAGCAAGATTTTCTTCTTTTTTTGCCTCAAGACCCA;MAPQ=60;MATEID=556135_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_220157001_220182001_261C;SPAN=3740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:9 DR:0 LR:-16.43 LO:20.02);ALT=T[chr1:220160482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220193563	+	chr1	220195689	+	.	4	4	556492_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=556492_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_220181501_220206501_58C;SPAN=2126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:101 GQ:3.9 PL:[0.0, 3.9, 250.8] SR:4 DR:4 LR:4.256 LO:12.41);ALT=A[chr1:220195689[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220203823	+	chr1	220205728	+	.	0	9	556531_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=556531_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_220181501_220206501_10C;SPAN=1905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:113 GQ:0.6 PL:[0.0, 0.6, 273.9] SR:9 DR:0 LR:0.9055 LO:16.52);ALT=C[chr1:220205728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220207002	+	chr1	220208256	+	.	0	6	557172_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=557172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_220206001_220231001_165C;SPAN=1254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:100 GQ:7.2 PL:[0.0, 7.2, 257.4] SR:6 DR:0 LR:7.287 LO:10.25);ALT=T[chr1:220208256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220208410	+	chr1	220219724	+	.	8	0	557180_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=557180_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:220208410(+)-1:220219724(-)__1_220206001_220231001D;SPAN=11314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=C[chr1:220219724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220213785	+	chr1	220219735	+	.	11	0	557221_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=557221_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:220213785(+)-1:220219735(-)__1_220206001_220231001D;SPAN=5950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:104 GQ:8.3 PL:[8.3, 0.0, 242.6] SR:0 DR:11 LR:-8.135 LO:21.61);ALT=A[chr1:220219735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	220273991	+	chr1	220275469	+	.	0	6	556845_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=556845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_220255001_220280001_112C;SPAN=1478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:83 GQ:2.4 PL:[0.0, 2.4, 204.6] SR:6 DR:0 LR:2.681 LO:10.75);ALT=G[chr1:220275469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	79165470	+	chr1	220426919	+	.	8	0	557622_1	0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=557622_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:220426919(-)-15:79165470(+)__1_220402001_220427001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:113 GQ:3.9 PL:[0.0, 3.9, 280.5] SR:0 DR:8 LR:4.207 LO:14.26);ALT=]chr15:79165470]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	221356192	+	chr11	22215160	+	.	10	0	4788723_1	20.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=4788723_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:221356192(+)-11:22215160(-)__11_22197001_22222001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:0 DR:10 LR:-20.82 LO:23.18);ALT=G[chr11:22215160[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	221913157	+	chr1	221915340	+	.	32	0	561828_1	78.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=561828_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:221913157(+)-1:221915340(-)__1_221896501_221921501D;SPAN=2183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:101 GQ:78.5 PL:[78.5, 0.0, 164.3] SR:0 DR:32 LR:-78.27 LO:80.03);ALT=A[chr1:221915340[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	222886284	+	chr1	222889025	+	.	4	2	565153_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=565153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_222876501_222901501_28C;SPAN=2741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:104 GQ:14.7 PL:[0.0, 14.7, 280.5] SR:2 DR:4 LR:14.97 LO:6.046);ALT=G[chr1:222889025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	224302100	+	chr1	224318173	+	.	2	9	570131_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=570131_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_224297501_224322501_232C;SPAN=16073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:129 GQ:1.4 PL:[1.4, 0.0, 311.6] SR:9 DR:2 LR:-1.362 LO:20.53);ALT=T[chr1:224318173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	224544693	+	chr1	224553578	+	.	11	0	571578_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=571578_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:224544693(+)-1:224553578(-)__1_224542501_224567501D;SPAN=8885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:113 GQ:5.9 PL:[5.9, 0.0, 266.6] SR:0 DR:11 LR:-5.697 LO:21.19);ALT=T[chr1:224553578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	224553693	+	chr1	224558984	+	.	3	4	571623_1	0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=571623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_224542501_224567501_197C;SPAN=5291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:108 GQ:6 PL:[0.0, 6.0, 273.9] SR:4 DR:3 LR:6.153 LO:12.2);ALT=G[chr1:224558984[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	224559125	+	chr1	224563495	+	.	0	8	571653_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=571653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_224542501_224567501_103C;SPAN=4370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:8 DR:0 LR:0.4135 LO:14.74);ALT=G[chr1:224563495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	224800120	+	chr1	224646603	+	CAAAACTTACTATAGCAGTTCTGTGAGCTGCTCTAGC	0	66	572074_1	99.0	.	EVDNC=ASSMB;INSERTION=CAAAACTTACTATAGCAGTTCTGTGAGCTGCTCTAGC;MAPQ=60;MATEID=572074_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_224640501_224665501_202C;SPAN=153517;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:63 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:66 DR:0 LR:-194.7 LO:194.7);ALT=]chr1:224800120]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr1	224782795	+	chr1	224786034	+	CTATAGTAGAACTTCTTTT	0	48	572731_1	99.0	.	EVDNC=ASSMB;INSERTION=CTATAGTAGAACTTCTTTT;MAPQ=60;MATEID=572731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_224763001_224788001_188C;SPAN=3239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:123 GQ:99 PL:[125.3, 0.0, 171.5] SR:48 DR:0 LR:-125.1 LO:125.6);ALT=C[chr1:224786034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	225133672	+	chr1	225248642	+	.	49	0	574239_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=574239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:225133672(+)-1:225248642(-)__1_225228501_225253501D;SPAN=114970;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:20 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:49 LR:-145.2 LO:145.2);ALT=C[chr1:225248642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	225235952	-	chr1	225236953	+	.	9	0	574257_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=574257_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:225235952(-)-1:225236953(-)__1_225228501_225253501D;SPAN=1001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:117 GQ:1.8 PL:[0.0, 1.8, 287.1] SR:0 DR:9 LR:1.989 LO:16.38);ALT=[chr1:225236953[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	225272506	+	chr15	27461950	-	.	8	44	574495_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=574495_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_225253001_225278001_96C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:19 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:44 DR:8 LR:-138.6 LO:138.6);ALT=C]chr15:27461950];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	225611815	+	chr1	225615668	+	.	18	0	575298_1	35.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=575298_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:225611815(+)-1:225615668(-)__1_225596001_225621001D;SPAN=3853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:0 DR:18 LR:-35.58 LO:40.99);ALT=T[chr1:225615668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	226110084	+	chr1	226111741	+	CTGAGCGCGGACACCGTGGGCAGGTTCATTTCTGGGGAGCTGGCTATTATCTTGTGAGCCGACAGGA	14	39	577198_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TGCCTGC;INSERTION=CTGAGCGCGGACACCGTGGGCAGGTTCATTTCTGGGGAGCTGGCTATTATCTTGTGAGCCGACAGGA;MAPQ=60;MATEID=577198_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_226110501_226135501_83C;SPAN=1657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:59 GQ:13.7 PL:[129.2, 0.0, 13.7] SR:39 DR:14 LR:-134.7 LO:134.7);ALT=C[chr1:226111741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79213215	+	chr1	226314956	+	.	14	0	6516536_1	32.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6516536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:226314956(-)-17:79213215(+)__17_79208501_79233501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:52 GQ:32.3 PL:[32.3, 0.0, 91.7] SR:0 DR:14 LR:-32.13 LO:33.82);ALT=]chr17:79213215]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	226578327	+	chr1	226579899	+	.	0	16	579255_1	22.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=579255_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_226576001_226601001_251C;SPAN=1572;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:114 GQ:22.1 PL:[22.1, 0.0, 253.1] SR:16 DR:0 LR:-21.93 LO:33.54);ALT=T[chr1:226579899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	226590082	+	chr1	226595511	+	.	0	23	579300_1	47.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=579300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_226576001_226601001_82C;SPAN=5429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:105 GQ:47.6 PL:[47.6, 0.0, 206.0] SR:23 DR:0 LR:-47.48 LO:53.16);ALT=T[chr1:226595511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	227128097	+	chr1	227149073	+	.	8	0	581748_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=581748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:227128097(+)-1:227149073(-)__1_227115001_227140001D;SPAN=20976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:0 DR:8 LR:-10.97 LO:16.77);ALT=C[chr1:227149073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228270547	+	chr1	228284776	+	.	140	0	585393_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=585393_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228270547(+)-1:228284776(-)__1_228266501_228291501D;SPAN=14229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:78 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:0 DR:140 LR:-415.9 LO:415.9);ALT=T[chr1:228284776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228295620	+	chr1	228296902	+	.	35	0	585862_1	93.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=585862_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228295620(+)-1:228296902(-)__1_228291001_228316001D;SPAN=1282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:80 GQ:93.8 PL:[93.8, 0.0, 100.4] SR:0 DR:35 LR:-93.86 LO:93.87);ALT=T[chr1:228296902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228302857	+	chr15	64380885	+	TCGCTGAAGTTTTACTCTTAAGCACAGC	0	7	5970659_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TCGCTGAAGTTTTACTCTTAAGCACAGC;MAPQ=54;MATEID=5970659_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_64361501_64386501_66C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:25 GQ:16.4 PL:[16.4, 0.0, 42.8] SR:7 DR:0 LR:-16.33 LO:17.05);ALT=A[chr15:64380885[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	228303103	+	chr15	64385933	+	.	9	0	5970663_1	16.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=5970663_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228303103(+)-15:64385933(-)__15_64361501_64386501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=C[chr15:64385933[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	228328065	+	chr1	228333211	+	.	50	15	585707_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=585707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_228315501_228340501_25C;SPAN=5146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:148 GQ:99 PL:[144.8, 0.0, 214.1] SR:15 DR:50 LR:-144.8 LO:145.5);ALT=G[chr1:228333211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228328100	+	chr1	228334539	+	.	56	0	585709_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=585709_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228328100(+)-1:228334539(-)__1_228315501_228340501D;SPAN=6439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:118 GQ:99 PL:[152.9, 0.0, 133.1] SR:0 DR:56 LR:-153.0 LO:153.0);ALT=G[chr1:228334539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228328109	+	chr1	228333726	+	.	17	0	585710_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=585710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:228328109(+)-1:228333726(-)__1_228315501_228340501D;SPAN=5617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:126 GQ:22.1 PL:[22.1, 0.0, 282.8] SR:0 DR:17 LR:-21.98 LO:35.32);ALT=G[chr1:228333726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228328990	+	chr1	228333210	+	.	0	10	585714_1	6.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=585714_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_228315501_228340501_332C;SPAN=4220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:10 DR:0 LR:-6.73 LO:19.53);ALT=G[chr1:228333210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	228333325	+	chr1	228334541	+	ATACCACGAGGAACCCGAGGCCCGGCGAGGAGAACGGCAA	3	130	585721_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATACCACGAGGAACCCGAGGCCCGGCGAGGAGAACGGCAA;MAPQ=60;MATEID=585721_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_228315501_228340501_241C;SPAN=1216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:130 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:130 DR:3 LR:-389.5 LO:389.5);ALT=C[chr1:228334541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	229407117	+	chr1	229424476	+	ATTTTTTGTTTAAGTTCTTGGTTATTGGAAATGCAGGAACTGGCAAATCTTGCTTACTTCATCAGTTTATTGAAAAAAAAT	0	40	589760_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATTTTTTGTTTAAGTTCTTGGTTATTGGAAATGCAGGAACTGGCAAATCTTGCTTACTTCATCAGTTTATTGAAAAAAAAT;MAPQ=60;MATEID=589760_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_229393501_229418501_136C;SPAN=17359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:40 DR:0 LR:-118.8 LO:118.8);ALT=G[chr1:229424476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	229407117	+	chr1	229422232	+	.	20	22	589646_1	85.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=589646_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTTTT;SCTG=c_1_229418001_229443001_378C;SPAN=15115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:22 DR:20 LR:-86.31 LO:86.31);ALT=G[chr1:229422232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	229434821	+	chr1	229438607	+	.	2	4	589690_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=589690_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_229418001_229443001_199C;SPAN=3786;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:96 GQ:9.3 PL:[0.0, 9.3, 250.8] SR:4 DR:2 LR:9.504 LO:8.227);ALT=T[chr1:229438607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	229812537	+	chr1	229820837	+	.	100	80	591106_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTGT;MAPQ=60;MATEID=591106_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_1_229810001_229835001_227C;SPAN=8300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:38 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:80 DR:100 LR:-435.7 LO:435.7);ALT=T[chr1:229820837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	230203153	+	chr1	230227334	+	.	16	5	594030_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=594030_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_1_230226501_230251501_282C;SPAN=24181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:57 GQ:40.7 PL:[40.7, 0.0, 96.8] SR:5 DR:16 LR:-40.67 LO:41.97);ALT=G[chr1:230227334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	230210996	+	chr12	51892570	-	.	4	42	5189841_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GGAGGCTGAGGCA;MAPQ=35;MATEID=5189841_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_12_51891001_51916001_132C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:46 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:42 DR:4 LR:-135.3 LO:135.3);ALT=C]chr12:51892570];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr1	230385017	+	chr1	230386203	+	.	0	5	594564_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=594564_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_230373501_230398501_257C;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:114 GQ:14.1 PL:[0.0, 14.1, 303.6] SR:5 DR:0 LR:14.38 LO:7.847);ALT=A[chr1:230386203[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	231374946	+	chr1	231376839	+	.	10	0	597974_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=597974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:231374946(+)-1:231376839(-)__1_231353501_231378501D;SPAN=1893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:108 GQ:3.8 PL:[3.8, 0.0, 257.9] SR:0 DR:10 LR:-3.75 LO:19.04);ALT=A[chr1:231376839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	231377202	+	chr1	231396252	+	.	2	2	597986_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=597986_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_231378001_231403001_186C;SPAN=19050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:46 GQ:0.8 PL:[0.8, 0.0, 109.7] SR:2 DR:2 LR:-0.7415 LO:7.501);ALT=G[chr1:231396252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	231377202	+	chr1	231386706	+	.	9	16	597985_1	46.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=597985_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_231378001_231403001_329C;SPAN=9504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:62 GQ:46.1 PL:[46.1, 0.0, 102.2] SR:16 DR:9 LR:-45.92 LO:47.18);ALT=G[chr1:231386706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	231658385	+	chr1	231664165	+	TCGTGCCAGAGCAGAACATGCCTTGTAGTTACTGCCATATTCTAGCCAAGTTACTCCATTTACTGTTCCTTTGTT	0	8	598948_1	2.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCGTGCCAGAGCAGAACATGCCTTGTAGTTACTGCCATATTCTAGCCAAGTTACTCCATTTACTGTTCCTTTGTT;MAPQ=60;MATEID=598948_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_231647501_231672501_139C;SPAN=5780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-2.025 LO:15.08);ALT=T[chr1:231664165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	231663161	+	chr1	231664165	+	.	2	4	598965_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=598965_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTTT;SCTG=c_1_231647501_231672501_139C;SPAN=1004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:94 GQ:10.2 PL:[0.0, 10.2, 221.9] SR:4 DR:2 LR:10.47 LO:6.784);ALT=C[chr1:231664165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235095664	+	chr1	235104135	+	.	3	23	610878_1	70.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=610878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_235102001_235127001_435C;SPAN=8471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:44 GQ:34.4 PL:[70.7, 0.0, 34.4] SR:23 DR:3 LR:-71.2 LO:71.2);ALT=C[chr1:235104135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235095711	+	chr1	235116436	+	.	9	0	610879_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=610879_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235095711(+)-1:235116436(-)__1_235102001_235127001D;SPAN=20725;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:0 DR:9 LR:-14.27 LO:19.37);ALT=A[chr1:235116436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235104238	+	chr1	235116403	+	.	13	5	610897_1	25.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=C;MAPQ=55;MATEID=610897_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_235102001_235127001_243C;SPAN=12165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:103 GQ:25.1 PL:[25.1, 0.0, 223.1] SR:5 DR:13 LR:-24.91 LO:34.31);ALT=C[chr1:235116403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235109071	+	chr1	235116402	+	.	9	1	610909_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=610909_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_235102001_235127001_346C;SPAN=7331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:1 DR:9 LR:-2.075 LO:16.94);ALT=C[chr1:235116402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66019165	+	chr1	235291963	+	.	22	0	611478_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=611478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235291963(-)-7:66019165(+)__1_235273501_235298501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:128 GQ:38 PL:[38.0, 0.0, 272.3] SR:0 DR:22 LR:-37.94 LO:48.24);ALT=]chr7:66019165]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	235291967	-	chrX	72443018	+	.	34	0	611479_1	77.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=611479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235291967(-)-23:72443018(-)__1_235273501_235298501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:130 GQ:77 PL:[77.0, 0.0, 238.7] SR:0 DR:34 LR:-77.01 LO:81.62);ALT=[chrX:72443018[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	235318429	+	chr1	235323825	+	.	3	4	611721_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=611721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_235322501_235347501_415C;SPAN=5396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:42 GQ:8.6 PL:[8.6, 0.0, 91.1] SR:4 DR:3 LR:-8.427 LO:12.63);ALT=T[chr1:235323825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235392702	+	chr1	235394428	+	.	2	5	611593_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=611593_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_1_235371501_235396501_37C;SPAN=1726;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:97 GQ:6.3 PL:[0.0, 6.3, 247.5] SR:5 DR:2 LR:6.474 LO:10.33);ALT=T[chr1:235394428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235491973	+	chr1	235498556	+	.	9	0	612154_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=612154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235491973(+)-1:235498556(-)__1_235494001_235519001D;SPAN=6583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=T[chr1:235498556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235992343	+	chr1	235993526	+	.	0	24	614258_1	45.0	.	EVDNC=ASSMB;HOMSEQ=CTGA;MAPQ=60;MATEID=614258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_235984001_236009001_139C;SPAN=1183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:124 GQ:45.8 PL:[45.8, 0.0, 253.7] SR:24 DR:0 LR:-45.63 LO:54.01);ALT=A[chr1:235993526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235993725	+	chr1	235996878	+	.	2	27	614262_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=614262_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_235984001_236009001_248C;SPAN=3153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:124 GQ:62.3 PL:[62.3, 0.0, 237.2] SR:27 DR:2 LR:-62.13 LO:67.97);ALT=C[chr1:235996878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235993764	+	chr1	236030139	+	.	58	0	614263_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=614263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235993764(+)-1:236030139(-)__1_235984001_236009001D;SPAN=36375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:45 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=C[chr1:236030139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	235996977	+	chr1	236030140	+	.	14	0	614274_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=614274_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:235996977(+)-1:236030140(-)__1_235984001_236009001D;SPAN=33163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:47 GQ:33.5 PL:[33.5, 0.0, 79.7] SR:0 DR:14 LR:-33.48 LO:34.55);ALT=A[chr1:236030140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	236549103	+	chr1	236551330	+	.	69	56	616486_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TAATAATTTGAAAGTTA;MAPQ=60;MATEID=616486_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_236547501_236572501_394C;SPAN=2227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:37 GQ:27 PL:[297.0, 27.0, 0.0] SR:56 DR:69 LR:-297.1 LO:297.1);ALT=A[chr1:236551330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	236687389	+	chr1	236689266	+	.	10	0	616952_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=616952_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:236687389(+)-1:236689266(-)__1_236670001_236695001D;SPAN=1877;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:117 GQ:1.4 PL:[1.4, 0.0, 281.9] SR:0 DR:10 LR:-1.312 LO:18.67);ALT=T[chr1:236689266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	244601072	+	chr1	244614936	+	.	0	16	643315_1	39.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=55;MATEID=643315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_244583501_244608501_295C;SPAN=13864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:16 DR:0 LR:-39.54 LO:40.27);ALT=T[chr1:244614936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	244999086	+	chr1	245006341	+	.	13	0	644962_1	24.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=644962_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:244999086(+)-1:245006341(-)__1_244975501_245000501D;SPAN=7255;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:68 GQ:24.5 PL:[24.5, 0.0, 140.0] SR:0 DR:13 LR:-24.49 LO:29.18);ALT=C[chr1:245006341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	244999096	+	chr2	231822463	+	.	9	0	1236167_1	16.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=1236167_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:244999096(+)-2:231822463(-)__2_231819001_231844001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=G[chr2:231822463[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr1	245018823	-	chr14	43769615	+	.	13	0	644838_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=644838_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:245018823(-)-14:43769615(-)__1_245000001_245025001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:0 DR:13 LR:-20.7 LO:28.0);ALT=[chr14:43769615[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	245023776	+	chr1	245025763	+	.	8	10	644974_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=644974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_245024501_245049501_1C;SPAN=1987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:46 GQ:33.8 PL:[33.8, 0.0, 76.7] SR:10 DR:8 LR:-33.75 LO:34.71);ALT=T[chr1:245025763[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	245912967	+	chr1	245927342	+	.	7	22	648360_1	64.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=648360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_245906501_245931501_109C;SPAN=14375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:115 GQ:64.7 PL:[64.7, 0.0, 213.2] SR:22 DR:7 LR:-64.57 LO:69.08);ALT=C[chr1:245927342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	245927454	+	chr1	246021797	+	.	2	6	648527_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=648527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246004501_246029501_232C;SPAN=94343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:6 DR:2 LR:-11.24 LO:16.84);ALT=G[chr1:246021797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246078944	+	chr1	246093172	+	CCTCTCCCACCTCGATGTCTCGGACTGCTCGCAGTAAGAGGTGGGGCCCATTGAACACAATCGAACAGTTGGGGTCACAGCTGTGATTGAGCAAAGAGATA	0	86	648781_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTGG;INSERTION=CCTCTCCCACCTCGATGTCTCGGACTGCTCGCAGTAAGAGGTGGGGCCCATTGAACACAATCGAACAGTTGGGGTCACAGCTGTGATTGAGCAAAGAGATA;MAPQ=60;MATEID=648781_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_246078001_246103001_398C;SPAN=14228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:129 GQ:64.1 PL:[248.9, 0.0, 64.1] SR:86 DR:0 LR:-255.0 LO:255.0);ALT=T[chr1:246093172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246078944	+	chr1	246091233	+	.	0	23	649822_1	66.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=649822_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_1_246347501_246372501_96C;SPAN=12289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:0 GQ:6 PL:[66.0, 6.0, 0.0] SR:23 DR:0 LR:-66.02 LO:66.02);ALT=T[chr1:246091233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246091389	+	chr1	246350042	+	.	37	0	649825_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=649825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:246091389(+)-1:246350042(-)__1_246347501_246372501D;SPAN=258653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:76 GQ:81.8 PL:[101.6, 0.0, 81.8] SR:0 DR:37 LR:-101.6 LO:101.6);ALT=A[chr1:246350042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246093239	+	chr1	246350043	+	.	0	38	649826_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=649826_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246347501_246372501_26C;SPAN=256804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:77 GQ:81.5 PL:[104.6, 0.0, 81.5] SR:38 DR:0 LR:-104.7 LO:104.7);ALT=C[chr1:246350043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246093241	+	chr1	246382744	+	.	0	20	649899_1	49.0	.	EVDNC=ASSMB;HOMSEQ=TCACCT;MAPQ=60;MATEID=649899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246372001_246397001_16C;SPAN=289503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:61 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:20 DR:0 LR:-49.49 LO:50.39);ALT=T[chr1:246382744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246518397	+	chr1	246670355	+	.	0	11	650981_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=650981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246666001_246691001_73C;SPAN=151958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:11 DR:0 LR:-26.02 LO:26.98);ALT=C[chr1:246670355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246729965	+	chr1	246754812	+	.	99	23	651890_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=651890_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_246715001_246740001_455C;SPAN=24847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:73 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:23 DR:99 LR:-359.8 LO:359.8);ALT=G[chr1:246754812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246733292	+	chr1	246754812	+	.	20	11	651948_1	53.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=651948_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_1_246739501_246764501_342C;SPAN=21520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:82 GQ:53.9 PL:[53.9, 0.0, 143.0] SR:11 DR:20 LR:-53.71 LO:56.04);ALT=G[chr1:246754812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	128868962	+	chr1	246806193	+	.	12	0	4445882_1	21.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4445882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:246806193(-)-9:128868962(+)__9_128845501_128870501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:0 DR:12 LR:-21.73 LO:26.64);ALT=]chr9:128868962]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr1	246887915	+	chr1	246890193	+	.	0	59	651632_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=651632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246886501_246911501_383C;SPAN=2278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:110 GQ:99 PL:[164.9, 0.0, 102.2] SR:59 DR:0 LR:-165.8 LO:165.8);ALT=G[chr1:246890193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246890306	+	chr1	246899277	+	.	0	17	651637_1	27.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=651637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246886501_246911501_56C;SPAN=8971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:105 GQ:27.8 PL:[27.8, 0.0, 225.8] SR:17 DR:0 LR:-27.67 LO:36.79);ALT=A[chr1:246899277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	246929442	+	chr1	246930497	+	.	0	16	652141_1	20.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=652141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_246911001_246936001_379C;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:119 GQ:20.6 PL:[20.6, 0.0, 268.1] SR:16 DR:0 LR:-20.58 LO:33.22);ALT=G[chr1:246930497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	247105771	-	chr7	124779379	+	.	29	0	3567703_1	89.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=3567703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:247105771(-)-7:124779379(-)__7_124778501_124803501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:35 GQ:2.7 PL:[89.1, 2.7, 0.0] SR:0 DR:29 LR:-91.93 LO:91.93);ALT=[chr7:124779379[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr1	247850475	+	chr1	247856516	+	.	100	60	655719_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=GAAAAGAAAGATC;MAPQ=60;MATEID=655719_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_247842001_247867001_25C;SPAN=6041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:49 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:60 DR:100 LR:-389.5 LO:389.5);ALT=C[chr1:247856516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	248051492	+	chr1	248057639	+	.	111	60	656454_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCATGTATTTATTT;MAPQ=60;MATEID=656454_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_1_248038001_248063001_31C;SPAN=6147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:42 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:60 DR:111 LR:-406.0 LO:406.0);ALT=T[chr1:248057639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	248839556	+	chr1	248840901	+	.	0	49	658794_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AAATTTAC;MAPQ=60;MATEID=658794_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_1_248822001_248847001_69C;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:31 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:49 DR:0 LR:-145.2 LO:145.2);ALT=C[chr1:248840901[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	265011	+	chr2	271865	+	.	79	11	660263_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTAA;MAPQ=60;MATEID=660263_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_245001_270001_312C;SPAN=6854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:55 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:11 DR:79 LR:-237.7 LO:237.7);ALT=A[chr2:271865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	669852	+	chr2	677289	+	CCAGTTCATCGCAGCCGCCTCATTGATGTATTCAGCACAGTAGACTAAGATGACTAGACACAGAAAGTGCCCGATCTGTAGTCTGTAGCTTCGGGAGGACAAGCAGGTGAGGAGCACGCAGAGCGCGTGGAAGGTGGCCAGCCCCATGAGCCAGGGCTCAGTCCAGTCCGTCTG	0	25	661440_1	64.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCAGTTCATCGCAGCCGCCTCATTGATGTATTCAGCACAGTAGACTAAGATGACTAGACACAGAAAGTGCCCGATCTGTAGTCTGTAGCTTCGGGAGGACAAGCAGGTGAGGAGCACGCAGAGCGCGTGGAAGGTGGCCAGCCCCATGAGCCAGGGCTCAGTCCAGTCCGTCTG;MAPQ=60;MATEID=661440_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_661501_686501_308C;SPAN=7437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:66 GQ:64.7 PL:[64.7, 0.0, 94.4] SR:25 DR:0 LR:-64.64 LO:64.97);ALT=T[chr2:677289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	675660	+	chr2	677344	+	.	21	0	661450_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=661450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:675660(+)-2:677344(-)__2_661501_686501D;SPAN=1684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:72 GQ:50 PL:[50.0, 0.0, 122.6] SR:0 DR:21 LR:-49.81 LO:51.6);ALT=G[chr2:677344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	1536483	+	chr2	1529454	+	.	0	26	664242_1	75.0	.	EVDNC=ASSMB;HOMSEQ=CCCCAAATCCCCC;MAPQ=60;MATEID=664242_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_2_1519001_1544001_147C;SPAN=7029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:37 GQ:13.1 PL:[75.8, 0.0, 13.1] SR:26 DR:0 LR:-78.22 LO:78.22);ALT=]chr2:1536483]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	1706799	+	chr2	1708435	+	.	9	0	663728_1	24.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=663728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:1706799(+)-2:1708435(-)__2_1690501_1715501D;SPAN=1636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:21 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.02 LO:24.03);ALT=G[chr2:1708435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	2577361	+	chr2	2576192	+	.	28	0	666407_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=666407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:2576192(-)-2:2577361(+)__2_2572501_2597501D;SPAN=1169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:28 DP:1259 GQ:99 PL:[0.0, 248.3, 3555.0] SR:0 DR:28 LR:248.7 LO:35.65);ALT=]chr2:2577361]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	2785137	+	chr2	2783804	+	.	14	0	666597_1	21.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=666597_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:2783804(-)-2:2785137(+)__2_2768501_2793501D;SPAN=1333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:0 DR:14 LR:-21.29 LO:29.89);ALT=]chr2:2785137]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	165894036	+	chr2	2973593	+	TTAGCTCCCACTTAAGTGAGAACATACGACATG	0	45	1075584_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TGGTTTTCCATTCCTGA;INSERTION=TTAGCTCCCACTTAAGTGAGAACATACGACATG;MAPQ=36;MATEID=1075584_2;MATENM=1;NM=0;NUMPARTS=4;SCTG=c_2_165889501_165914501_17C;SPAN=162920443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:23 GQ:12 PL:[132.0, 12.0, 0.0] SR:45 DR:0 LR:-132.0 LO:132.0);ALT=]chr2:165894036]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	3358407	+	chr2	3381418	+	.	0	11	668221_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=668221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3356501_3381501_243C;SPAN=23011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:97 GQ:10.1 PL:[10.1, 0.0, 224.6] SR:11 DR:0 LR:-10.03 LO:21.97);ALT=G[chr2:3381418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3383648	+	chr2	3391388	+	.	6	2	668048_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=668048_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3381001_3406001_265C;SPAN=7740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:2 DR:6 LR:1.547 LO:12.74);ALT=G[chr2:3391388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3504766	+	chr2	3517628	+	.	5	33	668437_1	96.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=668437_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3503501_3528501_22C;SPAN=12862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:82 GQ:96.8 PL:[96.8, 0.0, 100.1] SR:33 DR:5 LR:-96.62 LO:96.63);ALT=T[chr2:3517628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3504815	+	chr2	3523170	+	.	21	0	668438_1	45.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=668438_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:3504815(+)-2:3523170(-)__2_3503501_3528501D;SPAN=18355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:88 GQ:45.5 PL:[45.5, 0.0, 167.6] SR:0 DR:21 LR:-45.48 LO:49.44);ALT=G[chr2:3523170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3517749	+	chr2	3523139	+	.	0	40	668467_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=668467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3503501_3528501_90C;SPAN=5390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:84 GQ:92.9 PL:[109.4, 0.0, 92.9] SR:40 DR:0 LR:-109.3 LO:109.3);ALT=T[chr2:3523139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3579902	+	chr2	3581703	+	.	0	10	668509_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=668509_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3577001_3602001_258C;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:78 GQ:11.9 PL:[11.9, 0.0, 176.9] SR:10 DR:0 LR:-11.88 LO:20.54);ALT=T[chr2:3581703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3581846	+	chr2	3584312	+	.	20	7	668515_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=668515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3577001_3602001_61C;SPAN=2466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:83 GQ:47 PL:[47.0, 0.0, 152.6] SR:7 DR:20 LR:-46.83 LO:50.06);ALT=C[chr2:3584312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3593462	+	chr2	3595521	+	.	2	5	668553_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=668553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3577001_3602001_168C;SPAN=2059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:86 GQ:6.6 PL:[0.0, 6.6, 221.1] SR:5 DR:2 LR:6.795 LO:8.471);ALT=C[chr2:3595521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3604495	+	chr2	3605722	+	.	0	18	668710_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=668710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_3601501_3626501_70C;SPAN=1227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:86 GQ:36.2 PL:[36.2, 0.0, 171.5] SR:18 DR:0 LR:-36.12 LO:41.2);ALT=C[chr2:3605722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	3623018	+	chr17	26794855	+	.	30	0	6354006_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6354006_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:3623018(+)-17:26794855(-)__17_26778501_26803501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:30 DP:574 GQ:56.1 PL:[0.0, 56.1, 1505.0] SR:0 DR:30 LR:56.48 LO:49.41);ALT=G[chr17:26794855[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	3639922	-	chr16	31114886	+	.	6	19	6186437_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTCTCC;MAPQ=60;MATEID=6186437_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_16_31090501_31115501_105C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:50 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:19 DR:6 LR:-69.1 LO:69.1);ALT=[chr16:31114886[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	3688280	-	chr2	3689312	+	.	8	0	668933_1	2.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=668933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:3688280(-)-2:3689312(-)__2_3675001_3700001D;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=[chr2:3689312[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	4205269	-	chr2	4223479	+	CAT	19	22	670397_1	97.0	.	DISC_MAPQ=50;EVDNC=TSI_L;INSERTION=CAT;MAPQ=60;MATEID=670397_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_4189501_4214501_34C;SPAN=18210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:44 GQ:8 PL:[97.1, 0.0, 8.0] SR:22 DR:19 LR:-101.2 LO:101.2);ALT=[chr2:4223479[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	4205436	+	chr2	4212676	-	CAT	22	28	670399_1	99.0	.	DISC_MAPQ=51;EVDNC=TSI_L;HOMSEQ=CC;INSERTION=CAT;MAPQ=60;MATEID=670399_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_2_4189501_4214501_34C;SPAN=7240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:92 GQ:99 PL:[113.9, 0.0, 107.3] SR:28 DR:22 LR:-113.7 LO:113.7);ALT=C]chr2:4212676];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	4212676	+	chr2	4223479	+	CATAATTCTTCAATCTTTCATCGGTAGATTTTGGGATATAAGTAGAAAGCAAGGTGTTTTAACTAATGTCATATATCATAGAAAATAAAAGCAATATATTTATCCACTGCATTTAGAAGTATGAATGCTGGGGGGGGAGGAGCCAAGATGGCCGAATAGGAACAGCTC	0	46	670416_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CATAATTCTTCAATCTTTCATCGGTAGATTTTGGGATATAAGTAGAAAGCAAGGTGTTTTAACTAATGTCATATATCATAGAAAATAAAAGCAATATATTTATCCACTGCATTTAGAAGTATGAATGCTGGGGGGGGAGGAGCCAAGATGGCCGAATAGGAACAGCTC;MAPQ=60;MATEID=670416_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_4189501_4214501_34C;SPAN=10803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:45 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:46 DR:0 LR:-135.3 LO:135.3);ALT=G[chr2:4223479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	4781310	+	chr2	4787357	+	.	79	37	671921_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAGATACTGCA;MAPQ=60;MATEID=671921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_4777501_4802501_273C;SPAN=6047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:106 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:37 DR:79 LR:-312.5 LO:312.5);ALT=A[chr2:4787357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	7057754	+	chr2	7081077	+	.	8	11	676528_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=676528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_7080501_7105501_219C;SPAN=23323;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:57 GQ:37.4 PL:[37.4, 0.0, 100.1] SR:11 DR:8 LR:-37.37 LO:38.99);ALT=G[chr2:7081077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	7465154	+	chr12	123752727	+	.	11	0	5375570_1	26.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=5375570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:7465154(+)-12:123752727(-)__12_123749501_123774501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:0 DR:11 LR:-26.02 LO:26.98);ALT=C[chr12:123752727[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	26251322	+	chr11	64084948	+	.	19	0	4888395_1	41.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=4888395_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:26251322(+)-11:64084948(-)__11_64067501_64092501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:78 GQ:41.6 PL:[41.6, 0.0, 147.2] SR:0 DR:19 LR:-41.59 LO:44.92);ALT=G[chr11:64084948[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	26438045	+	chr2	26453059	+	.	0	14	725352_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=725352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_26435501_26460501_357C;SPAN=15014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:14 DR:0 LR:-18.58 LO:29.2);ALT=C[chr2:26453059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26455149	+	chr2	26457083	+	.	2	5	725417_1	3.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=725417_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_26435501_26460501_189C;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:5 DR:2 LR:-3.059 LO:13.4);ALT=T[chr2:26457083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26457223	+	chr2	26459723	+	.	2	16	725424_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=725424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_26435501_26460501_29C;SPAN=2500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:16 DR:2 LR:-32.87 LO:40.05);ALT=G[chr2:26459723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26459858	+	chr2	26461799	+	.	0	59	725438_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=725438_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_26460001_26485001_47C;SPAN=1941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:36 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:59 DR:0 LR:-174.9 LO:174.9);ALT=T[chr2:26461799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26459896	+	chr2	26467411	+	.	64	0	725439_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=725439_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:26459896(+)-2:26467411(-)__2_26460001_26485001D;SPAN=7515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:54 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=G[chr2:26467411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26467890	+	chr2	26486244	+	.	17	0	725971_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=725971_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:26467890(+)-2:26486244(-)__2_26484501_26509501D;SPAN=18354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:32 GQ:27.8 PL:[47.6, 0.0, 27.8] SR:0 DR:17 LR:-47.65 LO:47.65);ALT=G[chr2:26486244[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26467900	+	chr2	26477112	+	.	21	0	725479_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=725479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:26467900(+)-2:26477112(-)__2_26460001_26485001D;SPAN=9212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:57 GQ:53.9 PL:[53.9, 0.0, 83.6] SR:0 DR:21 LR:-53.88 LO:54.25);ALT=A[chr2:26477112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26507073	+	chr2	26508273	+	TGGTTTTTCTACCCATGTAGTTTTCTGCAAACCAATCAGAATCCATGGCTTTAAAATTTGCCAAAATCTGAC	2	12	726054_1	16.0	.	DISC_MAPQ=46;EVDNC=TSI_G;HOMSEQ=GACCAACCTGCAGCCAGTGGCTCCAAATGGGTGTCCCAGGGACAGAGATCCACCCCAGTTATTAAACTTCTCCAAAGGAGGCAATCCAACCTTGGTTTTTCTACCCATGTAGTTTTCTGCAAACCAATCAGAATCCATGGCTTTAAAATTTGCCAAAATCTGACCC;INSERTION=TGGTTTTTCTACCCATGTAGTTTTCTGCAAACCAATCAGAATCCATGGCTTTAAAATTTGCCAAAATCTGAC;MAPQ=60;MATEID=726054_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_26484501_26509501_350C;SECONDARY;SPAN=1200;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:97 GQ:16.7 PL:[16.7, 0.0, 218.0] SR:12 DR:2 LR:-16.63 LO:26.97);ALT=G[chr2:26508273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	26508440	+	chr2	26512783	+	.	6	10	726058_1	34.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=726058_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_26484501_26509501_252C;SPAN=4343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:55 GQ:34.7 PL:[34.7, 0.0, 97.4] SR:10 DR:6 LR:-34.61 LO:36.33);ALT=G[chr2:26512783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27435309	+	chr2	27438187	+	.	22	0	728180_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728180_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27435309(+)-2:27438187(-)__2_27415501_27440501D;SPAN=2878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:100 GQ:45.5 PL:[45.5, 0.0, 197.3] SR:0 DR:22 LR:-45.53 LO:50.89);ALT=G[chr2:27438187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27436167	+	chr2	27438188	+	.	2	49	728183_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=728183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27415501_27440501_265C;SPAN=2021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:117 GQ:99 PL:[133.4, 0.0, 149.9] SR:49 DR:2 LR:-133.4 LO:133.4);ALT=G[chr2:27438188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27535687	+	chr2	27545917	+	.	17	0	728691_1	39.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=728691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27535687(+)-2:27545917(-)__2_27513501_27538501D;SPAN=10230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:60 GQ:39.8 PL:[39.8, 0.0, 105.8] SR:0 DR:17 LR:-39.86 LO:41.51);ALT=G[chr2:27545917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27535688	+	chr2	27545340	+	.	8	0	728692_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27535688(+)-2:27545340(-)__2_27513501_27538501D;SPAN=9652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=G[chr2:27545340[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27535998	+	chr2	27545917	+	.	21	0	728695_1	59.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=728695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27535998(+)-2:27545917(-)__2_27513501_27538501D;SPAN=9919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:38 GQ:32.6 PL:[59.0, 0.0, 32.6] SR:0 DR:21 LR:-59.41 LO:59.41);ALT=T[chr2:27545917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27535999	+	chr2	27545344	+	.	10	0	728696_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728696_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27535999(+)-2:27545344(-)__2_27513501_27538501D;SPAN=9345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:38 GQ:22.7 PL:[22.7, 0.0, 68.9] SR:0 DR:10 LR:-22.72 LO:24.04);ALT=G[chr2:27545344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27593578	+	chr2	27595487	+	.	35	0	728801_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27593578(+)-2:27595487(-)__2_27587001_27612001D;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:0 DR:35 LR:-91.97 LO:92.16);ALT=T[chr2:27595487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27594210	+	chr2	27595488	+	.	0	52	728804_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=728804_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27587001_27612001_323C;SPAN=1278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:98 GQ:92.3 PL:[145.1, 0.0, 92.3] SR:52 DR:0 LR:-145.7 LO:145.7);ALT=G[chr2:27595488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27608748	+	chr2	27632169	+	TCTGTAGCTTGCCTTCCTTGTAGGCCTTCTGATCTTTGATGATATCAGGAAGATATTTGGCACAGTACAAGGCAACTTCCTCCCCTCCATGTCCATCGTAGACAGAAAACATGGCTGTCTCACTGTCCAGCTCAGGAATACAGTTGTGAGCAT	0	63	728855_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TCTGTAGCTTGCCTTCCTTGTAGGCCTTCTGATCTTTGATGATATCAGGAAGATATTTGGCACAGTACAAGGCAACTTCCTCCCCTCCATGTCCATCGTAGACAGAAAACATGGCTGTCTCACTGTCCAGCTCAGGAATACAGTTGTGAGCAT;MAPQ=60;MATEID=728855_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_27587001_27612001_63C;SPAN=23421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:34 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:63 DR:0 LR:-184.8 LO:184.8);ALT=T[chr2:27632169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27610073	+	chr2	27632224	+	.	16	0	728984_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=728984_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27610073(+)-2:27632224(-)__2_27611501_27636501D;SPAN=22151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:75 GQ:32.6 PL:[32.6, 0.0, 148.1] SR:0 DR:16 LR:-32.5 LO:36.77);ALT=T[chr2:27632224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27651632	+	chr2	27656113	+	.	39	0	729136_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=729136_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27651632(+)-2:27656113(-)__2_27636001_27661001D;SPAN=4481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:76 GQ:75.2 PL:[108.2, 0.0, 75.2] SR:0 DR:39 LR:-108.4 LO:108.4);ALT=A[chr2:27656113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27658094	+	chr2	27659619	+	.	2	6	729154_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=729154_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27636001_27661001_355C;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:6 DR:2 LR:3.764 LO:10.62);ALT=G[chr2:27659619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27806032	+	chr2	27820933	+	.	8	0	729931_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=729931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27806032(+)-2:27820933(-)__2_27807501_27832501D;SPAN=14901;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=T[chr2:27820933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27885149	+	chr2	27886195	+	.	5	6	729745_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=729745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27881001_27906001_184C;SPAN=1046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:73 GQ:13.4 PL:[13.4, 0.0, 161.9] SR:6 DR:5 LR:-13.23 LO:20.85);ALT=C[chr2:27886195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27994666	+	chr2	28002300	+	TTGCCAAGAGCAAGTCAAA	7	8	730463_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=TTGCCAAGAGCAAGTCAAA;MAPQ=60;MATEID=730463_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27979001_28004001_328C;SPAN=7634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:15 DP:221 GQ:10 PL:[0.0, 10.0, 554.5] SR:8 DR:7 LR:10.36 LO:26.45);ALT=T[chr2:28002300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27995247	+	chr2	27997290	+	.	25	0	730464_1	58.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=730464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:27995247(+)-2:27997290(-)__2_27979001_28004001D;SPAN=2043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:89 GQ:58.4 PL:[58.4, 0.0, 157.4] SR:0 DR:25 LR:-58.41 LO:60.94);ALT=G[chr2:27997290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27995252	+	chr2	28002300	+	TTGCCAAGAGCAAGTCAAA	148	7	730465_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTGCCAAGAGCAAGTCAAA;MAPQ=60;MATEID=730465_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_27979001_28004001_56C;SPAN=7048;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:133 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:7 DR:148 LR:-448.9 LO:448.9);ALT=G[chr2:28002300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	27997397	+	chr2	28002299	+	.	0	60	730467_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=730467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_27979001_28004001_343C;SPAN=4902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:138 GQ:99 PL:[160.7, 0.0, 173.9] SR:60 DR:0 LR:-160.7 LO:160.7);ALT=G[chr2:28002299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28081440	+	chr2	28113124	+	.	2	3	730562_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=730562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_28101501_28126501_186C;SPAN=31684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:50 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:3 DR:2 LR:-2.959 LO:9.695);ALT=T[chr2:28113124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28113759	+	chr2	28117396	+	.	33	0	730591_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=730591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:28113759(+)-2:28117396(-)__2_28101501_28126501D;SPAN=3637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:86 GQ:85.7 PL:[85.7, 0.0, 122.0] SR:0 DR:33 LR:-85.63 LO:86.0);ALT=G[chr2:28117396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28113768	+	chr2	28152697	+	.	9	0	730648_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=730648_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:28113768(+)-2:28152697(-)__2_28150501_28175501D;SPAN=38929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=A[chr2:28152697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28115315	+	chr2	28117398	+	.	0	7	730597_1	2.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=730597_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_2_28101501_28126501_227C;SPAN=2083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:7 DR:0 LR:-2.246 LO:13.27);ALT=G[chr2:28117398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28115315	+	chr2	28152698	+	TGGTGATTTACAAGTCAAGTTAAAATGTCCCCAGAAGTGGCCTTGAACCGAATATCTCCAATGCTCTCCCCTTTCATATCTAGCGTGGTCCGGAATGGAAAAGTGGGACTGGATGCTACAAACTGTTTGAGGATAACTGACTTAAAATCTG	0	25	730598_1	75.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TGGTGATTTACAAGTCAAGTTAAAATGTCCCCAGAAGTGGCCTTGAACCGAATATCTCCAATGCTCTCCCCTTTCATATCTAGCGTGGTCCGGAATGGAAAAGTGGGACTGGATGCTACAAACTGTTTGAGGATAACTGACTTAAAATCTG;MAPQ=60;MATEID=730598_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_28101501_28126501_227C;SPAN=37383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:30 GQ:1.5 PL:[75.9, 1.5, 0.0] SR:25 DR:0 LR:-79.42 LO:79.42);ALT=G[chr2:28152698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28627225	+	chr2	28631624	+	.	7	4	731966_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=731966_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_2_28616001_28641001_268C;SPAN=4399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:4 DR:7 LR:-5.276 LO:15.61);ALT=G[chr2:28631624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28975042	+	chr2	28999716	+	.	14	7	733131_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=733131_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_28983501_29008501_211C;SPAN=24674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:45 GQ:47.3 PL:[47.3, 0.0, 60.5] SR:7 DR:14 LR:-47.23 LO:47.34);ALT=G[chr2:28999716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28999849	+	chr2	29004604	+	AGATATTCATGGACAGTATACAGATTTACTGAGATTATTTGAATATGGAGGTTTCCCACCAGAAGCCAACTATCTTTTCTTAGGAGATTATGTGGACAGAGGAAAGCAGTCTTTGGAAACCATTTGTTTGCTATTGGCTTATAAAATCAAATATCCAGAGAACTTCTTTCTCTTAAGAGGAAACCATGAGTGTGCTAGCATCAATCGCATTTATGGATTCTATGATGAAT	0	11	733188_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AGATATTCATGGACAGTATACAGATTTACTGAGATTATTTGAATATGGAGGTTTCCCACCAGAAGCCAACTATCTTTTCTTAGGAGATTATGTGGACAGAGGAAAGCAGTCTTTGGAAACCATTTGTTTGCTATTGGCTTATAAAATCAAATATCCAGAGAACTTCTTTCTCTTAAGAGGAAACCATGAGTGTGCTAGCATCAATCGCATTTATGGATTCTATGATGAAT;MAPQ=60;MATEID=733188_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_28983501_29008501_164C;SPAN=4755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:71 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:11 DR:0 LR:-17.08 LO:23.58);ALT=G[chr2:29004604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	28999849	+	chr2	29001674	+	.	4	4	733187_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=733187_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_2_28983501_29008501_164C;SPAN=1825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:4 DR:4 LR:-7.985 LO:16.11);ALT=G[chr2:29001674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	29011677	+	chr2	29016726	+	.	2	4	733056_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGGT;MAPQ=60;MATEID=733056_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_29008001_29033001_177C;SPAN=5049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:78 GQ:1.2 PL:[0.0, 1.2, 191.4] SR:4 DR:2 LR:1.326 LO:10.92);ALT=T[chr2:29016726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	29016863	+	chr2	29022063	+	.	3	3	733075_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=733075_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_29008001_29033001_177C;SPAN=5200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:83 GQ:2.4 PL:[0.0, 2.4, 204.6] SR:3 DR:3 LR:2.681 LO:10.75);ALT=G[chr2:29022063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	29117790	+	chr2	29124851	+	.	0	10	733247_1	11.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=733247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_29106001_29131001_45C;SPAN=7061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:0 LR:-11.34 LO:20.42);ALT=G[chr2:29124851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	57976654	+	chr2	30294295	+	.	2	3	736526_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGAG;MAPQ=60;MATEID=736526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_30282001_30307001_56C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:48 GQ:3.5 PL:[3.5, 0.0, 112.4] SR:3 DR:2 LR:-3.501 LO:9.789);ALT=]chr8:57976654]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	30369930	+	chr2	30379493	+	.	11	16	736716_1	62.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=736716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_30355501_30380501_59C;SPAN=9563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:101 GQ:62 PL:[62.0, 0.0, 180.8] SR:16 DR:11 LR:-61.76 LO:65.12);ALT=T[chr2:30379493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	30369956	+	chr2	30378726	+	.	82	0	736719_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=736719_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:30369956(+)-2:30378726(-)__2_30355501_30380501D;SPAN=8770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:69 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=G[chr2:30378726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	30369965	+	chr2	30381481	+	.	28	0	736821_1	78.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=736821_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:30369965(+)-2:30381481(-)__2_30380001_30405001D;SPAN=11516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:52 GQ:45.5 PL:[78.5, 0.0, 45.5] SR:0 DR:28 LR:-78.73 LO:78.73);ALT=G[chr2:30381481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	30379660	+	chr2	30381483	+	.	0	36	736822_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=736822_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_30380001_30405001_194C;SPAN=1823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:53 GQ:22.1 PL:[104.6, 0.0, 22.1] SR:36 DR:0 LR:-107.3 LO:107.3);ALT=T[chr2:30381483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41238369	+	chr2	41250294	+	.	50	32	764464_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGA;MAPQ=60;MATEID=764464_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41233501_41258501_84C;SPAN=11925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:40 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:32 DR:50 LR:-204.7 LO:204.7);ALT=A[chr2:41250294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41775966	+	chr2	41781284	+	G	57	55	765669_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=765669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41772501_41797501_165C;SPAN=5318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:25 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:55 DR:57 LR:-267.4 LO:267.4);ALT=T[chr2:41781284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	41973156	+	chr2	41975866	+	.	79	54	766256_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAACCTCACATGC;MAPQ=60;MATEID=766256_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_41968501_41993501_127C;SPAN=2710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:46 GQ:27 PL:[297.0, 27.0, 0.0] SR:54 DR:79 LR:-297.1 LO:297.1);ALT=C[chr2:41975866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42052666	+	chr4	66413930	+	.	42	0	766432_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=766432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:42052666(+)-4:66413930(-)__2_42042001_42067001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:39 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=A[chr4:66413930[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	42217992	-	chr2	42219115	+	.	8	0	766820_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=766820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:42217992(-)-2:42219115(-)__2_42213501_42238501D;SPAN=1123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=[chr2:42219115[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	42346259	+	chr2	42347319	+	TGTA	32	20	767122_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTA;MAPQ=60;MATEID=767122_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_42336001_42361001_22C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:59 GQ:36.8 PL:[106.1, 0.0, 36.8] SR:20 DR:32 LR:-108.0 LO:108.0);ALT=C[chr2:42347319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42578501	+	chr2	42580352	+	.	5	101	767834_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=767834_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_42556501_42581501_12C;SPAN=1851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:132 GQ:4.1 PL:[314.3, 0.0, 4.1] SR:101 DR:5 LR:-332.3 LO:332.3);ALT=T[chr2:42580352[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42578554	+	chr2	42588232	+	.	62	0	767923_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=767923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:42578554(+)-2:42588232(-)__2_42581001_42606001D;SPAN=9678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:61 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:0 DR:62 LR:-181.5 LO:181.5);ALT=T[chr2:42588232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	42580486	+	chr2	42588229	+	.	165	41	767924_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=767924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_42581001_42606001_294C;SPAN=7743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:59 GQ:46 PL:[505.0, 46.0, 0.0] SR:41 DR:165 LR:-505.0 LO:505.0);ALT=G[chr2:42588229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	43200153	+	chr2	43207423	+	.	0	13	769918_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=769918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_43193501_43218501_182C;SPAN=7270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:13 DR:0 LR:-20.7 LO:28.0);ALT=G[chr2:43207423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	43228621	+	chr2	43231019	+	.	5	16	770267_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TCACC;MAPQ=60;MATEID=770267_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_2_43218001_43243001_42C;SPAN=2398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:80 GQ:37.7 PL:[37.7, 0.0, 156.5] SR:16 DR:5 LR:-37.74 LO:41.84);ALT=C[chr2:43231019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	43228622	+	chr2	43233177	+	.	20	3	770269_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=770269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_43218001_43243001_257C;SPAN=4555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:92 GQ:41.3 PL:[41.3, 0.0, 179.9] SR:3 DR:20 LR:-41.1 LO:46.15);ALT=T[chr2:43233177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	43231121	+	chr2	43233288	+	.	13	0	770281_1	19.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=770281_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:43231121(+)-2:43233288(-)__2_43218001_43243001D;SPAN=2167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:0 DR:13 LR:-19.34 LO:27.64);ALT=G[chr2:43233288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	44117016	+	chr2	44121684	+	.	4	4	772528_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=772528_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_44100001_44125001_87C;SPAN=4668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:4 DR:4 LR:-10.42 LO:16.64);ALT=C[chr2:44121684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	44169016	-	chr2	44170024	+	.	3	3	772582_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AATTAAAATAAAATAAAA;MAPQ=60;MATEID=772582_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_44149001_44174001_42C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:63 GQ:2.9 PL:[2.9, 0.0, 148.1] SR:3 DR:3 LR:-2.738 LO:11.5);ALT=[chr2:44170024[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	44209621	+	chr2	44223041	+	.	11	0	772950_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=772950_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:44209621(+)-2:44223041(-)__2_44222501_44247501D;SPAN=13420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:0 DR:11 LR:-23.31 LO:25.67);ALT=G[chr2:44223041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	44429185	+	chr2	44436347	+	.	0	8	773598_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=773598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_44418501_44443501_143C;SPAN=7162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:80 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:8 DR:0 LR:-4.734 LO:15.51);ALT=G[chr2:44436347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	44589286	+	chr2	44599853	+	.	9	8	774113_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=774113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_44565501_44590501_357C;SPAN=10567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:47 GQ:33.5 PL:[33.5, 0.0, 79.7] SR:8 DR:9 LR:-33.48 LO:34.55);ALT=T[chr2:44599853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	46842307	+	chr2	46844105	+	.	15	0	779826_1	26.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=779826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:46842307(+)-2:46844105(-)__2_46819501_46844501D;SPAN=1798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:87 GQ:26 PL:[26.0, 0.0, 184.4] SR:0 DR:15 LR:-25.94 LO:32.91);ALT=G[chr2:46844105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	46844441	+	chr2	46845912	+	.	6	5	779833_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GTGA;MAPQ=60;MATEID=779833_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=AA;SCTG=c_2_46819501_46844501_340C;SPAN=1471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:52 GQ:5.9 PL:[5.9, 0.0, 118.1] SR:5 DR:6 LR:-5.718 LO:12.03);ALT=A[chr2:46845912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	46844474	+	chr2	46846761	+	.	11	0	779835_1	23.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=779835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:46844474(+)-2:46846761(-)__2_46819501_46844501D;SPAN=2287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:49 GQ:23 PL:[23.0, 0.0, 95.6] SR:0 DR:11 LR:-23.04 LO:25.56);ALT=T[chr2:46846761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	46844484	+	chr2	46850899	+	.	18	0	779836_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=779836_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:46844484(+)-2:46850899(-)__2_46819501_46844501D;SPAN=6415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:47 GQ:46.7 PL:[46.7, 0.0, 66.5] SR:0 DR:18 LR:-46.68 LO:46.89);ALT=T[chr2:46850899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47136319	+	chr2	47168711	+	.	8	3	780692_1	23.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=780692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_47162501_47187501_307C;SPAN=32392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:23 GQ:23.6 PL:[23.6, 0.0, 30.2] SR:3 DR:8 LR:-23.48 LO:23.56);ALT=G[chr2:47168711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47220053	+	chr2	47229437	+	GTTGATTGCACATAGGAGAGA	15	63	780920_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;INSERTION=GTTGATTGCACATAGGAGAGA;MAPQ=60;MATEID=780920_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_47211501_47236501_242C;SPAN=9384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:240 GQ:99 PL:[156.1, 0.0, 426.8] SR:63 DR:15 LR:-156.1 LO:163.1);ALT=T[chr2:47229437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47389538	+	chr2	47403588	+	.	22	0	781614_1	24.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=781614_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:47389538(+)-2:47403588(-)__2_47383001_47408001D;SPAN=14050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:179 GQ:24.1 PL:[24.1, 0.0, 410.3] SR:0 DR:22 LR:-24.13 LO:44.76);ALT=T[chr2:47403588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47389830	+	chr2	47403577	+	.	106	0	781617_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=781617_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:47389830(+)-2:47403577(-)__2_47383001_47408001D;SPAN=13747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:81 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=T[chr2:47403577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	47403577	-	chr10	71923415	+	.	54	0	781682_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=781682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:47403577(-)-10:71923415(-)__2_47383001_47408001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:45 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=[chr10:71923415[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	48398167	-	chr2	48399193	+	.	9	0	784491_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=784491_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:48398167(-)-2:48399193(-)__2_48387501_48412501D;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:116 GQ:1.5 PL:[0.0, 1.5, 283.8] SR:0 DR:9 LR:1.718 LO:16.41);ALT=[chr2:48399193[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	48541953	+	chr2	48573339	+	.	40	7	784914_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=784914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48559001_48584001_122C;SPAN=31386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:65 GQ:32 PL:[124.4, 0.0, 32.0] SR:7 DR:40 LR:-127.2 LO:127.2);ALT=G[chr2:48573339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	48541953	+	chr2	48555699	+	.	12	2	784868_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=784868_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48534501_48559501_34C;SPAN=13746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:63 GQ:29.3 PL:[29.3, 0.0, 121.7] SR:2 DR:12 LR:-29.15 LO:32.46);ALT=G[chr2:48555699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	48781852	+	chr2	48784868	+	.	60	37	785747_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAAGTGCAAAATTTTTT;MAPQ=60;MATEID=785747_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48779501_48804501_359C;SPAN=3016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:60 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:37 DR:60 LR:-217.9 LO:217.9);ALT=T[chr2:48784868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	48851192	+	chr2	48857953	+	.	49	45	785640_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=785640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_48853001_48878001_52C;SPAN=6761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:22 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:45 DR:49 LR:-221.2 LO:221.2);ALT=A[chr2:48857953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	58688499	-	chr5	140035412	+	.	9	0	808333_1	20.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=808333_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:58688499(-)-5:140035412(-)__2_58677501_58702501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=[chr5:140035412[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	63555285	+	chr2	63549348	+	.	13	0	821250_1	30.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=821250_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63549348(-)-2:63555285(+)__2_63553001_63578001D;SPAN=5937;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:45 GQ:30.8 PL:[30.8, 0.0, 77.0] SR:0 DR:13 LR:-30.72 LO:31.88);ALT=]chr2:63555285]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	63816215	+	chr2	63824529	+	.	23	0	821675_1	65.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=821675_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63816215(+)-2:63824529(-)__2_63822501_63847501D;SPAN=8314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:38 GQ:26 PL:[65.6, 0.0, 26.0] SR:0 DR:23 LR:-66.53 LO:66.53);ALT=G[chr2:63824529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	63816227	+	chr2	63821669	+	.	59	0	821676_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=821676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:63816227(+)-2:63821669(-)__2_63822501_63847501D;SPAN=5442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:0 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=T[chr2:63821669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	63822653	+	chr2	63824531	+	.	0	33	821678_1	85.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=821678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_63822501_63847501_302C;SPAN=1878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:88 GQ:85.1 PL:[85.1, 0.0, 128.0] SR:33 DR:0 LR:-85.09 LO:85.58);ALT=G[chr2:63824531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	63824710	+	chr2	63826302	+	.	5	3	821681_1	5.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=821681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_63822501_63847501_139C;SPAN=1592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:3 DR:5 LR:-5.818 LO:15.7);ALT=T[chr2:63826302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	64068366	+	chr2	64083437	+	.	12	11	822337_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAG;MAPQ=60;MATEID=822337_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_64067501_64092501_188C;SPAN=15071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:92 GQ:34.7 PL:[34.7, 0.0, 186.5] SR:11 DR:12 LR:-34.49 LO:40.6);ALT=G[chr2:64083437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	64083567	+	chr2	64084961	+	.	0	10	822384_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=822384_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_64067501_64092501_138C;SPAN=1394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:10 DR:0 LR:-9.169 LO:19.98);ALT=G[chr2:64084961[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	64114780	+	chr2	64117212	+	.	6	3	822573_1	12.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=AAGGT;MAPQ=60;MATEID=822573_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_64092001_64117001_120C;SPAN=2432;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:41 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:3 DR:6 LR:-12.0 LO:15.33);ALT=T[chr2:64117212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	64335514	+	chr2	64371214	+	.	0	8	823236_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=823236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_64361501_64386501_40C;SPAN=35700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:8 DR:0 LR:-15.57 LO:18.13);ALT=C[chr2:64371214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	64864010	+	chr2	64880754	+	.	10	10	824474_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=824474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_64876001_64901001_310C;SPAN=16744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:35 GQ:36.8 PL:[36.8, 0.0, 46.7] SR:10 DR:10 LR:-36.73 LO:36.82);ALT=C[chr2:64880754[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40615708	+	chr2	65138905	+	.	18	29	6816193_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6816193_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_19_40596501_40621501_116C;SECONDARY;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:25 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:29 DR:18 LR:-112.2 LO:112.2);ALT=]chr19:40615708]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	65331940	+	chr2	65357027	+	.	0	13	826470_1	30.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=826470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_65317001_65342001_385C;SPAN=25087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:45 GQ:30.8 PL:[30.8, 0.0, 77.0] SR:13 DR:0 LR:-30.72 LO:31.88);ALT=A[chr2:65357027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	76970645	+	chr2	65432202	+	.	20	0	4633850_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4633850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:65432202(-)-10:76970645(+)__10_76954501_76979501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:30 GQ:14.9 PL:[57.8, 0.0, 14.9] SR:0 DR:20 LR:-59.31 LO:59.31);ALT=]chr10:76970645]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	65455058	+	chr19	20369162	+	.	11	0	6762570_1	23.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6762570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:65455058(+)-19:20369162(-)__19_20359501_20384501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:0 DR:11 LR:-23.85 LO:25.91);ALT=C[chr19:20369162[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	65455061	+	chr2	65466984	+	.	20	0	826201_1	54.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=826201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:65455061(+)-2:65466984(-)__2_65464001_65489001D;SPAN=11923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:43 GQ:47.9 PL:[54.5, 0.0, 47.9] SR:0 DR:20 LR:-54.38 LO:54.38);ALT=G[chr2:65466984[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	32800610	+	chr2	68290075	+	.	8	0	4567402_1	13.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4567402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:68290075(-)-10:32800610(+)__10_32781001_32806001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=]chr10:32800610]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	68592526	+	chr2	68607458	+	.	96	19	834109_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=834109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_68600001_68625001_162C;SPAN=14932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:48 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:19 DR:96 LR:-300.4 LO:300.4);ALT=G[chr2:68607458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	68592560	+	chr2	68607853	+	.	29	0	834110_1	82.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=834110_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:68592560(+)-2:68607853(-)__2_68600001_68625001D;SPAN=15293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:50 GQ:39.2 PL:[82.1, 0.0, 39.2] SR:0 DR:29 LR:-83.01 LO:83.01);ALT=G[chr2:68607853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	68613818	+	chr2	68615519	+	.	5	8	834147_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=834147_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_68600001_68625001_288C;SPAN=1701;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:8 DR:5 LR:-3.158 LO:17.1);ALT=T[chr2:68615519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	68914913	+	chr5	64468037	-	.	28	0	2488549_1	89.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2488549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:68914913(+)-5:64468037(+)__5_64459501_64484501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:28 LR:-89.12 LO:89.12);ALT=A]chr5:64468037];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	69650851	+	chr2	69659034	+	.	0	15	836527_1	37.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=836527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_69653501_69678501_6C;SPAN=8183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:45 GQ:37.4 PL:[37.4, 0.0, 70.4] SR:15 DR:0 LR:-37.32 LO:37.92);ALT=T[chr2:69659034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	69650888	+	chr2	69664506	+	.	11	0	836747_1	24.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=836747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:69650888(+)-2:69664506(-)__2_69629001_69654001D;SPAN=13618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:43 GQ:24.8 PL:[24.8, 0.0, 77.6] SR:0 DR:11 LR:-24.66 LO:26.28);ALT=A[chr2:69664506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	69659138	+	chr2	69664491	+	.	14	3	836553_1	23.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=836553_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_69653501_69678501_145C;SPAN=5353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:3 DR:14 LR:-23.73 LO:30.57);ALT=C[chr2:69664491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	69969349	+	chr2	70015183	+	.	27	0	837558_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=837558_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:69969349(+)-2:70015183(-)__2_69996501_70021501D;SPAN=45834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:44 GQ:27.8 PL:[77.3, 0.0, 27.8] SR:0 DR:27 LR:-78.37 LO:78.37);ALT=C[chr2:70015183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	69969349	+	chr2	70031662	+	.	34	0	837624_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=837624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:69969349(+)-2:70031662(-)__2_70021001_70046001D;SPAN=62313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:47 GQ:13.7 PL:[99.5, 0.0, 13.7] SR:0 DR:34 LR:-103.1 LO:103.1);ALT=C[chr2:70031662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70031760	+	chr2	70033516	+	.	0	17	837658_1	32.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=837658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_70021001_70046001_136C;SPAN=1756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:89 GQ:32 PL:[32.0, 0.0, 183.8] SR:17 DR:0 LR:-32.01 LO:38.15);ALT=G[chr2:70033516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70047954	+	chr2	70052586	+	.	3	7	837727_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=837727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_70045501_70070501_188C;SPAN=4632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:7 DR:3 LR:-6.089 LO:15.75);ALT=G[chr2:70052586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70121190	+	chr2	70123565	+	.	9	0	838047_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=838047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70121190(+)-2:70123565(-)__2_70119001_70144001D;SPAN=2375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:0 DR:9 LR:-5.868 LO:17.54);ALT=G[chr2:70123565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70121198	+	chr2	70122224	+	.	14	0	838048_1	19.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=838048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70121198(+)-2:70122224(-)__2_70119001_70144001D;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:98 GQ:19.7 PL:[19.7, 0.0, 217.7] SR:0 DR:14 LR:-19.66 LO:29.47);ALT=G[chr2:70122224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70122346	+	chr2	70124508	+	ATCTCCAAGACGACATAGATCCACATCTCCTTCCCCTTCTCGACTGAAAGAAAGAAGAGATGAGGAAAAGAAAGAAACAAAAGAAACAAAGAGCAAAGAACGGCAGATTACT	0	23	838051_1	53.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATCTCCAAGACGACATAGATCCACATCTCCTTCCCCTTCTCGACTGAAAGAAAGAAGAGATGAGGAAAAGAAAGAAACAAAAGAAACAAAGAGCAAAGAACGGCAGATTACT;MAPQ=60;MATEID=838051_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_70119001_70144001_0C;SPAN=2162;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:85 GQ:53 PL:[53.0, 0.0, 152.0] SR:23 DR:0 LR:-52.89 LO:55.62);ALT=G[chr2:70124508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70162597	+	chr2	70164365	+	.	3	3	838014_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=838014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_70143501_70168501_89C;SPAN=1768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:81 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:3 DR:3 LR:5.44 LO:8.605);ALT=G[chr2:70164365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70451761	+	chr2	70454867	+	.	0	7	838891_1	6.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=838891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_70437501_70462501_79C;SPAN=3106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:61 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:7 DR:0 LR:-6.581 LO:14.02);ALT=T[chr2:70454867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70457986	+	chr2	70475537	+	ATCCATAATCATTTTGCAGTTTTTACAAGGTCCAATCTGGCTAAAGAGTTGCAGAATTAGAGCTTCTGTCACATCTCTGGAAAGGTTACCGACGTAT	6	20	839080_1	58.0	.	DISC_MAPQ=60;EVDNC=TSI_G;INSERTION=ATCCATAATCATTTTGCAGTTTTTACAAGGTCCAATCTGGCTAAAGAGTTGCAGAATTAGAGCTTCTGTCACATCTCTGGAAAGGTTACCGACGTAT;MAPQ=60;MATEID=839080_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_70462001_70487001_128C;SPAN=17551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:53 GQ:58.4 PL:[58.4, 0.0, 68.3] SR:20 DR:6 LR:-58.26 LO:58.33);ALT=T[chr2:70475537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70463307	+	chr2	70475537	+	.	9	15	839085_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=839085_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_70462001_70487001_128C;SPAN=12230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:96 GQ:36.8 PL:[36.8, 0.0, 195.2] SR:15 DR:9 LR:-36.71 LO:42.96);ALT=T[chr2:70475537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70494166	+	chr6	31297451	-	.	16	0	2773970_1	45.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2773970_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70494166(+)-6:31297451(+)__6_31286501_31311501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:28 GQ:22.1 PL:[45.2, 0.0, 22.1] SR:0 DR:16 LR:-45.63 LO:45.63);ALT=G]chr6:31297451];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	70524612	+	chr2	70527971	+	.	0	44	839635_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=839635_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_70511001_70536001_278C;SPAN=3359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:105 GQ:99 PL:[116.9, 0.0, 136.7] SR:44 DR:0 LR:-116.8 LO:116.9);ALT=G[chr2:70527971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70524629	+	chr2	70529096	+	.	12	0	839636_1	7.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=839636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70524629(+)-2:70529096(-)__2_70511001_70536001D;SPAN=4467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:118 GQ:7.7 PL:[7.7, 0.0, 278.3] SR:0 DR:12 LR:-7.643 LO:23.36);ALT=C[chr2:70529096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	70662448	+	chr2	70661187	+	.	50	0	840263_1	99.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=840263_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:70661187(-)-2:70662448(+)__2_70658001_70683001D;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:78 GQ:44.9 PL:[143.9, 0.0, 44.9] SR:0 DR:50 LR:-146.7 LO:146.7);ALT=]chr2:70662448]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	71295863	+	chr2	71297869	+	.	8	0	841788_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=841788_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:71295863(+)-2:71297869(-)__2_71295001_71320001D;SPAN=2006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:0 DR:8 LR:0.6845 LO:14.7);ALT=G[chr2:71297869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	71357859	+	chr2	71360027	+	.	13	0	841547_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=841547_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:71357859(+)-2:71360027(-)__2_71344001_71369001D;SPAN=2168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:0 DR:13 LR:-20.7 LO:28.0);ALT=A[chr2:71360027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	71909807	+	chr2	71913583	+	.	5	5	842979_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=842979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_71907501_71932501_56C;SPAN=3776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:5 DR:5 LR:-5.326 LO:17.45);ALT=G[chr2:71913583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73460256	-	chr3	37017850	+	.	13	0	1354088_1	24.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1354088_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:73460256(-)-3:37017850(-)__3_36995001_37020001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:68 GQ:24.5 PL:[24.5, 0.0, 140.0] SR:0 DR:13 LR:-24.49 LO:29.18);ALT=[chr3:37017850[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	73461512	+	chr2	73466770	+	.	50	8	846958_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=846958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_73451001_73476001_311C;SPAN=5258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:108 GQ:99 PL:[145.7, 0.0, 116.0] SR:8 DR:50 LR:-145.9 LO:145.9);ALT=G[chr2:73466770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73461550	+	chr2	73467562	+	.	31	0	846961_1	77.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=846961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:73461550(+)-2:73467562(-)__2_73451001_73476001D;SPAN=6012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:93 GQ:77.3 PL:[77.3, 0.0, 146.6] SR:0 DR:31 LR:-77.14 LO:78.38);ALT=C[chr2:73467562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73467673	+	chr2	73470130	+	.	0	11	846969_1	16.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=846969_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_73451001_73476001_90C;SPAN=2457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:11 DR:0 LR:-15.99 LO:23.29);ALT=T[chr2:73470130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73478561	+	chr2	73479766	+	.	6	13	847027_1	42.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=847027_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_73475501_73500501_186C;SPAN=1205;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:76 GQ:42.2 PL:[42.2, 0.0, 141.2] SR:13 DR:6 LR:-42.13 LO:45.17);ALT=G[chr2:73479766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73957158	+	chr2	73961556	+	TTTTGACTTCTGTAATATTCATTATTTCAGGAAGATTTTTCAGAGAAACCTGATGACCTTCTACTTGAGATATTAGGTATTCTTGATTTATTTGTTTTTCTCCCTCTTCAATGTAAACAATTAGAATTGAAGTGTCATTTGCTGAGATACCAAATTTTTTCAAAGCCTCTGAAATATTGTTATTTGGGGAAAGGTTGAAAATAATTTCAGTAGATAGAGTTCTTGTCTTCATTTTTCCCAGTTTGTAGAGGTGAACTGCTTTGTTTGCTGCCACAAGTATCTGAAATGGATCAACAAT	0	36	848404_1	98.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTTTGACTTCTGTAATATTCATTATTTCAGGAAGATTTTTCAGAGAAACCTGATGACCTTCTACTTGAGATATTAGGTATTCTTGATTTATTTGTTTTTCTCCCTCTTCAATGTAAACAATTAGAATTGAAGTGTCATTTGCTGAGATACCAAATTTTTTCAAAGCCTCTGAAATATTGTTATTTGGGGAAAGGTTGAAAATAATTTCAGTAGATAGAGTTCTTGTCTTCATTTTTCCCAGTTTGTAGAGGTGAACTGCTTTGTTTGCTGCCACAAGTATCTGAAATGGATCAACAAT;MAPQ=60;MATEID=848404_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_2_73941001_73966001_58C;SPAN=4398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:77 GQ:88.1 PL:[98.0, 0.0, 88.1] SR:36 DR:0 LR:-98.0 LO:98.0);ALT=T[chr2:73961556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73957863	+	chr2	73959290	+	.	0	13	848407_1	26.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=848407_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_2_73941001_73966001_58C;SPAN=1427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:59 GQ:26.9 PL:[26.9, 0.0, 116.0] SR:13 DR:0 LR:-26.93 LO:30.08);ALT=T[chr2:73959290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	73959454	+	chr2	73961668	+	.	11	0	848410_1	11.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=848410_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:73959454(+)-2:73961668(-)__2_73941001_73966001D;SPAN=2214;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:0 DR:11 LR:-11.39 LO:22.24);ALT=C[chr2:73961668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74005505	+	chr2	74006999	+	.	0	6	848461_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=848461_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_73990001_74015001_289C;SPAN=1494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:79 GQ:1.5 PL:[0.0, 1.5, 194.7] SR:6 DR:0 LR:1.597 LO:10.88);ALT=T[chr2:74006999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74058187	+	chr2	74071940	+	.	0	17	848994_1	47.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=848994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74063501_74088501_67C;SPAN=13753;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:33 GQ:30.8 PL:[47.3, 0.0, 30.8] SR:17 DR:0 LR:-47.31 LO:47.31);ALT=G[chr2:74071940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74154100	+	chr2	74185270	+	.	9	0	849411_1	15.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=849411_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:74154100(+)-2:74185270(-)__2_74137001_74162001D;SPAN=31170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:0 DR:9 LR:-15.08 LO:19.6);ALT=C[chr2:74185270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74154179	+	chr2	74166036	+	.	0	20	849413_1	48.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=849413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74137001_74162001_71C;SPAN=11857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:64 GQ:48.8 PL:[48.8, 0.0, 104.9] SR:20 DR:0 LR:-48.68 LO:49.87);ALT=G[chr2:74166036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74154180	+	chr2	74173845	+	.	57	39	849414_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=849414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74137001_74162001_15C;SPAN=19665;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:63 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:39 DR:57 LR:-221.2 LO:221.2);ALT=G[chr2:74173845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74166150	+	chr2	74173846	+	.	0	7	849216_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=849216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74161501_74186501_120C;SPAN=7696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:108 GQ:6 PL:[0.0, 6.0, 273.9] SR:7 DR:0 LR:6.153 LO:12.2);ALT=G[chr2:74173846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74174034	+	chr2	74185271	+	.	0	10	849241_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=849241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74161501_74186501_90C;SPAN=11237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:10 DR:0 LR:-7.543 LO:19.68);ALT=G[chr2:74185271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74362787	+	chr2	74372315	+	.	0	10	849808_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=849808_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74357501_74382501_133C;SPAN=9528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:10 DR:0 LR:-13.5 LO:20.92);ALT=T[chr2:74372315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74362828	+	chr2	74374947	+	.	12	0	849809_1	15.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=849809_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:74362828(+)-2:74374947(-)__2_74357501_74382501D;SPAN=12119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:89 GQ:15.5 PL:[15.5, 0.0, 200.3] SR:0 DR:12 LR:-15.5 LO:24.93);ALT=T[chr2:74374947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74372431	+	chr2	74374948	+	.	5	3	849833_1	0	.	DISC_MAPQ=25;EVDNC=ASDIS;HOMSEQ=C;MAPQ=19;MATEID=849833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74357501_74382501_164C;SPAN=2517;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:3 DR:5 LR:1.818 LO:12.7);ALT=C[chr2:74374948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74399879	+	chr2	74405788	+	.	0	10	850121_1	14.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=850121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74382001_74407001_372C;SPAN=5909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:10 DR:0 LR:-13.77 LO:20.98);ALT=G[chr2:74405788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74425869	+	chr2	74432831	+	.	27	20	850265_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=850265_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74406501_74431501_184C;SPAN=6962;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:30 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:20 DR:27 LR:-138.6 LO:138.6);ALT=G[chr2:74432831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74425870	+	chr2	74428508	+	.	10	4	850267_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=850267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74406501_74431501_314C;SPAN=2638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:4 DR:10 LR:-14.05 LO:21.05);ALT=G[chr2:74428508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74590555	+	chr2	74592201	+	.	2	2	850617_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=850617_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_74578001_74603001_284C;SPAN=1646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:111 GQ:16.5 PL:[0.0, 16.5, 300.3] SR:2 DR:2 LR:16.87 LO:5.932);ALT=C[chr2:74592201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	74605406	+	chr2	74618920	+	.	19	0	850675_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=850675_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:74605406(+)-2:74618920(-)__2_74602501_74627501D;SPAN=13514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:87 GQ:39.2 PL:[39.2, 0.0, 171.2] SR:0 DR:19 LR:-39.15 LO:43.89);ALT=G[chr2:74618920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	75186552	+	chr2	75196534	+	ATAATGCAATAGAAGCTGTGGATGAATTTGCTTTTCTGGA	6	37	852291_1	99.0	.	DISC_MAPQ=47;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=ATAATGCAATAGAAGCTGTGGATGAATTTGCTTTTCTGGA;MAPQ=60;MATEID=852291_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_75166001_75191001_325C;SPAN=9982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:37 DR:6 LR:-125.4 LO:125.4);ALT=G[chr2:75196534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	75443089	+	chr2	77318914	-	.	9	0	857377_1	16.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=857377_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:75443089(+)-2:77318914(+)__2_77297501_77322501D;SPAN=1875825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-15.89 LO:19.85);ALT=C]chr2:77318914];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	75874347	+	chr2	75879265	+	.	0	11	853947_1	22.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=853947_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_75852001_75877001_94C;SPAN=4918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:50 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:11 DR:0 LR:-22.76 LO:25.45);ALT=T[chr2:75879265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	75878635	+	chr17	56429449	+	.	30	0	6446269_1	85.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6446269_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:75878635(+)-17:56429449(-)__17_56423501_56448501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:51 GQ:35.9 PL:[85.4, 0.0, 35.9] SR:0 DR:30 LR:-86.17 LO:86.17);ALT=A[chr17:56429449[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	76526512	+	chr2	76528894	+	.	48	40	855560_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTTTTCCATGTTTT;MAPQ=60;MATEID=855560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_76513501_76538501_253C;SPAN=2382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:34 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:40 DR:48 LR:-221.2 LO:221.2);ALT=T[chr2:76528894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	76773553	+	chr2	76775453	+	TTATTCTTTTA	0	23	856038_1	66.0	.	EVDNC=ASSMB;INSERTION=TTATTCTTTTA;MAPQ=60;MATEID=856038_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_76758501_76783501_60C;SPAN=1900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:15 GQ:6 PL:[66.0, 6.0, 0.0] SR:23 DR:0 LR:-66.02 LO:66.02);ALT=T[chr2:76775453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	76933615	+	chr2	76954376	+	.	12	0	856676_1	19.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=856676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:76933615(+)-2:76954376(-)__2_76930001_76955001D;SPAN=20761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:76 GQ:19.1 PL:[19.1, 0.0, 164.3] SR:0 DR:12 LR:-19.02 LO:25.83);ALT=C[chr2:76954376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	76954526	+	chr2	76933724	+	.	19	0	856677_1	46.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=856677_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:76933724(-)-2:76954526(+)__2_76930001_76955001D;SPAN=20802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:60 GQ:46.4 PL:[46.4, 0.0, 99.2] SR:0 DR:19 LR:-46.46 LO:47.51);ALT=]chr2:76954526]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	77007965	-	chr2	77023914	+	.	9	0	857025_1	11.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=857025_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:77007965(-)-2:77023914(-)__2_77003501_77028501D;SPAN=15949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=[chr2:77023914[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	84652727	+	chr2	84658631	+	.	0	17	872894_1	32.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=872894_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_84647501_84672501_313C;SPAN=5904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:88 GQ:32.3 PL:[32.3, 0.0, 180.8] SR:17 DR:0 LR:-32.28 LO:38.24);ALT=C[chr2:84658631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84668585	+	chr2	84670407	+	.	0	24	872927_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=872927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_84647501_84672501_132C;SPAN=1822;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:99 GQ:52.4 PL:[52.4, 0.0, 187.7] SR:24 DR:0 LR:-52.4 LO:56.69);ALT=T[chr2:84670407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84670527	+	chr2	84676772	+	.	0	57	873021_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=873021_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_84672001_84697001_349C;SPAN=6245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:53 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:57 DR:0 LR:-168.3 LO:168.3);ALT=G[chr2:84676772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84670575	+	chr2	84686302	+	.	71	0	873023_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=873023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:84670575(+)-2:84686302(-)__2_84672001_84697001D;SPAN=15727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:40 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=A[chr2:84686302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	84676876	+	chr2	84686297	+	.	35	10	873035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=873035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_84672001_84697001_74C;SPAN=9421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:67 GQ:61.1 PL:[100.7, 0.0, 61.1] SR:10 DR:35 LR:-101.2 LO:101.2);ALT=A[chr2:84686297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85329762	-	chr3	14239532	+	.	11	0	1288948_1	29.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=1288948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85329762(-)-3:14239532(-)__3_14234501_14259501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=[chr3:14239532[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	85337505	-	chr9	110537537	+	.	3	11	4384710_1	31.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCCTCTTTCTTTTCAATTACTGTGTCTCTTGTCT;MAPQ=60;MATEID=4384710_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_110519501_110544501_168C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:32 GQ:31.1 PL:[31.1, 0.0, 44.3] SR:11 DR:3 LR:-30.94 LO:31.12);ALT=[chr9:110537537[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	85549867	+	chr2	85553631	+	CTGGTCCAAACGTTGGTAGTCACTGGCCTTTGGCCGCCGGGTGACTTTAGATCTTTTTCCTTCCAGGACAAAAGCAATGAT	0	14	875524_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTGGTCCAAACGTTGGTAGTCACTGGCCTTTGGCCGCCGGGTGACTTTAGATCTTTTTCCTTCCAGGACAAAAGCAATGAT;MAPQ=60;MATEID=875524_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_85529501_85554501_19C;SPAN=3764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:64 GQ:29 PL:[29.0, 0.0, 124.7] SR:14 DR:0 LR:-28.88 LO:32.35);ALT=T[chr2:85553631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85549867	+	chr2	85552038	+	.	2	8	875523_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTT;MAPQ=60;MATEID=875523_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_2_85529501_85554501_19C;SPAN=2171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:8 DR:2 LR:-11.02 LO:18.56);ALT=T[chr2:85552038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85622750	+	chr2	85625142	+	.	3	36	875857_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=875857_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85603001_85628001_16C;SPAN=2392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:121 GQ:92.9 PL:[92.9, 0.0, 198.5] SR:36 DR:3 LR:-92.66 LO:94.86);ALT=C[chr2:85625142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85625908	+	chr2	85628288	+	GATCATCTCAGCAGGCTCCTCCCCATCAGTGACAATCTCCACCTGGGCCTTGCCCTGTCGCTCACTGTCCCGGATGGCCAGGGCCAGGTCCCTCGCCTTGTTGCGTTCCAGGATGTTGGACTTTCCACCACACCAGGCGAAGATGTT	0	32	875672_1	95.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GATCATCTCAGCAGGCTCCTCCCCATCAGTGACAATCTCCACCTGGGCCTTGCCCTGTCGCTCACTGTCCCGGATGGCCAGGGCCAGGTCCCTCGCCTTGTTGCGTTCCAGGATGTTGGACTTTCCACCACACCAGGCGAAGATGTT;MAPQ=60;MATEID=875672_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_85627501_85652501_87C;SPAN=2380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:39 GQ:0.6 PL:[95.7, 0.6, 0.0] SR:32 DR:0 LR:-101.1 LO:101.1);ALT=G[chr2:85628288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85626411	+	chr2	85628288	+	.	25	9	875673_1	91.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=875673_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_2_85627501_85652501_87C;SPAN=1877;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:39 GQ:2.6 PL:[91.7, 0.0, 2.6] SR:9 DR:25 LR:-96.83 LO:96.83);ALT=G[chr2:85628288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85629118	+	chr2	85637404	+	.	147	0	875683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=875683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85629118(+)-2:85637404(-)__2_85627501_85652501D;SPAN=8286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:85 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:0 DR:147 LR:-435.7 LO:435.7);ALT=A[chr2:85637404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85629142	+	chr2	85641105	+	.	42	0	875684_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=875684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85629142(+)-2:85641105(-)__2_85627501_85652501D;SPAN=11963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:97 GQ:99 PL:[112.4, 0.0, 122.3] SR:0 DR:42 LR:-112.4 LO:112.4);ALT=A[chr2:85641105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85766501	+	chr2	85768202	+	.	0	10	876007_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=876007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85750001_85775001_192C;SPAN=1701;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:10 DR:0 LR:-12.96 LO:20.79);ALT=G[chr2:85768202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85804773	+	chr2	85806131	+	.	106	5	876458_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=876458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85799001_85824001_256C;SPAN=1358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:143 DP:268 GQ:99 PL:[399.5, 0.0, 250.9] SR:5 DR:106 LR:-401.2 LO:401.2);ALT=G[chr2:85806131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85804826	+	chr2	85808698	+	.	94	0	876460_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=876460_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:85804826(+)-2:85808698(-)__2_85799001_85824001D;SPAN=3872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:161 GQ:99 PL:[266.9, 0.0, 121.7] SR:0 DR:94 LR:-269.5 LO:269.5);ALT=C[chr2:85808698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85806290	+	chr2	85808699	+	.	11	139	876464_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=876464_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85799001_85824001_108C;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:149 DP:266 GQ:99 PL:[419.9, 0.0, 225.1] SR:139 DR:11 LR:-422.9 LO:422.9);ALT=A[chr2:85808699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85822972	+	chr2	85824225	+	CTGCATTCTGCCCTGGCTAAGCA	2	47	876194_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGCATTCTGCCCTGGCTAAGCA;MAPQ=60;MATEID=876194_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85823501_85848501_315C;SPAN=1253;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:47 DR:2 LR:-160.5 LO:160.5);ALT=G[chr2:85824225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85843586	+	chr2	85846341	+	.	5	8	876257_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=876257_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_85823501_85848501_334C;SPAN=2755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:8 DR:5 LR:-7.543 LO:19.68);ALT=G[chr2:85846341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	85923179	+	chr2	85924626	+	.	0	5	876760_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=876760_2;MATENM=1;NM=0;NUMPARTS=4;SCTG=c_2_85921501_85946501_312C;SPAN=1447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:78 GQ:4.5 PL:[0.0, 4.5, 198.0] SR:5 DR:0 LR:4.627 LO:8.689);ALT=G[chr2:85924626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86333452	+	chr19	57686685	+	.	8	0	6876350_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6876350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:86333452(+)-19:57686685(-)__19_57673001_57698001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.59 LO:17.19);ALT=T[chr19:57686685[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	86406758	+	chr2	86422472	+	.	10	0	878100_1	23.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=878100_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:86406758(+)-2:86422472(-)__2_86411501_86436501D;SPAN=15714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:36 GQ:23.3 PL:[23.3, 0.0, 62.9] SR:0 DR:10 LR:-23.26 LO:24.32);ALT=A[chr2:86422472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86734718	+	chr2	86737480	+	.	3	2	879047_1	0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=879047_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_86730001_86755001_415C;SPAN=2762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:86 GQ:6.6 PL:[0.0, 6.6, 221.1] SR:2 DR:3 LR:6.795 LO:8.471);ALT=T[chr2:86737480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86737603	+	chr2	86756341	+	.	0	10	879059_1	20.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=879059_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_86730001_86755001_19C;SPAN=18738;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:10 DR:0 LR:-20.28 LO:22.97);ALT=C[chr2:86756341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86754365	+	chr2	86756341	+	.	0	7	879225_1	10.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=879225_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_86754501_86779501_75C;SPAN=1976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:7 DR:0 LR:-10.37 LO:14.87);ALT=C[chr2:86756341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	86756521	+	chr2	86790425	+	CCTTATTTGCCTGTCAACAACTCTCATTTCCTTTCTTATCTTCAATGACCACTCATTG	32	20	879231_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=CCTTATTTGCCTGTCAACAACTCTCATTTCCTTTCTTATCTTCAATGACCACTCATTG;MAPQ=60;MATEID=879231_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_86754501_86779501_183C;SPAN=33904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:20 DR:32 LR:-118.8 LO:118.8);ALT=C[chr2:86790425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	88333813	+	chr2	88355145	+	CATAATGCAAAATCCTTTGTTATTTGAACTGTAACACTACTCCACAGACATCTTTTATAAAAGGTATCTGTAAACAAAGTTCAGTCTTTGTTCATTCAATGTGGTAT	2	13	884968_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CATAATGCAAAATCCTTTGTTATTTGAACTGTAACACTACTCCACAGACATCTTTTATAAAAGGTATCTGTAAACAAAGTTCAGTCTTTGTTCATTCAATGTGGTAT;MAPQ=60;MATEID=884968_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_88322501_88347501_94C;SPAN=21332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:40 GQ:38.6 PL:[38.6, 0.0, 58.4] SR:13 DR:2 LR:-38.68 LO:38.9);ALT=T[chr2:88355145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	88336572	+	chr2	88355145	+	.	0	9	885080_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=885080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_88347001_88372001_240C;SPAN=18573;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:23 GQ:23.6 PL:[23.6, 0.0, 30.2] SR:9 DR:0 LR:-23.48 LO:23.56);ALT=T[chr2:88355145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	88689149	-	chr6	107399772	+	.	7	31	2974369_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=GGCTCACGCCTGTAATCCCAGCACTTTGGGAGGCTGAGG;MAPQ=34;MATEID=2974369_2;MATENM=1;NM=8;NUMPARTS=2;SCTG=c_6_107383501_107408501_144C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:60 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:31 DR:7 LR:-107.5 LO:107.5);ALT=[chr6:107399772[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	89029246	+	chr2	89032283	+	.	82	30	887260_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATATTAAAACTAAG;MAPQ=60;MATEID=887260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_89008501_89033501_104C;SPAN=3037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:99 DP:164 GQ:99 PL:[282.5, 0.0, 114.2] SR:30 DR:82 LR:-286.2 LO:286.2);ALT=G[chr2:89032283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	89835562	+	chr2	89830441	+	.	8	0	892315_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=892315_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:89830441(-)-2:89835562(+)__2_89817001_89842001D;SPAN=5121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:153 GQ:14.8 PL:[0.0, 14.8, 399.3] SR:0 DR:8 LR:15.04 LO:13.18);ALT=]chr2:89835562]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	89831994	+	chr2	89833326	+	.	0	35	892332_1	60.0	.	EVDNC=ASSMB;HOMSEQ=TGATGATTCCATTCGA;MAPQ=60;MATEID=892332_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_89817001_89842001_231C;SPAN=1332;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:203 GQ:60.7 PL:[60.7, 0.0, 430.4] SR:35 DR:0 LR:-60.54 LO:76.8);ALT=A[chr2:89833326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	89850662	+	chr2	89853637	+	.	44	25	893566_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATTTGAGTCCATTCCATCCCACTCCATT;MAPQ=60;MATEID=893566_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_89841501_89866501_311C;SPAN=2975;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:138 GQ:99 PL:[177.2, 0.0, 157.4] SR:25 DR:44 LR:-177.2 LO:177.2);ALT=T[chr2:89853637[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	89870200	-	chr2	89877008	+	.	12	0	891135_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=891135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:89870200(-)-2:89877008(-)__2_89866001_89891001D;SPAN=6808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:235 GQ:23.8 PL:[0.0, 23.8, 617.2] SR:0 DR:12 LR:24.06 LO:19.64);ALT=[chr2:89877008[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	95775786	+	chr2	95780811	+	.	2	10	899613_1	19.0	.	DISC_MAPQ=30;EVDNC=ASDIS;MAPQ=60;MATEID=899613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_95770501_95795501_207C;SPAN=5025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:10 DR:2 LR:-19.29 LO:25.9);ALT=A[chr2:95780811[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	95780949	+	chr2	95787477	+	ATTGCCGAGAACACTCTTCCATGCCAAAATGGAAGCTGCTGGTAAGGTGTTTAGGGAACACTGCCTCCCCAATAAATG	19	41	899636_1	99.0	.	DISC_MAPQ=49;EVDNC=TSI_G;HOMSEQ=ACCTGC;INSERTION=ATTGCCGAGAACACTCTTCCATGCCAAAATGGAAGCTGCTGGTAAGGTGTTTAGGGAACACTGCCTCCCCAATAAATG;MAPQ=60;MATEID=899636_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_95770501_95795501_214C;SPAN=6528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:83 GQ:60.2 PL:[139.4, 0.0, 60.2] SR:41 DR:19 LR:-140.9 LO:140.9);ALT=C[chr2:95787477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	95783694	+	chr2	95787477	+	.	8	15	899643_1	44.0	.	DISC_MAPQ=33;EVDNC=TSI_L;HOMSEQ=ACCTGC;MAPQ=60;MATEID=899643_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_95770501_95795501_214C;SPAN=3783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:78 GQ:44.9 PL:[44.9, 0.0, 143.9] SR:15 DR:8 LR:-44.89 LO:47.81);ALT=C[chr2:95787477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	96068621	+	chr2	96071298	+	.	10	7	900998_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=900998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_96064501_96089501_211C;SPAN=2677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:80 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:7 DR:10 LR:-24.54 LO:30.82);ALT=G[chr2:96071298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	96861289	+	chr2	96873883	+	.	9	3	903759_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=903759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_96873001_96898001_254C;SPAN=12594;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:3 DR:9 LR:-11.02 LO:18.56);ALT=T[chr2:96873883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	96969068	+	chr2	96970442	+	.	2	11	903672_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=903672_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_96946501_96971501_309C;SPAN=1374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:11 DR:2 LR:-18.21 LO:25.61);ALT=C[chr2:96970442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	97202601	+	chr2	97213137	+	.	9	0	904358_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=904358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97202601(+)-2:97213137(-)__2_97191501_97216501D;SPAN=10536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:0 DR:9 LR:-9.119 LO:18.15);ALT=C[chr2:97213137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	97519385	+	chr2	97523633	+	.	15	0	905374_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=905374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97519385(+)-2:97523633(-)__2_97510001_97535001D;SPAN=4248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:86 GQ:26.3 PL:[26.3, 0.0, 181.4] SR:0 DR:15 LR:-26.22 LO:33.0);ALT=G[chr2:97523633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	97520205	+	chr2	97523623	+	.	9	0	905375_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=905375_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97520205(+)-2:97523623(-)__2_97510001_97535001D;SPAN=3418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:0 DR:9 LR:-8.577 LO:18.05);ALT=A[chr2:97523623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	97873675	+	chr2	97875508	+	.	30	0	906475_1	92.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=906475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:97873675(+)-2:97875508(-)__2_97853001_97878001D;SPAN=1833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:32 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:30 LR:-92.42 LO:92.42);ALT=C[chr2:97875508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	98262654	+	chr2	98264459	+	GGTGTTCCCACTGATGAAGAGCAGGCGACTGGGTTGGAGAGGGAGATCATGCTGGCTGCAAAGAAGGGACTGGACCCATACAATGTACTGGCCCCAAAGGGAGCTTCAGGCACCAGGGAAGACCCTAATTTAGTCCCCTCCATCTCCAACAAGAGAATAGTAGGCTGCATCT	0	202	908428_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=GGTGTTCCCACTGATGAAGAGCAGGCGACTGGGTTGGAGAGGGAGATCATGCTGGCTGCAAAGAAGGGACTGGACCCATACAATGTACTGGCCCCAAAGGGAGCTTCAGGCACCAGGGAAGACCCTAATTTAGTCCCCTCCATCTCCAACAAGAGAATAGTAGGCTGCATCT;MAPQ=60;MATEID=908428_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_98245001_98270001_178C;SPAN=1805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:202 DP:170 GQ:54.4 PL:[597.4, 54.4, 0.0] SR:202 DR:0 LR:-597.4 LO:597.4);ALT=T[chr2:98264459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	98278409	+	chr2	98280305	+	.	5	4	908043_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=908043_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=CC;SCTG=c_2_98269501_98294501_323C;SPAN=1896;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:55 GQ:8.3 PL:[8.3, 0.0, 123.8] SR:4 DR:5 LR:-8.206 LO:14.35);ALT=C[chr2:98280305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99217257	+	chr2	99224769	+	ACTGATCTTTTACACTCAAAAAATGCGTACTTCAAAGAGTTGCAGTATCCTTCCTTCAAACACTGCCGAGGTGATTTTCCTT	7	35	910566_1	95.0	.	DISC_MAPQ=37;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=ACTGATCTTTTACACTCAAAAAATGCGTACTTCAAAGAGTTGCAGTATCCTTCCTTCAAACACTGCCGAGGTGATTTTCCTT;MAPQ=60;MATEID=910566_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_99200501_99225501_182C;SPAN=7512;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:85 GQ:95.9 PL:[95.9, 0.0, 109.1] SR:35 DR:7 LR:-95.81 LO:95.87);ALT=C[chr2:99224769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99220687	+	chr2	99224865	+	.	16	0	910573_1	35.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=910573_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:99220687(+)-2:99224865(-)__2_99200501_99225501D;SPAN=4178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:66 GQ:35 PL:[35.0, 0.0, 124.1] SR:0 DR:16 LR:-34.94 LO:37.79);ALT=T[chr2:99224865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99343031	+	chr2	99347510	+	.	32	3	910762_1	97.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=910762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_99323001_99348001_166C;SPAN=4479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:55 GQ:34.7 PL:[97.4, 0.0, 34.7] SR:3 DR:32 LR:-98.87 LO:98.87);ALT=C[chr2:99347510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99790520	+	chr2	99797390	+	.	13	0	911929_1	24.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=911929_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:99790520(+)-2:99797390(-)__2_99788501_99813501D;SPAN=6870;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:67 GQ:24.8 PL:[24.8, 0.0, 137.0] SR:0 DR:13 LR:-24.76 LO:29.27);ALT=T[chr2:99797390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99868361	+	chr6	119043030	+	.	12	24	3001826_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGAGTCTCACTCTGTCGCCCAGGCTGGAGTGCAGTGGC;MAPQ=60;MATEID=3001826_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_119021001_119046001_263C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:50 GQ:22.7 PL:[98.6, 0.0, 22.7] SR:24 DR:12 LR:-101.4 LO:101.4);ALT=C[chr6:119043030[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	99949723	+	chr2	99952723	+	.	13	0	912595_1	21.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=912595_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:99949723(+)-2:99952723(-)__2_99935501_99960501D;SPAN=3000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:78 GQ:21.8 PL:[21.8, 0.0, 167.0] SR:0 DR:13 LR:-21.78 LO:28.31);ALT=A[chr2:99952723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	99954052	+	chr2	99976697	+	.	0	36	912604_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=912604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_99935501_99960501_31C;SPAN=22645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:57 GQ:34.1 PL:[103.4, 0.0, 34.1] SR:36 DR:0 LR:-105.3 LO:105.3);ALT=G[chr2:99976697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	100512454	+	chr12	7108135	-	.	13	13	913643_1	75.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GGTTCAAGCAATTCTCCTGCCTCAGCCTCC;MAPQ=16;MATEID=913643_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_100499001_100524001_337C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:38 GQ:16.1 PL:[75.5, 0.0, 16.1] SR:13 DR:13 LR:-77.64 LO:77.64);ALT=C]chr12:7108135];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	100754401	+	chr2	100758946	+	.	25	7	914294_1	67.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=914294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_100744001_100769001_58C;SPAN=4545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:93 GQ:67.4 PL:[67.4, 0.0, 156.5] SR:7 DR:25 LR:-67.23 LO:69.27);ALT=T[chr2:100758946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	101179561	+	chr3	101431300	+	.	25	0	1558979_1	66.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1558979_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:101179561(+)-3:101431300(-)__3_101430001_101455001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:61 GQ:66.2 PL:[66.2, 0.0, 79.4] SR:0 DR:25 LR:-66.0 LO:66.1);ALT=G[chr3:101431300[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	101941207	+	chr14	73761581	-	.	0	32	5796825_1	80.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GCACTTT;MAPQ=60;MATEID=5796825_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCTTCT;SCTG=c_14_73745001_73770001_26C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:37 GQ:7.2 PL:[80.6, 7.2, 0.0] SR:32 DR:0 LR:-80.85 LO:80.85);ALT=C]chr14:73761581];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	104694509	+	chr7	135542434	+	.	6	31	924199_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGTGGAGGGTGAGCAAGATGA;MAPQ=60;MATEID=924199_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_104688501_104713501_287C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:25 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:31 DR:6 LR:-102.3 LO:102.3);ALT=A[chr7:135542434[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	105654648	+	chr2	105665626	+	.	13	0	926367_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=926367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:105654648(+)-2:105665626(-)__2_105644001_105669001D;SPAN=10978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:83 GQ:20.6 PL:[20.6, 0.0, 179.0] SR:0 DR:13 LR:-20.43 LO:27.93);ALT=C[chr2:105665626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	116974340	-	chr2	116981887	+	ACT	23	16	958731_1	95.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ACT;MAPQ=60;MATEID=958731_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_172C;SPAN=7547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:87 GQ:95.3 PL:[95.3, 0.0, 115.1] SR:16 DR:23 LR:-95.27 LO:95.38);ALT=[chr2:116981887[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	116974634	+	chr2	116978304	+	.	24	22	958733_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=958733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_95C;SPAN=3670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:79 GQ:84.2 PL:[107.3, 0.0, 84.2] SR:22 DR:24 LR:-107.5 LO:107.5);ALT=T[chr2:116978304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	116978299	+	chr2	116982310	-	.	27	17	958741_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATA;MAPQ=60;MATEID=958741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_116963001_116988001_61C;SPAN=4011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:79 GQ:84.2 PL:[107.3, 0.0, 84.2] SR:17 DR:27 LR:-107.5 LO:107.5);ALT=A]chr2:116982310];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	117853169	-	chr10	3139269	+	.	14	0	4495967_1	39.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=4495967_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:117853169(-)-10:3139269(-)__10_3136001_3161001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:6 GQ:3.6 PL:[39.6, 3.6, 0.0] SR:0 DR:14 LR:-39.61 LO:39.61);ALT=[chr10:3139269[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	117853389	+	chr10	3139011	-	.	18	0	4495968_1	52.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4495968_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:117853389(+)-10:3139011(+)__10_3136001_3161001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:15 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=C]chr10:3139011];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	118572439	+	chr2	118575019	+	.	36	34	962222_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=962222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_118555501_118580501_305C;SPAN=2580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:89 GQ:18.8 PL:[197.0, 0.0, 18.8] SR:34 DR:36 LR:-205.7 LO:205.7);ALT=G[chr2:118575019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	119653329	+	chr2	119659369	+	.	63	48	964901_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CGGCACTGGCTT;MAPQ=60;MATEID=964901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_119633501_119658501_153C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:28 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:48 DR:63 LR:-274.0 LO:274.0);ALT=T[chr2:119659369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	119711274	-	chr2	119712441	+	.	9	0	964610_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=964610_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:119711274(-)-2:119712441(-)__2_119707001_119732001D;SPAN=1167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:93 GQ:4.7 PL:[4.7, 0.0, 219.2] SR:0 DR:9 LR:-4.513 LO:17.32);ALT=[chr2:119712441[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	120124668	+	chr2	120125759	+	.	63	0	965746_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=965746_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:120124668(+)-2:120125759(-)__2_120123501_120148501D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:97 GQ:53 PL:[181.7, 0.0, 53.0] SR:0 DR:63 LR:-185.5 LO:185.5);ALT=T[chr2:120125759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120124670	+	chr2	120128313	+	.	29	0	965747_1	62.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=965747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:120124670(+)-2:120128313(-)__2_120123501_120148501D;SPAN=3643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:124 GQ:62.3 PL:[62.3, 0.0, 237.2] SR:0 DR:29 LR:-62.13 LO:67.97);ALT=C[chr2:120128313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120124677	+	chr2	120129818	+	.	15	0	965748_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=965748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:120124677(+)-2:120129818(-)__2_120123501_120148501D;SPAN=5141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:121 GQ:17 PL:[17.0, 0.0, 274.4] SR:0 DR:15 LR:-16.73 LO:30.57);ALT=C[chr2:120129818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120125881	+	chr2	120128314	+	.	0	213	965754_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=965754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_120123501_120148501_16C;SPAN=2433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:213 DP:158 GQ:57.4 PL:[630.4, 57.4, 0.0] SR:213 DR:0 LR:-630.5 LO:630.5);ALT=G[chr2:120128314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	120128379	+	chr2	120129819	+	.	7	219	965759_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=965759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_120123501_120148501_15C;SPAN=1440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:225 DP:144 GQ:60.7 PL:[666.7, 60.7, 0.0] SR:219 DR:7 LR:-666.8 LO:666.8);ALT=G[chr2:120129819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	102085249	+	chr2	120149146	+	GCACCTCAGCCTCCTGACCAGCTGGGATTACAGACATTCACCACAGAGCCTGGCTAATT	2	68	2117706_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;INSERTION=GCACCTCAGCCTCCTGACCAGCTGGGATTACAGACATTCACCACAGAGCCTGGCTAATT;MAPQ=60;MATEID=2117706_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_4_102067001_102092001_231C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:56 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:68 DR:2 LR:-208.0 LO:208.0);ALT=]chr4:102085249]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	120418488	+	chr2	120417080	+	GGC	37	72	966609_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GGC;MAPQ=60;MATEID=966609_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_2_120417501_120442501_334C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:25 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:72 DR:37 LR:-260.8 LO:260.8);ALT=]chr2:120418488]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	120417200	+	chr2	120418496	+	.	30	49	966610_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCC;MAPQ=60;MATEID=966610_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_120417501_120442501_249C;SPAN=1296;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:22 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:49 DR:30 LR:-194.7 LO:194.7);ALT=C[chr2:120418496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	121010556	+	chr2	121036193	+	.	20	8	968319_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=968319_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_121030001_121055001_104C;SPAN=25637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:58 GQ:56.9 PL:[56.9, 0.0, 83.3] SR:8 DR:20 LR:-56.91 LO:57.19);ALT=G[chr2:121036193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	121036354	+	chr2	121043448	+	.	7	9	968338_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=968338_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_121030001_121055001_232C;SPAN=7094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:9 DR:7 LR:-12.74 LO:22.52);ALT=G[chr2:121043448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	121361006	+	chr2	121362068	-	.	9	0	968954_1	7.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=968954_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:121361006(+)-2:121362068(+)__2_121348501_121373501D;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:82 GQ:7.7 PL:[7.7, 0.0, 189.2] SR:0 DR:9 LR:-7.493 LO:17.84);ALT=T]chr2:121362068];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	125766561	+	chr2	125768248	+	.	20	26	979655_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=979655_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_125758501_125783501_140C;SPAN=1687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:94 GQ:99 PL:[106.7, 0.0, 119.9] SR:26 DR:20 LR:-106.6 LO:106.6);ALT=C[chr2:125768248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	125768401	+	chr2	125766562	+	TCTATACTCACTACTACACTAT	0	30	979657_1	70.0	.	EVDNC=ASSMB;INSERTION=TCTATACTCACTACTACACTAT;MAPQ=60;MATEID=979657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_125758501_125783501_280C;SPAN=1839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:105 GQ:70.7 PL:[70.7, 0.0, 182.9] SR:30 DR:0 LR:-70.58 LO:73.39);ALT=]chr2:125768401]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	126443251	+	chr2	126451832	+	.	95	53	981173_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAAC;MAPQ=60;MATEID=981173_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_126444501_126469501_206C;SPAN=8581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:13 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:53 DR:95 LR:-373.0 LO:373.0);ALT=C[chr2:126451832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	127413860	+	chr2	127451435	+	.	16	0	983307_1	39.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=983307_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:127413860(+)-2:127451435(-)__2_127449001_127474001D;SPAN=37575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:50 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.27 LO:40.1);ALT=C[chr2:127451435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	127674758	+	chr2	127677273	+	.	85	53	983779_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=983779_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_127669501_127694501_17C;SPAN=2515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:27 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:53 DR:85 LR:-343.3 LO:343.3);ALT=C[chr2:127677273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	128528625	+	chr2	128568654	+	.	33	0	986631_1	95.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=986631_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:128528625(+)-2:128568654(-)__2_128527001_128552001D;SPAN=40029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:33 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:0 DR:33 LR:-95.72 LO:95.72);ALT=C[chr2:128568654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	128839986	+	chr12	22808468	+	.	24	0	987895_1	75.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=987895_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:128839986(+)-12:22808468(-)__2_128821001_128846001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:28 GQ:4.2 PL:[75.9, 4.2, 0.0] SR:0 DR:24 LR:-77.12 LO:77.12);ALT=T[chr12:22808468[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	129546068	-	chr2	129550109	+	.	9	1	989362_1	0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TGTGTGC;MAPQ=60;MATEID=989362_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_129531501_129556501_65C;SPAN=4041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:125 GQ:0.6 PL:[0.0, 0.6, 303.6] SR:1 DR:9 LR:0.8556 LO:18.37);ALT=[chr2:129550109[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	138722133	+	chr2	138724663	+	.	9	0	1014275_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1014275_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:138722133(+)-2:138724663(-)__2_138719001_138744001D;SPAN=2530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:91 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.055 LO:17.41);ALT=C[chr2:138724663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	139046347	+	chr17	1303411	+	.	35	0	6282323_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6282323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:139046347(+)-17:1303411(-)__17_1298501_1323501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:56 GQ:34.4 PL:[100.4, 0.0, 34.4] SR:0 DR:35 LR:-102.1 LO:102.1);ALT=T[chr17:1303411[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	153512932	+	chr2	153514401	+	.	9	0	1047145_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1047145_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:153512932(+)-2:153514401(-)__2_153492501_153517501D;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:0 DR:9 LR:-9.661 LO:18.26);ALT=A[chr2:153514401[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	153529558	+	chr2	153532919	+	TTTCTTTCAATAATTCTTTAAAAGCTTGCTTTGCCTCTTCCTTTGTATTCCAAGTGTATGTTTTCTTTGCTGGTTGGCTCTCCTCCTCTTCTTTTTTGGGAGTAAAA	0	21	1047210_1	49.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTTCTTTCAATAATTCTTTAAAAGCTTGCTTTGCCTCTTCCTTTGTATTCCAAGTGTATGTTTTCTTTGCTGGTTGGCTCTCCTCCTCTTCTTTTTTGGGAGTAAAA;MAPQ=60;MATEID=1047210_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_153517001_153542001_15C;SPAN=3361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:75 GQ:49.1 PL:[49.1, 0.0, 131.6] SR:21 DR:0 LR:-49.0 LO:51.15);ALT=T[chr2:153532919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	153551136	+	chr2	153572509	+	.	0	47	1047461_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1047461_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_153566001_153591001_129C;SPAN=21373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:39 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:47 DR:0 LR:-138.6 LO:138.6);ALT=T[chr2:153572509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	153551182	+	chr2	153573869	+	.	20	0	1047462_1	56.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1047462_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:153551182(+)-2:153573869(-)__2_153566001_153591001D;SPAN=22687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:36 GQ:29.9 PL:[56.3, 0.0, 29.9] SR:0 DR:20 LR:-56.66 LO:56.66);ALT=A[chr2:153573869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	153572641	+	chr2	153573870	+	.	34	6	1047485_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1047485_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_153566001_153591001_334C;SPAN=1229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:75 GQ:72.2 PL:[108.5, 0.0, 72.2] SR:6 DR:34 LR:-108.8 LO:108.8);ALT=C[chr2:153573870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	155006887	-	chr2	167547093	+	A	21	64	1079412_1	99.0	.	DISC_MAPQ=21;EVDNC=ASDIS;INSERTION=A;MAPQ=47;MATEID=1079412_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_167531001_167556001_372C;SPAN=12540206;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:24 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:64 DR:21 LR:-211.3 LO:211.3);ALT=[chr2:167547093[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	155007024	+	chr2	167545932	-	.	36	0	1079414_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=1079414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:155007024(+)-2:167545932(+)__2_167531001_167556001D;SPAN=12538908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:10 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=T]chr2:167545932];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	156126148	-	chr18	43666350	+	GCCACGACTCAAAAGTTGTTGAGTGGCAGCATCGAGGTCAGAACCGAACTGGGCAAAAGCAGCAACCTCACGATACTGAGCCAATTCCAGCTTCATGGTACCTGC	0	21	6609427_1	59.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TACCTGC;INSERTION=GCCACGACTCAAAAGTTGTTGAGTGGCAGCATCGAGGTCAGAACCGAACTGGGCAAAAGCAGCAACCTCACGATACTGAGCCAATTCCAGCTTCATGGTACCTGC;MAPQ=57;MATEID=6609427_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_18_43659001_43684001_85C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:37 GQ:29.6 PL:[59.3, 0.0, 29.6] SR:21 DR:0 LR:-59.79 LO:59.79);ALT=[chr18:43666350[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	164520323	+	chr2	203199395	-	.	19	16	1163927_1	89.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=GCCTCCCGGGTTCAAGCAATTCTCCTGCCTCAGCATCCTGAG;MAPQ=42;MATEID=1163927_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_2_203178501_203203501_124C;SPAN=38679072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:22 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:16 DR:19 LR:-89.12 LO:89.12);ALT=C]chr2:203199395];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	165430267	-	chr8	109228638	+	.	11	0	1074318_1	18.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1074318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:165430267(-)-8:109228638(-)__2_165424001_165449001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:0 DR:11 LR:-18.7 LO:24.04);ALT=[chr8:109228638[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	166888737	+	chr18	47205588	-	.	6	5	1077604_1	1.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACACACACACACACACACACACACA;MAPQ=60;MATEID=1077604_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=ACACACACACACACACACACACAC;SCTG=c_2_166869501_166894501_320C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:1 PL:[1.0, 0.0, 39.6] SR:5 DR:6 LR:-0.2054 LO:4.362);ALT=A]chr18:47205588];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	167545960	+	chr2	167547086	+	.	31	0	1079442_1	89.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=1079442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:167545960(+)-2:167547086(-)__2_167531001_167556001D;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:16 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=T[chr2:167547086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170105133	+	chr2	170111163	+	.	51	21	1085145_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAACAGCAATGTTGA;MAPQ=60;MATEID=1085145_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_170103501_170128501_12C;SPAN=6030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:55 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:21 DR:51 LR:-171.6 LO:171.6);ALT=A[chr2:170111163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170428682	+	chr2	170430179	+	.	0	7	1085979_1	2.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1085979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_170422001_170447001_99C;SPAN=1497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:76 GQ:2.6 PL:[2.6, 0.0, 180.8] SR:7 DR:0 LR:-2.517 LO:13.31);ALT=C[chr2:170430179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170441041	+	chr2	170460533	+	.	30	0	1086009_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1086009_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170441041(+)-2:170460533(-)__2_170422001_170447001D;SPAN=19492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:49 GQ:32.9 PL:[85.7, 0.0, 32.9] SR:0 DR:30 LR:-87.03 LO:87.03);ALT=T[chr2:170460533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170441407	+	chr2	170460533	+	.	14	0	1086012_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1086012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170441407(+)-2:170460533(-)__2_170422001_170447001D;SPAN=19126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:35 GQ:36.8 PL:[36.8, 0.0, 46.7] SR:0 DR:14 LR:-36.73 LO:36.82);ALT=G[chr2:170460533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170460773	+	chr2	170462547	+	.	0	16	1085899_1	31.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=45;MATEID=1085899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_170446501_170471501_268C;SPAN=1774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:80 GQ:31.1 PL:[31.1, 0.0, 163.1] SR:16 DR:0 LR:-31.14 LO:36.26);ALT=T[chr2:170462547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170465268	+	chr2	170471094	+	AACAACGAAACCAACTCCTCATTTAGATG	4	16	1085919_1	49.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TGACTTCAGTGAAGGAAATGGACGAGGAGGGGAATCTATCTATGGAGGATTTTTTGAAG;INSERTION=AACAACGAAACCAACTCCTCATTTAGATG;MAPQ=2;MATEID=1085919_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_170446501_170471501_114C;SPAN=5826;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:63 GQ:49.1 PL:[49.1, 0.0, 101.9] SR:16 DR:4 LR:-48.95 LO:50.04);ALT=T[chr2:170471094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170488443	+	chr2	170489669	+	.	0	4	1085817_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1085817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_170471001_170496001_221C;SPAN=1226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:4 DR:0 LR:6.844 LO:6.647);ALT=G[chr2:170489669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170551172	+	chr2	170553868	+	.	9	0	1085618_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1085618_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170551172(+)-2:170553868(-)__2_170544501_170569501D;SPAN=2696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:75 GQ:9.5 PL:[9.5, 0.0, 171.2] SR:0 DR:9 LR:-9.39 LO:18.21);ALT=T[chr2:170553868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170641518	+	chr2	170643952	+	.	70	41	1086336_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=TCATTATTTTC;MAPQ=60;MATEID=1086336_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_170618001_170643001_86C;SPAN=2434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:31 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:41 DR:70 LR:-280.6 LO:280.6);ALT=C[chr2:170643952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170655507	+	chr2	170661981	+	.	36	0	1086235_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1086235_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170655507(+)-2:170661981(-)__2_170642501_170667501D;SPAN=6474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:79 GQ:94.1 PL:[97.4, 0.0, 94.1] SR:0 DR:36 LR:-97.44 LO:97.44);ALT=A[chr2:170661981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170678569	+	chr2	170680999	+	.	0	13	1086749_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1086749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_170667001_170692001_382C;SPAN=2430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:13 DR:0 LR:-19.34 LO:27.64);ALT=T[chr2:170680999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	170678609	+	chr2	170681332	+	.	12	0	1086751_1	20.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1086751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:170678609(+)-2:170681332(-)__2_170667001_170692001D;SPAN=2723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:0 DR:12 LR:-20.92 LO:26.38);ALT=A[chr2:170681332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	171608279	-	chr20	32699970	+	.	15	0	6984855_1	30.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6984855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:171608279(-)-20:32699970(-)__20_32683001_32708001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:72 GQ:30.2 PL:[30.2, 0.0, 142.4] SR:0 DR:15 LR:-30.01 LO:34.3);ALT=[chr20:32699970[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	171785897	+	chr2	171804852	+	.	10	0	1089319_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1089319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:171785897(+)-2:171804852(-)__2_171769501_171794501D;SPAN=18955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:40 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-22.17 LO:23.78);ALT=G[chr2:171804852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	171804940	+	chr2	171806049	+	.	0	10	1089224_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1089224_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_171794001_171819001_83C;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:79 GQ:11.6 PL:[11.6, 0.0, 179.9] SR:10 DR:0 LR:-11.61 LO:20.48);ALT=A[chr2:171806049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172379248	+	chr2	172398094	+	.	0	11	1091049_1	24.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1091049_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172382001_172407001_7C;SPAN=18846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:11 DR:0 LR:-24.12 LO:26.03);ALT=G[chr2:172398094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172725335	+	chr2	172749715	+	.	4	6	1092110_1	22.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1092110_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_2_172749501_172774501_69C;SPAN=24380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:38 GQ:22.7 PL:[22.7, 0.0, 68.9] SR:6 DR:4 LR:-22.72 LO:24.04);ALT=T[chr2:172749715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172725335	+	chr2	172750710	+	GTAGAAATATGTTTCTTAACTCATGAGGATCCCCTCGCTTAGTTGTCTG	23	7	1092111_1	80.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CACCT;INSERTION=GTAGAAATATGTTTCTTAACTCATGAGGATCCCCTCGCTTAGTTGTCTG;MAPQ=60;MATEID=1092111_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_2_172749501_172774501_69C;SPAN=25375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:46 GQ:30.5 PL:[80.0, 0.0, 30.5] SR:7 DR:23 LR:-81.11 LO:81.11);ALT=T[chr2:172750710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172779018	+	chr2	172782046	+	.	6	3	1092051_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1092051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172774001_172799001_2C;SPAN=3028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:3 DR:6 LR:2.902 LO:12.57);ALT=G[chr2:172782046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172779066	+	chr2	172803225	+	.	10	0	1092277_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1092277_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:172779066(+)-2:172803225(-)__2_172798501_172823501D;SPAN=24159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:36 GQ:23.3 PL:[23.3, 0.0, 62.9] SR:0 DR:10 LR:-23.26 LO:24.32);ALT=G[chr2:172803225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172779069	+	chr2	172809396	+	.	10	0	1092278_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1092278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:172779069(+)-2:172809396(-)__2_172798501_172823501D;SPAN=30327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:26 GQ:26 PL:[26.0, 0.0, 35.9] SR:0 DR:10 LR:-25.97 LO:26.07);ALT=T[chr2:172809396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172782151	+	chr2	172803226	+	.	3	15	1092280_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1092280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172798501_172823501_184C;SPAN=21075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:37 GQ:42.8 PL:[42.8, 0.0, 46.1] SR:15 DR:3 LR:-42.79 LO:42.8);ALT=G[chr2:172803226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172782152	+	chr2	172793489	+	.	3	4	1092063_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAGG;MAPQ=60;MATEID=1092063_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172774001_172799001_24C;SPAN=11337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:4 DR:3 LR:-3.059 LO:13.4);ALT=G[chr2:172793489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172803303	+	chr2	172809399	+	.	0	15	1092298_1	34.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1092298_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172798501_172823501_73C;SPAN=6096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:55 GQ:34.7 PL:[34.7, 0.0, 97.4] SR:15 DR:0 LR:-34.61 LO:36.33);ALT=A[chr2:172809399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172864947	+	chr2	172926231	+	.	13	0	1092454_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1092454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:172864947(+)-2:172926231(-)__2_172921001_172946001D;SPAN=61284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:42 GQ:31.7 PL:[31.7, 0.0, 68.0] SR:0 DR:13 LR:-31.53 LO:32.35);ALT=T[chr2:172926231[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172864954	+	chr2	172928435	+	.	8	0	1092455_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1092455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:172864954(+)-2:172928435(-)__2_172921001_172946001D;SPAN=63481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=G[chr2:172928435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	172926383	+	chr2	172928436	+	.	0	12	1092471_1	11.0	.	EVDNC=ASSMB;HOMSEQ=AAG;MAPQ=60;MATEID=1092471_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172921001_172946001_62C;SPAN=2053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:106 GQ:11 PL:[11.0, 0.0, 245.3] SR:12 DR:0 LR:-10.89 LO:23.95);ALT=G[chr2:172928436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	173004263	+	chr2	173007481	+	.	85	36	1092750_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GTAGAGATGGGGTTT;MAPQ=60;MATEID=1092750_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_172994501_173019501_230C;SPAN=3218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:25 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:36 DR:85 LR:-290.5 LO:290.5);ALT=T[chr2:173007481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41576288	+	chr2	173030023	+	.	10	0	5933266_1	23.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5933266_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:173030023(-)-15:41576288(+)__15_41552001_41577001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:34 GQ:23.9 PL:[23.9, 0.0, 56.9] SR:0 DR:10 LR:-23.8 LO:24.62);ALT=]chr15:41576288]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	173940730	+	chr2	173955723	+	.	9	5	1095311_1	24.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1095311_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_173925501_173950501_130C;SPAN=14993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:31 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:5 DR:9 LR:-24.61 LO:25.11);ALT=G[chr2:173955723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	175094189	+	chr2	175113178	+	.	58	0	1098190_1	99.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=1098190_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:175094189(+)-2:175113178(-)__2_175101501_175126501D;SPAN=18989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:31 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=A[chr2:175113178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42504992	+	chr2	175113176	+	.	61	0	7311591_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7311591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:175113176(-)-22:42504992(+)__22_42483001_42508001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:66 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:0 DR:61 LR:-194.7 LO:194.7);ALT=]chr22:42504992]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	175213903	+	chr2	175215387	+	.	0	5	1098284_1	0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=1098284_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_175199501_175224501_280C;SPAN=1484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:76 GQ:3.9 PL:[0.0, 3.9, 191.4] SR:5 DR:0 LR:4.085 LO:8.747);ALT=G[chr2:175215387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	175252507	+	chr2	175260277	+	.	13	9	1098520_1	40.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=48;MATEID=1098520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_175248501_175273501_140C;SPAN=7770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:83 GQ:40.4 PL:[40.4, 0.0, 159.2] SR:9 DR:13 LR:-40.23 LO:44.33);ALT=C[chr2:175260277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	175348648	-	chr2	175349684	+	.	14	0	1098830_1	23.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1098830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:175348648(-)-2:175349684(-)__2_175346501_175371501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:85 GQ:23.3 PL:[23.3, 0.0, 181.7] SR:0 DR:14 LR:-23.19 LO:30.41);ALT=[chr2:175349684[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	175446168	+	chr2	175462329	+	AGTGCAAACGTCGGGGGCGGCGGGGGTGCTGGAGGGGGAGGGACAGGCATCTTGGGCAGTTATGCGTTCAACAGTCTTGCTGATAAAT	0	20	1099108_1	46.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGTGCAAACGTCGGGGGCGGCGGGGGTGCTGGAGGGGGAGGGACAGGCATCTTGGGCAGTTATGCGTTCAACAGTCTTGCTGATAAAT;MAPQ=60;MATEID=1099108_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_175444501_175469501_221C;SPAN=16161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:72 GQ:46.7 PL:[46.7, 0.0, 125.9] SR:20 DR:0 LR:-46.51 LO:48.63);ALT=C[chr2:175462329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176043980	+	chr2	176046083	+	CTCCAGTCCTACTAGCCTCTGGTCGAGATAACACTGATGCAGAAATTGGTCTGTATGCAACTCTGGATCCAGCTCGGAT	13	217	1100780_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTCCAGTCCTACTAGCCTCTGGTCGAGATAACACTGATGCAGAAATTGGTCTGTATGCAACTCTGGATCCAGCTCGGAT;MAPQ=60;MATEID=1100780_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_176032501_176057501_37C;SPAN=2103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:224 DP:193 GQ:60.4 PL:[663.4, 60.4, 0.0] SR:217 DR:13 LR:-663.5 LO:663.5);ALT=T[chr2:176046083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176044031	+	chr2	176046382	+	.	87	0	1100781_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1100781_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:176044031(+)-2:176046382(-)__2_176032501_176057501D;SPAN=2351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:210 GQ:99 PL:[230.3, 0.0, 279.8] SR:0 DR:87 LR:-230.3 LO:230.6);ALT=T[chr2:176046382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176044907	+	chr2	176046083	+	.	4	99	1100785_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1100785_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_2_176032501_176057501_37C;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:103 DP:187 GQ:99 PL:[289.4, 0.0, 164.0] SR:99 DR:4 LR:-291.2 LO:291.2);ALT=C[chr2:176046083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176044956	+	chr2	176046382	+	.	97	0	1100786_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1100786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:176044956(+)-2:176046382(-)__2_176032501_176057501D;SPAN=1426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:201 GQ:99 PL:[266.0, 0.0, 219.8] SR:0 DR:97 LR:-265.9 LO:265.9);ALT=T[chr2:176046382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	176335115	+	chr2	176336296	-	.	2	28	1101594_1	50.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGTCC;MAPQ=60;MATEID=1101594_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_2_176326501_176351501_163C;SPAN=1181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:167 GQ:50.6 PL:[50.6, 0.0, 354.2] SR:28 DR:2 LR:-50.49 LO:63.73);ALT=C]chr2:176336296];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	177265645	+	chr2	177272041	+	.	97	76	1103493_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATT;MAPQ=60;MATEID=1103493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_177257501_177282501_173C;SPAN=6396;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:39 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:76 DR:97 LR:-412.6 LO:412.6);ALT=T[chr2:177272041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	177355934	-	chr2	177357086	+	.	8	0	1103684_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1103684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:177355934(-)-2:177357086(-)__2_177355501_177380501D;SPAN=1152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=[chr2:177357086[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	181880746	+	chr22	22250027	-	.	3	37	1114398_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GAATTG;MAPQ=60;MATEID=1114398_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_181863501_181888501_310C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:43 GQ:8.1 PL:[118.8, 8.1, 0.0] SR:37 DR:3 LR:-119.1 LO:119.1);ALT=C]chr22:22250027];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	182322579	+	chr2	182339686	+	CTCCTAGTGGGTGCGCCCACTGCCAACTGGCTCGCCAACGCTTCAGTGATCAATCCCGGGGCGATTTACAGATGCAGGATCGGAAAGAATCCCGGCCAGACGTGCGAACAGCTCCAGCTG	0	49	1115478_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=CTCCTAGTGGGTGCGCCCACTGCCAACTGGCTCGCCAACGCTTCAGTGATCAATCCCGGGGCGATTTACAGATGCAGGATCGGAAAGAATCCCGGCCAGACGTGCGAACAGCTCCAGCTG;MAPQ=60;MATEID=1115478_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_182304501_182329501_54C;SPAN=17107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:36 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:49 DR:0 LR:-145.2 LO:145.2);ALT=G[chr2:182339686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	182323046	+	chr2	182339686	+	.	22	25	1115479_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=1115479_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_182304501_182329501_54C;SPAN=16640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:60 GQ:23.3 PL:[122.3, 0.0, 23.3] SR:25 DR:22 LR:-126.2 LO:126.2);ALT=T[chr2:182339686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	182340015	+	chr2	182344862	+	ATTATGTGAAAAAATTTGGAGAAAATTTTGCATCATGTCAAGCTGGAATATCCAGTTTTTACACAA	9	16	1115328_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTATGTGAAAAAATTTGGAGAAAATTTTGCATCATGTCAAGCTGGAATATCCAGTTTTTACACAA;MAPQ=60;MATEID=1115328_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_182329001_182354001_323C;SPAN=4847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:84 GQ:43.4 PL:[43.4, 0.0, 158.9] SR:16 DR:9 LR:-43.26 LO:47.06);ALT=G[chr2:182344862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	182343552	+	chr2	182344862	+	.	5	7	1115336_1	9.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=1115336_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_2_182329001_182354001_323C;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:7 DR:5 LR:-9.119 LO:18.15);ALT=G[chr2:182344862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	182344994	+	chr2	182346323	+	.	2	23	1115345_1	60.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1115345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_182329001_182354001_83C;SPAN=1329;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:81 GQ:60.8 PL:[60.8, 0.0, 133.4] SR:23 DR:2 LR:-60.58 LO:62.17);ALT=G[chr2:182346323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	182387069	+	chr2	182388163	+	.	10	4	1115514_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1115514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_182378001_182403001_243C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:65 GQ:25.4 PL:[25.4, 0.0, 131.0] SR:4 DR:10 LR:-25.3 LO:29.46);ALT=G[chr2:182388163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	183028730	+	chr2	183029749	+	.	25	26	1117031_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=1117031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_183015001_183040001_226C;SPAN=1019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:74 GQ:65.9 PL:[112.1, 0.0, 65.9] SR:26 DR:25 LR:-112.6 LO:112.6);ALT=G[chr2:183029749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	183581212	+	chr2	183582666	+	ATATTTTTGTGGAATGAAAAGGAAGTATTAGAAATGAGCTGAAGACCATTCAC	0	18	1118129_1	42.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATATTTTTGTGGAATGAAAAGGAAGTATTAGAAATGAGCTGAAGACCATTCAC;MAPQ=60;MATEID=1118129_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_183578501_183603501_202C;SPAN=1454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:63 GQ:42.5 PL:[42.5, 0.0, 108.5] SR:18 DR:0 LR:-42.35 LO:44.03);ALT=T[chr2:183582666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	183583017	+	chr2	183584733	+	.	3	2	1118134_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1118134_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_183578501_183603501_296C;SPAN=1716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:2 DR:3 LR:4.677 LO:6.851);ALT=G[chr2:183584733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	183594669	+	chr2	183595755	+	.	0	5	1118179_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1118179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_183578501_183603501_280C;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:65 GQ:0.9 PL:[0.0, 0.9, 158.4] SR:5 DR:0 LR:1.105 LO:9.099);ALT=G[chr2:183595755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187351185	+	chr2	187359960	+	.	59	72	1126341_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1126341_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_187327001_187352001_151C;SPAN=8775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:57 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:72 DR:59 LR:-283.9 LO:283.9);ALT=G[chr2:187359960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187351190	+	chr2	187364906	+	.	20	0	1126343_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1126343_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:187351190(+)-2:187364906(-)__2_187327001_187352001D;SPAN=13716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:0 DR:20 LR:-52.2 LO:52.37);ALT=T[chr2:187364906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187360064	+	chr2	187364907	+	.	0	36	1126349_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AGGTA;MAPQ=60;MATEID=1126349_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CACA;SCTG=c_2_187327001_187352001_151C;SPAN=4843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:0 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:36 DR:0 LR:-105.6 LO:105.6);ALT=A[chr2:187364907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187367316	+	chr2	187368759	+	.	0	30	1126258_1	72.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=1126258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_187351501_187376501_181C;SPAN=1443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:99 GQ:72.2 PL:[72.2, 0.0, 167.9] SR:30 DR:0 LR:-72.21 LO:74.32);ALT=T[chr2:187368759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	187368941	+	chr2	187370176	+	.	12	4	1126267_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1126267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_187351501_187376501_89C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:78 GQ:21.8 PL:[21.8, 0.0, 167.0] SR:4 DR:12 LR:-21.78 LO:28.31);ALT=G[chr2:187370176[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	188296092	+	chr2	188312765	+	.	7	4	1128594_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1128594_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_188307001_188332001_351C;SPAN=16673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:52 GQ:12.5 PL:[12.5, 0.0, 111.5] SR:4 DR:7 LR:-12.32 LO:17.12);ALT=C[chr2:188312765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	188368553	+	chr2	188418987	+	.	9	0	1128903_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1128903_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:188368553(+)-2:188418987(-)__2_188405001_188430001D;SPAN=50434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:0 DR:9 LR:-16.16 LO:19.94);ALT=T[chr2:188418987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	188394212	+	chr2	188418926	+	.	0	8	1128723_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1128723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_188380501_188405501_121C;SPAN=24714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:8 DR:0 LR:-14.76 LO:17.85);ALT=C[chr2:188418926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	188649775	+	chr2	195455676	+	.	16	0	1129472_1	43.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=1129472_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:188649775(+)-2:195455676(-)__2_188625501_188650501D;SPAN=6805901;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:36 GQ:43.1 PL:[43.1, 0.0, 43.1] SR:0 DR:16 LR:-43.06 LO:43.06);ALT=G[chr2:195455676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	189119678	+	chr2	189120982	+	.	17	0	1130365_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1130365_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:189119678(+)-2:189120982(-)__2_189115501_189140501D;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.57 LO:43.16);ALT=C[chr2:189120982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	190306304	+	chr2	190313116	+	.	10	0	1132814_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1132814_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:190306304(+)-2:190313116(-)__2_190291501_190316501D;SPAN=6812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:0 DR:10 LR:-9.711 LO:20.09);ALT=A[chr2:190313116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	190426918	+	chr2	190428308	+	.	2	3	1133232_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1133232_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_190414001_190439001_286C;SPAN=1390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:61 GQ:3 PL:[0.0, 3.0, 151.8] SR:3 DR:2 LR:3.322 LO:6.992);ALT=C[chr2:190428308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	190647370	+	chr2	190648994	+	.	15	0	1133798_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1133798_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:190647370(+)-2:190648994(-)__2_190634501_190659501D;SPAN=1624;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:81 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:0 DR:15 LR:-27.57 LO:33.43);ALT=C[chr2:190648994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	190649313	+	chr2	190656513	+	.	13	0	1133802_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1133802_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:190649313(+)-2:190656513(-)__2_190634501_190659501D;SPAN=7200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:75 GQ:22.7 PL:[22.7, 0.0, 158.0] SR:0 DR:13 LR:-22.59 LO:28.56);ALT=C[chr2:190656513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	2788642	+	chr2	191184440	+	.	5	5	2402816_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTCGACATGAGCCTCC;MAPQ=60;MATEID=2402816_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_2768501_2793501_92C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:35 GQ:10.4 PL:[10.4, 0.0, 73.1] SR:5 DR:5 LR:-10.32 LO:13.15);ALT=]chr5:2788642]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	194324817	-	chr4	131114465	+	.	12	25	2207260_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=2207260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_131099501_131124501_350C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:30 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:25 DR:12 LR:-102.3 LO:102.3);ALT=[chr4:131114465[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	194545044	+	chr14	65447291	+	TTTTTTTTTTATTTTTATTTTTTTTTTTTTTTT	43	47	5775820_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TTTTA;INSERTION=TTTTTTTTTTATTTTTATTTTTTTTTTTTTTTT;MAPQ=60;MATEID=5775820_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_65439501_65464501_193C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:36 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:47 DR:43 LR:-224.5 LO:224.5);ALT=A[chr14:65447291[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	194689502	+	chr2	194698766	+	.	60	50	1142905_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1142905_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_194677001_194702001_27C;SPAN=9264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:25 GQ:24 PL:[264.0, 24.0, 0.0] SR:50 DR:60 LR:-264.1 LO:264.1);ALT=G[chr2:194698766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198051833	+	chr2	198175302	+	.	11	9	1150775_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=1150775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198156001_198181001_150C;SPAN=123469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:12 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:9 DR:11 LR:-42.91 LO:42.91);ALT=G[chr2:198175302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198115016	+	chr2	198175310	+	.	16	0	1150777_1	49.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1150777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198115016(+)-2:198175310(-)__2_198156001_198181001D;SPAN=60294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:17 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:16 LR:-49.51 LO:49.51);ALT=G[chr2:198175310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198261053	+	chr2	198262709	+	.	6	4	1151047_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1151047_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198254001_198279001_176C;SPAN=1656;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:4 DR:6 LR:-7.222 LO:17.79);ALT=C[chr2:198262709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198263309	+	chr2	198264774	+	.	7	3	1151056_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CATACCTAT;MAPQ=60;MATEID=1151056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198254001_198279001_11C;SPAN=1465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:3 DR:7 LR:-6.73 LO:19.53);ALT=T[chr2:198264774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198268513	+	chr2	198269798	+	.	21	0	1151071_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1151071_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198268513(+)-2:198269798(-)__2_198254001_198279001D;SPAN=1285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:69 GQ:50.6 PL:[50.6, 0.0, 116.6] SR:0 DR:21 LR:-50.63 LO:52.07);ALT=G[chr2:198269798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198270198	+	chr2	198273091	+	TATATCCTTCTGGGAACATAGCATCTAATTCCTCATCAGAAAGTGGGCGATTTCTCTCATCAATTTCTCTTTCCCACCGCCAAGCCTGAAGCTGTTCAGGAGTCATACTCATTATGTG	0	23	1151077_1	51.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=TATATCCTTCTGGGAACATAGCATCTAATTCCTCATCAGAAAGTGGGCGATTTCTCTCATCAATTTCTCTTTCCCACCGCCAAGCCTGAAGCTGTTCAGGAGTCATACTCATTATGTG;MAPQ=60;MATEID=1151077_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_198254001_198279001_304C;SPAN=2893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:89 GQ:51.8 PL:[51.8, 0.0, 164.0] SR:23 DR:0 LR:-51.81 LO:55.07);ALT=T[chr2:198273091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198270198	+	chr2	198272719	+	.	3	12	1151076_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TACCT;MAPQ=60;MATEID=1151076_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ATAT;SCTG=c_2_198254001_198279001_304C;SPAN=2521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:72 GQ:30.2 PL:[30.2, 0.0, 142.4] SR:12 DR:3 LR:-30.01 LO:34.3);ALT=T[chr2:198272719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198273307	+	chr2	198274494	+	.	4	3	1151086_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1151086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198254001_198279001_31C;SPAN=1187;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:3 DR:4 LR:0.1925 LO:12.92);ALT=T[chr2:198274494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198285857	+	chr2	198288531	+	.	5	36	1151294_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1151294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198278501_198303501_167C;SPAN=2674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:95 GQ:99 PL:[109.7, 0.0, 119.6] SR:36 DR:5 LR:-109.6 LO:109.6);ALT=C[chr2:198288531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198285908	+	chr2	198299692	+	.	26	0	1151295_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1151295_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198285908(+)-2:198299692(-)__2_198278501_198303501D;SPAN=13784;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:97 GQ:59.6 PL:[59.6, 0.0, 175.1] SR:0 DR:26 LR:-59.55 LO:62.74);ALT=A[chr2:198299692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198288700	+	chr2	198299696	+	.	37	12	1151306_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1151306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198278501_198303501_370C;SPAN=10996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:102 GQ:99 PL:[127.7, 0.0, 117.8] SR:12 DR:37 LR:-127.5 LO:127.5);ALT=T[chr2:198299696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198318388	+	chr2	198324653	+	.	9	8	1151406_1	26.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1151406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198303001_198328001_358C;SPAN=6265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:73 GQ:26.6 PL:[26.6, 0.0, 148.7] SR:8 DR:9 LR:-26.44 LO:31.44);ALT=G[chr2:198324653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198360415	+	chr2	198361606	+	.	0	6	1151930_1	0	.	EVDNC=ASSMB;HOMSEQ=CCTGGGCT;MAPQ=60;MATEID=1151930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_198352001_198377001_306C;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:90 GQ:4.5 PL:[0.0, 4.5, 227.7] SR:6 DR:0 LR:4.577 LO:10.53);ALT=T[chr2:198361606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	198362139	+	chr2	198364504	+	.	39	0	1151938_1	88.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=1151938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198362139(+)-2:198364504(-)__2_198352001_198377001D;SPAN=2365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:149 GQ:88.4 PL:[88.4, 0.0, 273.2] SR:0 DR:39 LR:-88.37 LO:93.64);ALT=G[chr2:198364504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	36810206	+	chr2	198364504	+	.	17	0	1151947_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1151947_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198364504(-)-3:36810206(+)__2_198352001_198377001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:99 GQ:29.3 PL:[29.3, 0.0, 210.8] SR:0 DR:17 LR:-29.3 LO:37.27);ALT=]chr3:36810206]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	198365192	+	chr14	64068293	+	.	29	0	1151960_1	82.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1151960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:198365192(+)-14:64068293(-)__2_198352001_198377001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:50 GQ:39.2 PL:[82.1, 0.0, 39.2] SR:0 DR:29 LR:-83.01 LO:83.01);ALT=A[chr14:64068293[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	200713715	+	chr2	200715473	+	.	14	0	1157026_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1157026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:200713715(+)-2:200715473(-)__2_200704001_200729001D;SPAN=1758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:0 DR:14 LR:-28.06 LO:32.03);ALT=A[chr2:200715473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201676743	+	chr2	201680061	+	.	55	0	1159312_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1159312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201676743(+)-2:201680061(-)__2_201659501_201684501D;SPAN=3318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:77 GQ:25.4 PL:[160.7, 0.0, 25.4] SR:0 DR:55 LR:-166.2 LO:166.2);ALT=C[chr2:201680061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201678004	+	chr2	201680062	+	.	0	28	1159316_1	71.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1159316_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_201659501_201684501_379C;SPAN=2058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:78 GQ:71.3 PL:[71.3, 0.0, 117.5] SR:28 DR:0 LR:-71.3 LO:71.93);ALT=G[chr2:201680062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201726207	+	chr2	201729313	+	.	8	0	1159397_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1159397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201726207(+)-2:201729313(-)__2_201708501_201733501D;SPAN=3106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=A[chr2:201729313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201726597	+	chr2	201729316	+	.	10	0	1159398_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1159398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201726597(+)-2:201729316(-)__2_201708501_201733501D;SPAN=2719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:96 GQ:7.1 PL:[7.1, 0.0, 224.9] SR:0 DR:10 LR:-7.001 LO:19.58);ALT=G[chr2:201729316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201746213	+	chr2	201752336	+	GTTGGATCTCCTGTTTGAACCATGAAACCCTTGATATTCCTATGAAATATACAGCCATTGTAGTAATTACTGGCACAAAGAGCCAAGAAATTCTCACATGTTTTGGGTGTCCTCTCACAGAAGACTTCAATTTTAATATCACCTACATCTGTATGCAGTGTCACAGA	0	19	1159569_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTGGATCTCCTGTTTGAACCATGAAACCCTTGATATTCCTATGAAATATACAGCCATTGTAGTAATTACTGGCACAAAGAGCCAAGAAATTCTCACATGTTTTGGGTGTCCTCTCACAGAAGACTTCAATTTTAATATCACCTACATCTGTATGCAGTGTCACAGA;MAPQ=60;MATEID=1159569_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_201733001_201758001_328C;SPAN=6123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:73 GQ:43.1 PL:[43.1, 0.0, 132.2] SR:19 DR:0 LR:-42.94 LO:45.56);ALT=T[chr2:201752336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201936814	+	chr2	201950180	+	.	19	0	1160233_1	42.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=1160233_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201936814(+)-2:201950180(-)__2_201929001_201954001D;SPAN=13366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:76 GQ:42.2 PL:[42.2, 0.0, 141.2] SR:0 DR:19 LR:-42.13 LO:45.17);ALT=A[chr2:201950180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201936830	+	chr2	201943601	+	.	17	0	1160234_1	33.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=1160234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:201936830(+)-2:201943601(-)__2_201929001_201954001D;SPAN=6771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:85 GQ:33.2 PL:[33.2, 0.0, 171.8] SR:0 DR:17 LR:-33.09 LO:38.53);ALT=A[chr2:201943601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201981204	+	chr2	201994451	+	.	4	4	1160301_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1160301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_201978001_202003001_188C;SPAN=13247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:4 DR:4 LR:-3.921 LO:15.38);ALT=G[chr2:201994451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	201983624	+	chr2	201994452	+	.	13	10	1160313_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1160313_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_201978001_202003001_335C;SPAN=10828;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:89 GQ:28.7 PL:[28.7, 0.0, 187.1] SR:10 DR:13 LR:-28.7 LO:35.43);ALT=C[chr2:201994452[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	202048032	+	chr2	202050492	+	.	10	9	1160530_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1160530_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_202027001_202052001_306C;SPAN=2460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:68 GQ:31.1 PL:[31.1, 0.0, 133.4] SR:9 DR:10 LR:-31.09 LO:34.72);ALT=G[chr2:202050492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	202125373	+	chr2	202131181	+	.	20	0	1161095_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1161095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:202125373(+)-2:202131181(-)__2_202100501_202125501D;SPAN=5808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:46 GQ:53.6 PL:[53.6, 0.0, 56.9] SR:0 DR:20 LR:-53.56 LO:53.57);ALT=T[chr2:202131181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	202146658	+	chr2	202149441	+	.	79	50	1160930_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCAAATTCTT;MAPQ=60;MATEID=1160930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_202149501_202174501_306C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:7 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:50 DR:79 LR:-333.4 LO:333.4);ALT=T[chr2:202149441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135347363	+	chr2	203104274	+	.	66	0	3621391_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=3621391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:203104274(-)-7:135347363(+)__7_135338001_135363001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:98 GQ:46.1 PL:[191.3, 0.0, 46.1] SR:0 DR:66 LR:-196.2 LO:196.2);ALT=]chr7:135347363]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	203130580	+	chr2	203139829	+	.	9	0	1163640_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1163640_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:203130580(+)-2:203139829(-)__2_203129501_203154501D;SPAN=9249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:77 GQ:8.9 PL:[8.9, 0.0, 177.2] SR:0 DR:9 LR:-8.848 LO:18.1);ALT=G[chr2:203139829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	203165090	+	chr2	203167642	+	.	3	7	1163502_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1163502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_203154001_203179001_156C;SPAN=2552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:7 DR:3 LR:-6.901 LO:15.9);ALT=G[chr2:203167642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	203638956	+	chr4	89444837	+	.	33	0	2080293_1	89.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=2080293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:203638956(+)-4:89444837(-)__4_89425001_89450001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:71 GQ:80 PL:[89.9, 0.0, 80.0] SR:0 DR:33 LR:-89.71 LO:89.71);ALT=T[chr4:89444837[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	203772682	+	chr2	203776159	+	.	0	10	1165659_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1165659_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_203766501_203791501_127C;SPAN=3477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:81 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:0 LR:-11.07 LO:20.36);ALT=T[chr2:203776159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	204103858	+	chr2	204110568	+	.	3	2	1166818_1	6.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1166818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_204109501_204134501_331C;SPAN=6710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:36 GQ:6.8 PL:[6.8, 0.0, 79.4] SR:2 DR:3 LR:-6.752 LO:10.46);ALT=G[chr2:204110568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	208474495	+	chr2	208476785	+	.	77	33	1177710_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGAAAACCTATTC;MAPQ=60;MATEID=1177710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_208470501_208495501_63C;SPAN=2290;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:35 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:33 DR:77 LR:-287.2 LO:287.2);ALT=C[chr2:208476785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209002677	+	chr10	13283671	+	AAAGTGCTAGGATTACAGGCATGCACCACCACATGTGGCTGGGGTCATTTTTTGAAACGTAAACATTGAAGGAGGTAGCACCCTATATCCTGATCTCTGTGGAAAGGTAGGGGCATGAATTCAGCAGACACCCTACTCTGAGTTGTGAGGACCAAACATAGTGGCCTATGATTACCAACCCCTGAAGCTCTTTAAACCACTCCAGCTCTTTAGTTCAGCAGAATCGAGCCCAGGTTCTCTCCTCTATTGCACAAGTCTTTTATTATTATTATTTTTAAAATAGAGACGGGGGT	12	60	4518281_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;HOMSEQ=CTCCTGGGCTCAAGCAATCCT;INSERTION=AAAGTGCTAGGATTACAGGCATGCACCACCACATGTGGCTGGGGTCATTTTTTGAAACGTAAACATTGAAGGAGGTAGCACCCTATATCCTGATCTCTGTGGAAAGGTAGGGGCATGAATTCAGCAGACACCCTACTCTGAGTTGTGAGGACCAAACATAGTGGCCTATGATTACCAACCCCTGAAGCTCTTTAAACCACTCCAGCTCTTTAGTTCAGCAGAATCGAGCCCAGGTTCTCTCCTCTATTGCACAAGTCTTTTATTATTATTATTTTTAAAATAGAGACGGGGGT;MAPQ=60;MATEID=4518281_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_13279001_13304001_174C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:53 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:60 DR:12 LR:-184.8 LO:184.8);ALT=T[chr10:13283671[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	209033773	+	chr17	19995679	-	.	39	0	6342394_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6342394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:209033773(+)-17:19995679(+)__17_19992001_20017001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:32 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:39 LR:-115.5 LO:115.5);ALT=T]chr17:19995679];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	209116293	+	chr2	209118608	+	.	0	29	1179607_1	71.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=1179607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_209107501_209132501_362C;SPAN=2315;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:91 GQ:71.3 PL:[71.3, 0.0, 147.2] SR:29 DR:0 LR:-71.08 LO:72.62);ALT=T[chr2:209118608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209116339	+	chr2	209119695	+	.	26	0	1179609_1	63.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=1179609_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:209116339(+)-2:209119695(-)__2_209107501_209132501D;SPAN=3356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:83 GQ:63.5 PL:[63.5, 0.0, 136.1] SR:0 DR:26 LR:-63.34 LO:64.87);ALT=A[chr2:209119695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209131139	+	chr2	209136232	+	.	34	20	1179659_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1179659_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_209132001_209157001_38C;SPAN=5093;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:52 GQ:2.6 PL:[121.4, 0.0, 2.6] SR:20 DR:34 LR:-127.7 LO:127.7);ALT=G[chr2:209136232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	209191156	+	chr2	209192902	+	.	2	5	1179829_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=1179829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_209181001_209206001_285C;SPAN=1746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:89 GQ:4.2 PL:[0.0, 4.2, 224.4] SR:5 DR:2 LR:4.306 LO:10.56);ALT=G[chr2:209192902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216176920	+	chr2	216182875	+	.	22	0	1195689_1	55.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1195689_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:216176920(+)-2:216182875(-)__2_216163501_216188501D;SPAN=5955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:63 GQ:55.7 PL:[55.7, 0.0, 95.3] SR:0 DR:22 LR:-55.55 LO:56.18);ALT=C[chr2:216182875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216177347	+	chr2	216182876	+	.	0	24	1195691_1	57.0	.	EVDNC=ASSMB;HOMSEQ=TCAG;MAPQ=60;MATEID=1195691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_216163501_216188501_62C;SPAN=5529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:81 GQ:57.5 PL:[57.5, 0.0, 136.7] SR:24 DR:0 LR:-57.28 LO:59.17);ALT=G[chr2:216182876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216203630	+	chr2	216209502	+	.	3	5	1195547_1	3.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=1195547_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_216188001_216213001_324C;SPAN=5872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:72 GQ:3.8 PL:[3.8, 0.0, 168.8] SR:5 DR:3 LR:-3.6 LO:13.48);ALT=T[chr2:216209502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216211665	+	chr2	216213815	+	.	3	2	1195576_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1195576_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_216188001_216213001_122C;SPAN=2150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:50 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:2 DR:3 LR:0.3422 LO:7.35);ALT=G[chr2:216213815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216845659	+	chr17	8650195	-	.	11	12	6306999_1	52.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=TTCCCTTCCCTTCCCT;MAPQ=57;MATEID=6306999_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_8648501_8673501_176C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:12 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:12 DR:11 LR:-52.81 LO:52.81);ALT=A]chr17:8650195];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	216974181	+	chr2	216990638	+	CAGCTGTTGTGCTGTGTATGGACGTGGGCTTTACCATGAGTAACTCCATTCCTGGTATAGAATCCCCATTTGAACAAGCAAAGAAGGTGATAACCATGTTTGTACAGCGACAGGTGTTTGCTGAGAACAAGGATGAGATTGCTTTAGTCCTGTTTGGTACAGATGGCACTGACAATCCCCTTTCTGGTGGGGATCAGTATCAGAACATCACAGTGCACAGACATCTGATGCTACCAGATTTTGATTTGCTGGAGGACATTGAAAGCAAAATCCAACCAGGTTCTCAACAGGCTGACTTCCTGGATGCACTAATCGTGAGCATGGATGTGATTCAACATGAAACAATAGGAAAGAAGTTTGAGAAGAGGCATATTGAAATATTCACTGACCTCAGCAGCCGATTCAGCAAAAGTCAGCTGGATATTATAATTCATAGCTTGAAGAAATGTGACATCTCCCTGCAATTCTTCTTGCCTTTCTCACTTGGCAAGGAAGATGGAAGTGGGGACAGAGGAGATGGCCCCTTTCGCTTAGGTGGCCATGGGCCTTCCTTTCCACTAAAAGGAATTACCGAACAGCAAAAAGAAGGTCTTGAGATAGTGAAAATGGTGATGATATCTTTAGAAGGTGAAGATGGGTTGGATGAAATTTATTCATTC	0	30	1198043_1	76.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAGCTGTTGTGCTGTGTATGGACGTGGGCTTTACCATGAGTAACTCCATTCCTGGTATAGAATCCCCATTTGAACAAGCAAAGAAGGTGATAACCATGTTTGTACAGCGACAGGTGTTTGCTGAGAACAAGGATGAGATTGCTTTAGTCCTGTTTGGTACAGATGGCACTGACAATCCCCTTTCTGGTGGGGATCAGTATCAGAACATCACAGTGCACAGACATCTGATGCTACCAGATTTTGATTTGCTGGAGGACATTGAAAGCAAAATCCAACCAGGTTCTCAACAGGCTGACTTCCTGGATGCACTAATCGTGAGCATGGATGTGATTCAACATGAAACAATAGGAAAGAAGTTTGAGAAGAGGCATATTGAAATATTCACTGACCTCAGCAGCCGATTCAGCAAAAGTCAGCTGGATATTATAATTCATAGCTTGAAGAAATGTGACATCTCCCTGCAATTCTTCTTGCCTTTCTCACTTGGCAAGGAAGATGGAAGTGGGGACAGAGGAGATGGCCCCTTTCGCTTAGGTGGCCATGGGCCTTCCTTTCCACTAAAAGGAATTACCGAACAGCAAAAAGAAGGTCTTGAGATAGTGAAAATGGTGATGATATCTTTAGAAGGTGAAGATGGGTTGGATGAAATTTATTCATTC;MAPQ=60;MATEID=1198043_2;MATENM=0;NM=0;NUMPARTS=7;SCTG=c_2_216972001_216997001_267C;SPAN=16457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:85 GQ:76.1 PL:[76.1, 0.0, 128.9] SR:30 DR:0 LR:-76.0 LO:76.78);ALT=G[chr2:216990638[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216974181	+	chr2	216977737	+	.	35	9	1198042_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=1198042_2;MATENM=0;NM=0;NUMPARTS=7;REPSEQ=GG;SCTG=c_2_216972001_216997001_267C;SPAN=3556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:103 GQ:99 PL:[110.9, 0.0, 137.3] SR:9 DR:35 LR:-110.7 LO:110.9);ALT=G[chr2:216977737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216974226	+	chr2	216981379	+	.	36	0	1198045_1	91.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1198045_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:216974226(+)-2:216981379(-)__2_216972001_216997001D;SPAN=7153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:102 GQ:91.4 PL:[91.4, 0.0, 154.1] SR:0 DR:36 LR:-91.2 LO:92.14);ALT=C[chr2:216981379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216977854	+	chr2	216981380	+	.	4	56	1198052_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=1198052_2;MATENM=0;NM=0;NUMPARTS=7;REPSEQ=TTT;SCTG=c_2_216972001_216997001_267C;SPAN=3526;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:121 GQ:99 PL:[158.9, 0.0, 132.5] SR:56 DR:4 LR:-158.8 LO:158.8);ALT=T[chr2:216981380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	216983888	+	chr2	216986785	+	.	8	7	1198065_1	28.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=1198065_2;MATENM=0;NM=0;NUMPARTS=7;REPSEQ=TT;SCTG=c_2_216972001_216997001_267C;SPAN=2897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:79 GQ:28.1 PL:[28.1, 0.0, 163.4] SR:7 DR:8 LR:-28.11 LO:33.61);ALT=T[chr2:216986785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217057458	+	chr2	217059641	+	.	2	6	1198007_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1198007_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_2_217045501_217070501_210C;SPAN=2183;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:6 DR:2 LR:1.005 LO:12.81);ALT=G[chr2:217059641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217057458	+	chr2	217069043	+	ATGGAATTACTCTGATCACCAAAGAGGAAGCCTCTGGAAGTTCTGTCACAGCTGAGGAAGCCAAAA	4	17	1198008_1	34.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATGGAATTACTCTGATCACCAAAGAGGAAGCCTCTGGAAGTTCTGTCACAGCTGAGGAAGCCAAAA;MAPQ=60;MATEID=1198008_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_217045501_217070501_210C;SPAN=11585;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:79 GQ:34.7 PL:[34.7, 0.0, 156.8] SR:17 DR:4 LR:-34.71 LO:39.14);ALT=G[chr2:217069043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217089943	+	chr2	217092499	+	.	79	45	1198277_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GCCATGTGTTCTT;MAPQ=60;MATEID=1198277_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_2_217070001_217095001_328C;SPAN=2556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:322 GQ:99 PL:[249.7, 0.0, 530.3] SR:45 DR:79 LR:-249.5 LO:255.1);ALT=T[chr2:217092499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217089968	+	chr2	217093111	+	.	9	0	1198278_1	0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=1198278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:217089968(+)-2:217093111(-)__2_217070001_217095001D;SPAN=3143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:472 GQ:97.8 PL:[0.0, 97.8, 1340.0] SR:0 DR:9 LR:98.17 LO:10.86);ALT=T[chr2:217093111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	217475711	+	chr17	36909097	-	.	15	0	6386400_1	40.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6386400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:217475711(+)-17:36909097(+)__17_36897001_36922001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:35 GQ:40.1 PL:[40.1, 0.0, 43.4] SR:0 DR:15 LR:-40.03 LO:40.05);ALT=T]chr17:36909097];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	217955896	+	chr2	217957267	+	.	41	33	1200419_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTGG;MAPQ=60;MATEID=1200419_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_217952001_217977001_18C;SPAN=1371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:45 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:33 DR:41 LR:-184.8 LO:184.8);ALT=G[chr2:217957267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219081977	+	chr2	219104114	+	CCGCCGCCATGATCCTGCTGGAGGTGAACAACCGCATCATCGAGGAGACGCTCGCGCTCAAGTTCGAGAACGCGGCCGCCGGAAACAAACCGGAAGCAGTAGAAGTAACATTTGCAGATTTCGATGGGGTCCTCTATCATATTTCAAATCCTAATGGAGACAAAACAAAAGTGATGGTCAGTATTTCTTTGAAATTCTACAAGGAACTTCAGGCACATGGTGCTGATGAGTTATTAAAGAGGGTGTACGGGAGTTTCTTGGTAAATCCAGAATCAGGATACAATGTCTCTTTGCTATATGACCTTGAAAATCTTCCGGCATCCAAGGATTCCATTGTGCATCAAGCTGGCATGTTGAAGCGAAATTGTTTTGCCTCTGTCTTTGAAAAATACTTCCAATTCCAAGAAGAGGGCAAGGAAGGAGAGAACAGGGCAGTTATCCATTATAGGGATGATGAGACCAT	2	33	1203179_1	78.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=CCGCCGCCATGATCCTGCTGGAGGTGAACAACCGCATCATCGAGGAGACGCTCGCGCTCAAGTTCGAGAACGCGGCCGCCGGAAACAAACCGGAAGCAGTAGAAGTAACATTTGCAGATTTCGATGGGGTCCTCTATCATATTTCAAATCCTAATGGAGACAAAACAAAAGTGATGGTCAGTATTTCTTTGAAATTCTACAAGGAACTTCAGGCACATGGTGCTGATGAGTTATTAAAGAGGGTGTACGGGAGTTTCTTGGTAAATCCAGAATCAGGATACAATGTCTCTTTGCTATATGACCTTGAAAATCTTCCGGCATCCAAGGATTCCATTGTGCATCAAGCTGGCATGTTGAAGCGAAATTGTTTTGCCTCTGTCTTTGAAAAATACTTCCAATTCCAAGAAGAGGGCAAGGAAGGAGAGAACAGGGCAGTTATCCATTATAGGGATGATGAGACCAT;MAPQ=60;MATEID=1203179_2;MATENM=0;NM=0;NUMPARTS=7;SCTG=c_2_219079001_219104001_51C;SPAN=22137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:138 GQ:78.2 PL:[78.2, 0.0, 256.4] SR:33 DR:2 LR:-78.15 LO:83.47);ALT=G[chr2:219104114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219082015	+	chr2	219099072	+	.	11	0	1203181_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1203181_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219082015(+)-2:219099072(-)__2_219079001_219104001D;SPAN=17057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:136 GQ:0.3 PL:[0.0, 0.3, 330.0] SR:0 DR:11 LR:0.5347 LO:20.27);ALT=C[chr2:219099072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219082086	+	chr2	219093456	+	.	104	0	1203182_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1203182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219082086(+)-2:219093456(-)__2_219079001_219104001D;SPAN=11370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:104 DP:160 GQ:88.7 PL:[299.9, 0.0, 88.7] SR:0 DR:104 LR:-306.3 LO:306.3);ALT=C[chr2:219093456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219093521	+	chr2	219104113	+	.	2	3	1203441_1	4.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1203441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219103501_219128501_345C;SPAN=10592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:44 GQ:4.7 PL:[4.7, 0.0, 100.4] SR:3 DR:2 LR:-4.584 LO:9.99);ALT=T[chr2:219104113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219103622	+	chr2	219110138	+	.	11	0	1203448_1	11.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1203448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219103622(+)-2:219110138(-)__2_219103501_219128501D;SPAN=6516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:91 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:0 DR:11 LR:-11.66 LO:22.29);ALT=C[chr2:219110138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219104208	+	chr2	219110139	+	.	15	27	1203450_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GCAGG;MAPQ=60;MATEID=1203450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219103501_219128501_268C;SPAN=5931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:97 GQ:99 PL:[105.8, 0.0, 128.9] SR:27 DR:15 LR:-105.8 LO:105.9);ALT=G[chr2:219110139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219104258	+	chr2	219114085	+	.	12	0	1203451_1	11.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1203451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219104258(+)-2:219114085(-)__2_219103501_219128501D;SPAN=9827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:106 GQ:11 PL:[11.0, 0.0, 245.3] SR:0 DR:12 LR:-10.89 LO:23.95);ALT=T[chr2:219114085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219110269	+	chr2	219114542	+	TGCTGTTCCCTCGTCACACCAATGCCAGTGCTCGAGACAACACCATCAACCTGATCCACACGTTCCGGGACTACCTGCACTACCACATCAAGTGCTCTA	13	154	1203468_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TGCTGTTCCCTCGTCACACCAATGCCAGTGCTCGAGACAACACCATCAACCTGATCCACACGTTCCGGGACTACCTGCACTACCACATCAAGTGCTCTA;MAPQ=60;MATEID=1203468_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_219103501_219128501_31C;SPAN=4273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:161 DP:132 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:154 DR:13 LR:-475.3 LO:475.3);ALT=G[chr2:219114542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219110322	+	chr2	219114085	+	.	12	0	1203469_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1203469_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219110322(+)-2:219114085(-)__2_219103501_219128501D;SPAN=3763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:101 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:0 DR:12 LR:-12.25 LO:24.22);ALT=A[chr2:219114085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219114213	+	chr2	219118613	+	.	12	0	1203482_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1203482_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219114213(+)-2:219118613(-)__2_219103501_219128501D;SPAN=4400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:147 GQ:0 PL:[0.0, 0.0, 356.4] SR:0 DR:12 LR:0.2139 LO:22.16);ALT=C[chr2:219118613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219114645	+	chr2	219118614	+	.	30	86	1203484_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1203484_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219103501_219128501_77C;SPAN=3969;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:165 GQ:77.6 PL:[321.8, 0.0, 77.6] SR:86 DR:30 LR:-330.0 LO:330.0);ALT=G[chr2:219118614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219131711	+	chr2	219134105	+	GCACACTCAAAGAGCAGCTCCCCATCGCTGAGCCGCCATACGAAGGCTTTGTCATCTTCACCCCCGGTCACTGCCAAGGTATTGGTCTTGGGGTCCAGGCTCACACAAAACACAGATG	3	11	1203272_1	22.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GCACACTCAAAGAGCAGCTCCCCATCGCTGAGCCGCCATACGAAGGCTTTGTCATCTTCACCCCCGGTCACTGCCAAGGTATTGGTCTTGGGGTCCAGGCTCACACAAAACACAGATG;MAPQ=60;MATEID=1203272_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_219128001_219153001_233C;SPAN=2394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:65 GQ:22.1 PL:[22.1, 0.0, 134.3] SR:11 DR:3 LR:-22.0 LO:26.73);ALT=T[chr2:219134105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219132339	+	chr2	219134105	+	.	4	5	1203273_1	12.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=1203273_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_219128001_219153001_233C;SPAN=1766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:5 DR:4 LR:-12.1 LO:18.81);ALT=G[chr2:219134105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219135336	+	chr2	219137294	+	.	13	0	1203280_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1203280_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219135336(+)-2:219137294(-)__2_219128001_219153001D;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:95 GQ:17.3 PL:[17.3, 0.0, 212.0] SR:0 DR:13 LR:-17.18 LO:27.1);ALT=G[chr2:219137294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219144850	+	chr2	219146662	+	.	0	7	1203312_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1203312_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_2_219128001_219153001_317C;SPAN=1812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:7 DR:0 LR:-2.788 LO:13.35);ALT=C[chr2:219146662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219146907	+	chr2	219157188	+	.	29	12	1203348_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=1203348_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_219152501_219177501_148C;SPAN=10281;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:36 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:12 DR:29 LR:-104.7 LO:104.7);ALT=G[chr2:219157188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219188156	+	chr2	219204505	+	.	9	7	1204241_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1204241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219177001_219202001_100C;SPAN=16349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:35 GQ:30.2 PL:[30.2, 0.0, 53.3] SR:7 DR:9 LR:-30.13 LO:30.52);ALT=T[chr2:219204505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219264882	+	chr2	219266285	+	.	9	3	1203642_1	16.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1203642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219250501_219275501_362C;SPAN=1403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:3 DR:9 LR:-16.48 LO:21.7);ALT=T[chr2:219266285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219275809	+	chr2	219276877	-	.	8	0	1203774_1	10.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1203774_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:219275809(+)-2:219276877(+)__2_219275001_219300001D;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-9.882 LO:16.52);ALT=A]chr2:219276877];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	219433701	+	chr2	219445283	+	.	4	3	1204514_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1204514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_219422001_219447001_272C;SPAN=11582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:89 GQ:7.5 PL:[0.0, 7.5, 231.0] SR:3 DR:4 LR:7.607 LO:8.395);ALT=G[chr2:219445283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	219797359	+	chr7	37333349	+	.	4	14	3256124_1	52.0	.	DISC_MAPQ=18;EVDNC=ASDIS;HOMSEQ=AAAA;MAPQ=60;MATEID=3256124_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_37313501_37338501_83C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:14 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:14 DR:4 LR:-52.81 LO:52.81);ALT=A[chr7:37333349[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	220023085	+	chr2	220025442	+	.	6	2	1206333_1	0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1206333_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_220010001_220035001_111C;SPAN=2357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:94 GQ:5.4 PL:[0.0, 5.4, 237.6] SR:2 DR:6 LR:5.661 LO:10.42);ALT=C[chr2:220025442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	220052366	+	chr2	220056242	+	.	11	0	1206271_1	22.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1206271_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:220052366(+)-2:220056242(-)__2_220034501_220059501D;SPAN=3876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:52 GQ:22.4 PL:[22.4, 0.0, 101.6] SR:0 DR:11 LR:-22.22 LO:25.23);ALT=C[chr2:220056242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	220239746	+	chr2	220246056	+	.	4	9	1207273_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1207273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_220230501_220255501_242C;SPAN=6310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:80 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:9 DR:4 LR:-17.94 LO:25.53);ALT=T[chr2:220246056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	221278223	-	chr5	39787751	+	C	8	25	2458234_1	94.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=2458234_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_39763501_39788501_132C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:42 GQ:5.3 PL:[94.4, 0.0, 5.3] SR:25 DR:8 LR:-98.59 LO:98.59);ALT=[chr5:39787751[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	221616224	-	chr2	221617278	+	.	8	0	1210464_1	3.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=1210464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:221616224(-)-2:221617278(-)__2_221602501_221627501D;SPAN=1054;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:0 DR:8 LR:-3.379 LO:15.29);ALT=[chr2:221617278[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr2	222809057	-	chr12	66524482	+	.	9	0	5229061_1	15.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=5229061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:222809057(-)-12:66524482(-)__12_66517501_66542501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:52 GQ:15.8 PL:[15.8, 0.0, 108.2] SR:0 DR:9 LR:-15.62 LO:19.77);ALT=[chr12:66524482[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	222826521	-	chr5	137910933	+	.	19	0	2592707_1	51.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2592707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:222826521(-)-5:137910933(-)__5_137910501_137935501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:40 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:0 DR:19 LR:-51.91 LO:51.91);ALT=[chr5:137910933[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr2	223507724	+	chr2	223520735	+	AATTTCATCAAGCTCCAGACCAAATTCAAAACATAGTTCATCAAATTCTTCGTCAG	14	9	1215007_1	57.0	.	DISC_MAPQ=58;EVDNC=TSI_G;INSERTION=AATTTCATCAAGCTCCAGACCAAATTCAAAACATAGTTCATCAAATTCTTCGTCAG;MAPQ=60;MATEID=1215007_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_223513501_223538501_11C;SPAN=13011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:43 GQ:44.6 PL:[57.8, 0.0, 44.6] SR:9 DR:14 LR:-57.73 LO:57.73);ALT=T[chr2:223520735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	223513514	+	chr2	223520735	+	.	6	6	1215009_1	6.0	.	DISC_MAPQ=58;EVDNC=TSI_L;MAPQ=60;MATEID=1215009_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_223513501_223538501_11C;SPAN=7221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:6 DR:6 LR:-6.139 LO:17.59);ALT=G[chr2:223520735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	223760191	+	chr2	223762672	+	.	28	17	1215833_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACTTTGTTCTTT;MAPQ=60;MATEID=1215833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_223758501_223783501_345C;SPAN=2481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:51 GQ:9.5 PL:[111.8, 0.0, 9.5] SR:17 DR:28 LR:-116.3 LO:116.3);ALT=T[chr2:223762672[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	224039700	+	chr9	109426677	+	.	24	21	4381014_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=4381014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_109417001_109442001_253C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:46 GQ:5.7 PL:[122.1, 5.7, 0.0] SR:21 DR:24 LR:-124.8 LO:124.8);ALT=T[chr9:109426677[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	109426854	+	chr2	224039705	+	AAATTTTAAAATTTAAAATATAAAG	20	32	4381015_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAATTTTAAAATTTAAAATATAAAG;MAPQ=60;MATEID=4381015_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_109417001_109442001_87C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:35 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:32 DR:20 LR:-128.7 LO:128.7);ALT=]chr9:109426854]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	224315277	+	chr2	224316406	-	.	8	0	1217126_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1217126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:224315277(+)-2:224316406(+)__2_224297501_224322501D;SPAN=1129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=C]chr2:224316406];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	224822368	+	chr2	224824250	+	.	0	18	1218478_1	36.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1218478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_224812001_224837001_82C;SPAN=1882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:84 GQ:36.8 PL:[36.8, 0.0, 165.5] SR:18 DR:0 LR:-36.66 LO:41.41);ALT=G[chr2:224824250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	228067531	+	chr6	29903883	-	CAC	2	6	1226378_1	16.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=CAC;MAPQ=60;MATEID=1226378_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_228046001_228071001_312C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:6 DP:2 GQ:1.5 PL:[16.5, 1.5, 0.0] SR:6 DR:2 LR:-16.5 LO:16.5);ALT=A]chr6:29903883];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	228190086	+	chr2	228195334	+	.	11	0	1226773_1	26.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=1226773_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:228190086(+)-2:228195334(-)__2_228193001_228218001D;SPAN=5248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:0 DR:11 LR:-26.29 LO:27.14);ALT=A[chr2:228195334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	228190144	+	chr2	228193393	+	.	21	25	1226762_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=17;MATEID=1226762_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_228168501_228193501_298C;SPAN=3249;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:101 GQ:99 PL:[108.2, 0.0, 134.6] SR:25 DR:21 LR:-108.0 LO:108.2);ALT=G[chr2:228193393[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	228190144	+	chr2	228197134	+	.	0	8	1226776_1	15.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=1226776_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_228193001_228218001_71C;SPAN=6990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:8 DR:0 LR:-15.03 LO:17.94);ALT=G[chr2:228197134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	228258379	+	chr2	228241100	+	.	51	23	1227072_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CACTTT;MAPQ=60;MATEID=1227072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_228242001_228267001_31C;SPAN=17279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:40 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:23 DR:51 LR:-191.4 LO:191.4);ALT=]chr2:228258379]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	230877120	+	chr2	230879677	+	.	69	49	1233472_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCTG;MAPQ=60;MATEID=1233472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_230863501_230888501_111C;SPAN=2557;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:62 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:49 DR:69 LR:-270.7 LO:270.7);ALT=G[chr2:230879677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231072776	+	chr2	231077062	+	TTCTTGTCTGAAGGTGTGCTGGACACCTCCTGGGGCTCTTCTGGGTCATTTGGTTCTGGAGAATTATCTCTTATCTCTGGCATAGAGCCCAAGGGAGAGTGGGGCATCTCTTGAGGGTCTTCTTTATCTCTTATTTGGGGGATCAGGTTGTCACTGGCCA	0	33	1234207_1	88.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTCTTGTCTGAAGGTGTGCTGGACACCTCCTGGGGCTCTTCTGGGTCATTTGGTTCTGGAGAATTATCTCTTATCTCTGGCATAGAGCCCAAGGGAGAGTGGGGCATCTCTTGAGGGTCTTCTTTATCTCTTATTTGGGGGATCAGGTTGTCACTGGCCA;MAPQ=60;MATEID=1234207_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_231059501_231084501_316C;SPAN=4286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:77 GQ:88.1 PL:[88.1, 0.0, 98.0] SR:33 DR:0 LR:-88.07 LO:88.11);ALT=T[chr2:231077062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231077743	+	chr2	231079665	+	.	2	5	1234220_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1234220_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_231059501_231084501_33C;SPAN=1922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:5 DR:2 LR:1.005 LO:12.81);ALT=C[chr2:231079665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231081645	+	chr2	231084588	+	.	25	8	1234283_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1234283_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231084001_231109001_124C;SPAN=2943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:26 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:8 DR:25 LR:-75.92 LO:75.92);ALT=T[chr2:231084588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231192000	+	chr2	231222517	+	.	9	0	1234621_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1234621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231192000(+)-2:231222517(-)__2_231182001_231207001D;SPAN=30517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:36 GQ:20 PL:[20.0, 0.0, 66.2] SR:0 DR:9 LR:-19.96 LO:21.4);ALT=A[chr2:231222517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231192017	+	chr2	231193470	+	.	5	4	1234622_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1234622_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231182001_231207001_187C;SPAN=1453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:65 GQ:5.6 PL:[5.6, 0.0, 150.8] SR:4 DR:5 LR:-5.497 LO:13.81);ALT=G[chr2:231193470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231193547	+	chr2	231222518	+	.	0	7	1234623_1	15.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1234623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231182001_231207001_290C;SPAN=28971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:27 GQ:15.8 PL:[15.8, 0.0, 48.8] SR:7 DR:0 LR:-15.79 LO:16.77);ALT=G[chr2:231222518[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231281044	+	chr2	231282304	+	.	14	9	1234795_1	28.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1234795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231280001_231305001_176C;SPAN=1260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:78 GQ:28.4 PL:[28.4, 0.0, 160.4] SR:9 DR:14 LR:-28.38 LO:33.71);ALT=G[chr2:231282304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231281045	+	chr2	231307648	+	.	19	0	1234796_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1234796_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231281045(+)-2:231307648(-)__2_231280001_231305001D;SPAN=26603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:41 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:0 DR:19 LR:-51.62 LO:51.62);ALT=T[chr2:231307648[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231282381	+	chr2	231307650	+	.	0	19	1234798_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1234798_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231280001_231305001_258C;SPAN=25269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:47 GQ:50 PL:[50.0, 0.0, 63.2] SR:19 DR:0 LR:-49.99 LO:50.08);ALT=G[chr2:231307650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231307815	+	chr2	231308893	+	.	2	3	1234738_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1234738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231304501_231329501_22C;SPAN=1078;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:59 GQ:0.5 PL:[0.5, 0.0, 142.4] SR:3 DR:2 LR:-0.5205 LO:9.318);ALT=G[chr2:231308893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231729788	+	chr2	231738130	+	.	53	0	1235889_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1235889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231729788(+)-2:231738130(-)__2_231721001_231746001D;SPAN=8342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:92 GQ:71 PL:[150.2, 0.0, 71.0] SR:0 DR:53 LR:-151.5 LO:151.5);ALT=C[chr2:231738130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231729911	+	chr2	231740324	+	.	10	0	1235892_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1235892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231729911(+)-2:231740324(-)__2_231721001_231746001D;SPAN=10413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:66 GQ:15.2 PL:[15.2, 0.0, 143.9] SR:0 DR:10 LR:-15.13 LO:21.33);ALT=C[chr2:231740324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231738272	+	chr2	231740332	+	.	0	17	1235916_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1235916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_231721001_231746001_324C;SPAN=2060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:73 GQ:36.5 PL:[36.5, 0.0, 138.8] SR:17 DR:0 LR:-36.34 LO:39.81);ALT=G[chr2:231740332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231921720	+	chr2	231926955	+	.	15	0	1236238_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1236238_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:231921720(+)-2:231926955(-)__2_231917001_231942001D;SPAN=5235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:83 GQ:27.2 PL:[27.2, 0.0, 172.4] SR:0 DR:15 LR:-27.03 LO:33.26);ALT=G[chr2:231926955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231921755	+	chr2	231927220	+	CTGGAATTATTTCTCTTCTGGATGAAGATGAACCACAGCTTAAGGAATTTGCACTACACAAATTGAATGCAGTTGTTAATGACTTCTGGGCAGAAATTTCCGAGTCCGTAGACAAAAT	0	27	1236240_1	66.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTGGAATTATTTCTCTTCTGGATGAAGATGAACCACAGCTTAAGGAATTTGCACTACACAAATTGAATGCAGTTGTTAATGACTTCTGGGCAGAAATTTCCGAGTCCGTAGACAAAAT;MAPQ=60;MATEID=1236240_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_231917001_231942001_135C;SPAN=5465;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:84 GQ:66.5 PL:[66.5, 0.0, 135.8] SR:27 DR:0 LR:-66.37 LO:67.73);ALT=G[chr2:231927220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	231921755	+	chr2	231925980	+	.	3	10	1236239_1	9.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1236239_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_231917001_231942001_135C;SPAN=4225;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:10 DR:3 LR:-9.169 LO:19.98);ALT=G[chr2:231925980[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232018382	+	chr2	232026051	+	.	3	4	1236535_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=1236535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_232015001_232040001_144C;SPAN=7669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:4 DR:3 LR:0.1925 LO:12.92);ALT=T[chr2:232026051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232026223	+	chr2	232028347	+	.	2	11	1236550_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1236550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_232015001_232040001_269C;SPAN=2124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:11 DR:2 LR:-13.55 LO:22.7);ALT=G[chr2:232028347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232321836	+	chr2	232322976	+	ACTCCAAGTGCTATTCTTTCCACCTCTATAGTCTTGATTTTGACCTTTCTCTCCAGTATAGTACAGGGAAATAGATCGCCCATCGATCTCTGTTCCCTGCTTTTCTTCAAAGGTTTTCTCTGCATCAGCTTCTGTCTTAAATTCAATATAAGCAAT	3	18	1237710_1	44.0	.	DISC_MAPQ=49;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=ACTCCAAGTGCTATTCTTTCCACCTCTATAGTCTTGATTTTGACCTTTCTCTCCAGTATAGTACAGGGAAATAGATCGCCCATCGATCTCTGTTCCCTGCTTTTCTTCAAAGGTTTTCTCTGCATCAGCTTCTGTCTTAAATTCAATATAAGCAAT;MAPQ=60;MATEID=1237710_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_232309001_232334001_165C;SPAN=1140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:78 GQ:44.9 PL:[44.9, 0.0, 143.9] SR:18 DR:3 LR:-44.89 LO:47.81);ALT=C[chr2:232322976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232323838	+	chr2	232324862	+	.	10	27	1237721_1	81.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1237721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_232309001_232334001_204C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:103 GQ:81.2 PL:[81.2, 0.0, 167.0] SR:27 DR:10 LR:-81.03 LO:82.73);ALT=T[chr2:232324862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232323883	+	chr2	232325187	+	.	13	0	1237722_1	18.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=1237722_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232323883(+)-2:232325187(-)__2_232309001_232334001D;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=A[chr2:232325187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232326730	+	chr2	232327909	+	.	27	91	1237733_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=1237733_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_2_232309001_232334001_332C;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:136 GQ:6.9 PL:[343.2, 6.9, 0.0] SR:91 DR:27 LR:-358.6 LO:358.6);ALT=T[chr2:232327909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232326730	+	chr2	232329046	+	CTTCTCCACTGCTATCATCTTCTTCATCTTCTGACATTTCCTCATCTTCACTATCTTCTTCTACCTCCTTTGGAGGAGGAGCCATTTTCTTGGGGTCACCTTGATTTTTACCTG	49	162	1237734_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTTCTCCACTGCTATCATCTTCTTCATCTTCTGACATTTCCTCATCTTCACTATCTTCTTCTACCTCCTTTGGAGGAGGAGCCATTTTCTTGGGGTCACCTTGATTTTTACCTG;MAPQ=60;MATEID=1237734_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_232309001_232334001_332C;SPAN=2316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:181 DP:130 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:162 DR:49 LR:-534.7 LO:534.7);ALT=T[chr2:232329046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232328079	+	chr2	232329114	+	.	106	0	1237741_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1237741_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232328079(+)-2:232329114(-)__2_232309001_232334001D;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:99 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=A[chr2:232329114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	232603948	+	chr2	232645896	+	.	15	0	1238672_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1238672_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:232603948(+)-2:232645896(-)__2_232627501_232652501D;SPAN=41948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:42 GQ:38.3 PL:[38.3, 0.0, 61.4] SR:0 DR:15 LR:-38.14 LO:38.49);ALT=T[chr2:232645896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233271097	+	chr2	233242971	+	.	19	0	1240239_1	49.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1240239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:233242971(-)-2:233271097(+)__2_233240001_233265001D;SPAN=28126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:51 GQ:49.1 PL:[49.1, 0.0, 72.2] SR:0 DR:19 LR:-48.9 LO:49.2);ALT=]chr2:233271097]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	233415486	+	chr2	233421137	+	.	11	0	1240761_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1240761_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:233415486(+)-2:233421137(-)__2_233411501_233436501D;SPAN=5651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:93 GQ:11.3 PL:[11.3, 0.0, 212.6] SR:0 DR:11 LR:-11.12 LO:22.18);ALT=T[chr2:233421137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233415489	+	chr2	233422591	+	.	20	0	1240762_1	38.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1240762_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:233415489(+)-2:233422591(-)__2_233411501_233436501D;SPAN=7102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:102 GQ:38.6 PL:[38.6, 0.0, 206.9] SR:0 DR:20 LR:-38.39 LO:45.13);ALT=C[chr2:233422591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233421241	+	chr2	233428957	+	CTGTTGTCCCTGGACCGGCAGAGCATCCCCTGCAGTACAACTACACTTTTTGGTACTCCAGGAGAACCCCCGGCCGTCCCACGAGCTCACAGAGCTATGAACAGAATATCAAACAGATTGGCACCTTTGCCTCT	0	35	1240784_1	94.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GTG;INSERTION=CTGTTGTCCCTGGACCGGCAGAGCATCCCCTGCAGTACAACTACACTTTTTGGTACTCCAGGAGAACCCCCGGCCGTCCCACGAGCTCACAGAGCTATGAACAGAATATCAAACAGATTGGCACCTTTGCCTCT;MAPQ=60;MATEID=1240784_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_2_233411501_233436501_376C;SPAN=7716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:79 GQ:94.1 PL:[94.1, 0.0, 97.4] SR:35 DR:0 LR:-94.13 LO:94.14);ALT=G[chr2:233428957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233422731	+	chr2	233428957	+	.	0	8	1240791_1	4.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GTG;MAPQ=60;MATEID=1240791_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_2_233411501_233436501_376C;SPAN=6226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:8 DR:0 LR:-4.192 LO:15.42);ALT=G[chr2:233428957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233562154	+	chr2	233599857	+	.	8	0	1241386_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1241386_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:233562154(+)-2:233599857(-)__2_233583001_233608001D;SPAN=37703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:0 DR:8 LR:-16.11 LO:18.33);ALT=G[chr2:233599857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	233677201	+	chr2	233680342	+	.	2	3	1241513_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TACAG;MAPQ=60;MATEID=1241513_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_2_233656501_233681501_272C;SPAN=3141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:85 GQ:6.3 PL:[0.0, 6.3, 217.8] SR:3 DR:2 LR:6.524 LO:8.497);ALT=G[chr2:233680342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124704272	+	chr2	235414066	+	.	5	17	1246105_1	59.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=ATATATATATA;MAPQ=16;MATEID=1246105_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_235396001_235421001_72C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:21 DP:18 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:17 DR:5 LR:-59.41 LO:59.41);ALT=]chr11:124704272]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr2	237994645	+	chr3	68194175	+	.	15	0	1465891_1	36.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1465891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:237994645(+)-3:68194175(-)__3_68183501_68208501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:48 GQ:36.5 PL:[36.5, 0.0, 79.4] SR:0 DR:15 LR:-36.51 LO:37.4);ALT=T[chr3:68194175[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr2	238601165	+	chr2	238617186	+	.	0	33	1254675_1	94.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=1254675_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_238605501_238630501_190C;SPAN=16021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:54 GQ:35 PL:[94.4, 0.0, 35.0] SR:33 DR:0 LR:-95.68 LO:95.68);ALT=G[chr2:238617186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	238601169	+	chr3	178978986	-	.	9	0	1811902_1	11.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1811902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:238601169(+)-3:178978986(+)__3_178972501_178997501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=G]chr3:178978986];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	238875775	+	chr2	238881731	+	.	53	13	1255559_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=1255559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_238875001_238900001_298C;SPAN=5956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:54 GQ:15 PL:[165.0, 15.0, 0.0] SR:13 DR:53 LR:-165.0 LO:165.0);ALT=G[chr2:238881731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	238875793	+	chr20	3276848	-	.	19	0	6893536_1	47.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6893536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:238875793(+)-20:3276848(+)__20_3258501_3283501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:57 GQ:47.3 PL:[47.3, 0.0, 90.2] SR:0 DR:19 LR:-47.28 LO:48.04);ALT=G]chr20:3276848];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr2	238944582	+	chr2	238949927	+	.	0	12	1255792_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1255792_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_238948501_238973501_206C;SPAN=5345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:40 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:12 DR:0 LR:-28.78 LO:29.66);ALT=G[chr2:238949927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	239098616	+	chr2	239112139	+	AATCGCCACTGCTAGCGGGTGGGAGATCATCAAAAAGCAAAGGTCCCCCTGATCCTGAGTCAGTACTGCTGGCCGGAGGGAGGTCATCAAAGAGCAGGGGTCCTTTCTGAGCTTCTTTC	0	24	1256086_1	61.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AATCGCCACTGCTAGCGGGTGGGAGATCATCAAAAAGCAAAGGTCCCCCTGATCCTGAGTCAGTACTGCTGGCCGGAGGGAGGTCATCAAAGAGCAGGGGTCCTTTCTGAGCTTCTTTC;MAPQ=60;MATEID=1256086_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_2_239095501_239120501_152C;SPAN=13523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:65 GQ:61.7 PL:[61.7, 0.0, 94.7] SR:24 DR:0 LR:-61.61 LO:62.03);ALT=G[chr2:239112139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	239103022	+	chr2	239112214	+	.	8	0	1256104_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1256104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:239103022(+)-2:239112214(-)__2_239095501_239120501D;SPAN=9192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:52 GQ:12.5 PL:[12.5, 0.0, 111.5] SR:0 DR:8 LR:-12.32 LO:17.12);ALT=T[chr2:239112214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	239103561	+	chr2	239112234	+	.	15	0	1256108_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1256108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=2:239103561(+)-2:239112234(-)__2_239095501_239120501D;SPAN=8673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:0 DR:15 LR:-35.16 LO:36.62);ALT=A[chr2:239112234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9432182	+	chr3	9433361	+	.	0	10	1280158_1	24.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=1280158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_9408001_9433001_31C;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:31 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:10 DR:0 LR:-24.61 LO:25.11);ALT=C[chr3:9433361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9691428	+	chr3	9695303	+	.	0	16	1280713_1	35.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=1280713_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_9677501_9702501_234C;SPAN=3875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:63 GQ:35.9 PL:[35.9, 0.0, 115.1] SR:16 DR:0 LR:-35.75 LO:38.17);ALT=T[chr3:9695303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9710479	+	chr3	9712731	+	GGGTGCAGATGATGCCTGGGCAGATGTGGAGGACGTCACGGAGGAGGACTGTGCTCTTC	0	7	1280476_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GGGTGCAGATGATGCCTGGGCAGATGTGGAGGACGTCACGGAGGAGGACTGTGCTCTTC;MAPQ=60;MATEID=1280476_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_9702001_9727001_124C;SPAN=2252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:55 GQ:8.3 PL:[8.3, 0.0, 123.8] SR:7 DR:0 LR:-8.206 LO:14.35);ALT=G[chr3:9712731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9834861	+	chr3	9843341	+	.	14	0	1281016_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1281016_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:9834861(+)-3:9843341(-)__3_9824501_9849501D;SPAN=8480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:0 DR:14 LR:-28.06 LO:32.03);ALT=A[chr3:9843341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9834868	+	chr3	9839341	+	.	25	0	1281017_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1281017_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:9834868(+)-3:9839341(-)__3_9824501_9849501D;SPAN=4473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:116 GQ:51.2 PL:[51.2, 0.0, 229.4] SR:0 DR:25 LR:-51.1 LO:57.58);ALT=C[chr3:9839341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9834882	+	chr3	9841864	+	.	57	0	1281018_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1281018_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:9834882(+)-3:9841864(-)__3_9824501_9849501D;SPAN=6982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:90 GQ:54.8 PL:[163.7, 0.0, 54.8] SR:0 DR:57 LR:-166.8 LO:166.8);ALT=G[chr3:9841864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9839462	+	chr3	9843342	+	AGTAGCAAAGAGCTCCTGTTACAACCTGTGACCATCAGCAGGAATGAGAAGGAAAAGGTTCTGATTGAGGGCTCCATCAACTCTGTCCGGGTCAGCATTGCTGTGAAA	15	147	1281027_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=AGTAGCAAAGAGCTCCTGTTACAACCTGTGACCATCAGCAGGAATGAGAAGGAAAAGGTTCTGATTGAGGGCTCCATCAACTCTGTCCGGGTCAGCATTGCTGTGAAA;MAPQ=60;MATEID=1281027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_9824501_9849501_273C;SPAN=3880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:89 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:147 DR:15 LR:-435.7 LO:435.7);ALT=G[chr3:9843342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9839462	+	chr3	9841865	+	.	31	68	1281026_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TCAGG;MAPQ=60;MATEID=1281026_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_3_9824501_9849501_273C;SPAN=2403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:112 GQ:6.2 PL:[263.6, 0.0, 6.2] SR:68 DR:31 LR:-278.0 LO:278.0);ALT=G[chr3:9841865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9841981	+	chr3	9843342	+	.	2	52	1281034_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=1281034_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGATGA;SCTG=c_3_9824501_9849501_273C;SPAN=1361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:85 GQ:34.4 PL:[117.6, 0.0, 34.4] SR:52 DR:2 LR:-120.4 LO:120.4);ALT=G[chr3:9843342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9843441	+	chr3	9845525	+	.	4	18	1281038_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1281038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_9824501_9849501_306C;SPAN=2084;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:60 GQ:53 PL:[53.0, 0.0, 92.6] SR:18 DR:4 LR:-53.07 LO:53.65);ALT=G[chr3:9845525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9845697	+	chr3	9847894	+	.	11	9	1281054_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1281054_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_9824501_9849501_291C;SPAN=2197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:9 DR:11 LR:-39.54 LO:40.27);ALT=T[chr3:9847894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	9932495	+	chr3	9934606	+	TGTGACC	17	10	1281156_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTGACC;MAPQ=60;MATEID=1281156_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_9922501_9947501_158C;SPAN=2111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:68 GQ:50.9 PL:[50.9, 0.0, 113.6] SR:10 DR:17 LR:-50.9 LO:52.23);ALT=G[chr3:9934606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10157503	+	chr3	10167309	+	.	72	83	1281931_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1281931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_10143001_10168001_182C;SPAN=9806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:109 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:83 DR:72 LR:-379.6 LO:379.6);ALT=G[chr3:10167309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10157503	+	chr3	10160589	+	.	4	8	1281930_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1281930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_10143001_10168001_131C;SPAN=3086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:8 DR:4 LR:-9.982 LO:20.14);ALT=G[chr3:10160589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10157541	+	chr3	10167951	+	.	71	0	1281932_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1281932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10157541(+)-3:10167951(-)__3_10143001_10168001D;SPAN=10410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:90 GQ:8.6 PL:[209.9, 0.0, 8.6] SR:0 DR:71 LR:-221.2 LO:221.2);ALT=G[chr3:10167951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10354415	+	chr3	10357005	+	.	0	46	1282485_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1282485_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_10339001_10364001_107C;SPAN=2590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:74 GQ:46.1 PL:[131.9, 0.0, 46.1] SR:46 DR:0 LR:-134.0 LO:134.0);ALT=C[chr3:10357005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10354437	+	chr3	33075435	-	.	8	0	1341593_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1341593_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10354437(+)-3:33075435(+)__3_33075001_33100001D;SPAN=22720998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=G]chr3:33075435];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	10354465	+	chr3	10362729	+	.	32	0	1282488_1	87.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1282488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10354465(+)-3:10362729(-)__3_10339001_10364001D;SPAN=8264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:66 GQ:71.3 PL:[87.8, 0.0, 71.3] SR:0 DR:32 LR:-87.83 LO:87.83);ALT=T[chr3:10362729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10357120	+	chr3	10359734	+	.	2	12	1282490_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1282490_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_10339001_10364001_277C;SPAN=2614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:41 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:12 DR:2 LR:-35.11 LO:35.58);ALT=G[chr3:10359734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	10357149	+	chr3	10362730	+	.	34	0	1282492_1	97.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1282492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:10357149(+)-3:10362730(-)__3_10339001_10364001D;SPAN=5581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:54 GQ:31.7 PL:[97.7, 0.0, 31.7] SR:0 DR:34 LR:-99.33 LO:99.33);ALT=T[chr3:10362730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	11955824	+	chr3	12913431	+	.	12	0	1284848_1	35.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=1284848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:11955824(+)-3:12913431(-)__3_11931501_11956501D;SPAN=957607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:17 GQ:5.3 PL:[35.0, 0.0, 5.3] SR:0 DR:12 LR:-36.15 LO:36.15);ALT=C[chr3:12913431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	12913579	+	chr3	11956085	+	.	13	0	1285034_1	36.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=1285034_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:11956085(-)-3:12913579(+)__3_11956001_11981001D;SPAN=957494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:25 GQ:23 PL:[36.2, 0.0, 23.0] SR:0 DR:13 LR:-36.26 LO:36.26);ALT=]chr3:12913579]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	12369506	-	chr5	139682623	+	.	19	0	2596077_1	52.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2596077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:12369506(-)-5:139682623(-)__5_139674501_139699501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:38 GQ:39.2 PL:[52.4, 0.0, 39.2] SR:0 DR:19 LR:-52.52 LO:52.52);ALT=[chr5:139682623[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	12610502	+	chr3	12611568	+	.	0	5	1286192_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1286192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_12593001_12618001_161C;SPAN=1066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:62 GQ:0 PL:[0.0, 0.0, 148.5] SR:5 DR:0 LR:0.2923 LO:9.206);ALT=G[chr3:12611568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	12881854	+	chr3	12882992	+	.	22	0	1287018_1	46.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=1287018_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:12881854(+)-3:12882992(-)__3_12862501_12887501D;SPAN=1138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:98 GQ:46.1 PL:[46.1, 0.0, 191.3] SR:0 DR:22 LR:-46.07 LO:51.12);ALT=T[chr3:12882992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	13359281	+	chr3	13360572	+	.	3	4	1287652_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1287652_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_13352501_13377501_65C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:64 GQ:2.6 PL:[2.6, 0.0, 151.1] SR:4 DR:3 LR:-2.467 LO:11.46);ALT=T[chr3:13360572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	13455613	+	chr3	13461558	+	.	0	10	1287724_1	16.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=1287724_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_13450501_13475501_42C;SPAN=5945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:10 DR:0 LR:-16.48 LO:21.7);ALT=C[chr3:13461558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	14212053	+	chr3	14214366	+	.	0	8	1289280_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=1289280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_14210001_14235001_155C;SPAN=2313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:8 DR:0 LR:-8.527 LO:16.22);ALT=G[chr3:14214366[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	14214563	+	chr3	14219966	+	.	15	11	1289285_1	51.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1289285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_14210001_14235001_111C;SPAN=5403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:66 GQ:51.5 PL:[51.5, 0.0, 107.6] SR:11 DR:15 LR:-51.44 LO:52.57);ALT=C[chr3:14219966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	14220420	+	chr3	14225434	+	.	12	0	1289298_1	27.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=1289298_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:14220420(+)-3:14225434(-)__3_14210001_14235001D;SPAN=5014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=T[chr3:14225434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	14220424	+	chr3	14239535	+	.	14	0	1289299_1	40.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=1289299_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:14220424(+)-3:14239535(-)__3_14210001_14235001D;SPAN=19111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:20 GQ:7.7 PL:[40.7, 0.0, 7.7] SR:0 DR:14 LR:-42.07 LO:42.07);ALT=C[chr3:14239535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	14693385	+	chr3	14695932	+	.	7	7	1289702_1	22.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1289702_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_14675501_14700501_255C;SPAN=2547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:7 DR:7 LR:-22.49 LO:25.34);ALT=G[chr3:14695932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15094976	+	chr3	15106567	+	AAGTAGAATCGCAGGAAGGGTGACGGCGTCATGTTCTTAAACATCATGATCTGCACCCAAGGGTTTTTGTATTGAATCTGAGGTATGTTGAAAAACACAAACTT	0	57	1290471_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=AAGTAGAATCGCAGGAAGGGTGACGGCGTCATGTTCTTAAACATCATGATCTGCACCCAAGGGTTTTTGTATTGAATCTGAGGTATGTTGAAAAACACAAACTT;MAPQ=60;MATEID=1290471_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_15092001_15117001_41C;SPAN=11591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:72 GQ:3.8 PL:[168.8, 0.0, 3.8] SR:57 DR:0 LR:-177.8 LO:177.8);ALT=T[chr3:15106567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15101032	+	chr3	15106696	+	.	30	0	1290487_1	80.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1290487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:15101032(+)-3:15106696(-)__3_15092001_15117001D;SPAN=5664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:71 GQ:80 PL:[80.0, 0.0, 89.9] SR:0 DR:30 LR:-79.8 LO:79.85);ALT=A[chr3:15106696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15138211	+	chr3	15140573	+	.	11	0	1290438_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1290438_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:15138211(+)-3:15140573(-)__3_15116501_15141501D;SPAN=2362;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=A[chr3:15140573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	6978180	+	chr3	15180686	+	.	12	0	3728710_1	26.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=3728710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:15180686(-)-8:6978180(+)__8_6958001_6983001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:50 GQ:26 PL:[26.0, 0.0, 95.3] SR:0 DR:12 LR:-26.07 LO:28.28);ALT=]chr8:6978180]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	15617606	-	chr16	865370	+	.	2	10	6074006_1	25.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=AGGCTGGAGTGCAGTGGTGTGATCTCGGCTCA;MAPQ=60;MATEID=6074006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_857501_882501_188C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:10 DR:2 LR:-25.75 LO:26.84);ALT=[chr16:865370[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	15712064	+	chr3	15717404	+	.	4	4	1291503_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1291503_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15704501_15729501_263C;SPAN=5340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:50 GQ:6.2 PL:[6.2, 0.0, 115.1] SR:4 DR:4 LR:-6.26 LO:12.14);ALT=C[chr3:15717404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15749573	+	chr3	15751175	+	.	3	3	1291691_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1291691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15729001_15754001_52C;SPAN=1602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:3 DR:3 LR:6.844 LO:6.647);ALT=T[chr3:15751175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15836813	+	chr3	15838556	+	.	2	3	1291978_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1291978_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15827001_15852001_158C;SPAN=1743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:138 GQ:20.7 PL:[0.0, 20.7, 376.2] SR:3 DR:2 LR:20.88 LO:7.427);ALT=G[chr3:15838556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15836814	+	chr3	15837912	+	.	8	15	1291979_1	45.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1291979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15827001_15852001_28C;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:87 GQ:45.8 PL:[45.8, 0.0, 164.6] SR:15 DR:8 LR:-45.75 LO:49.56);ALT=C[chr3:15837912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	15836814	+	chr3	15839478	+	.	9	5	1291980_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1291980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_15827001_15852001_119C;SPAN=2664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:13 DP:165 GQ:1.6 PL:[0.0, 1.6, 402.6] SR:5 DR:9 LR:1.79 LO:23.8);ALT=C[chr3:15839478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	16302338	+	chr3	16306275	+	.	11	5	1292572_1	27.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1292572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_16292501_16317501_128C;SPAN=3937;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:56 GQ:27.8 PL:[27.8, 0.0, 107.0] SR:5 DR:11 LR:-27.74 LO:30.42);ALT=T[chr3:16306275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	16535385	+	chr3	16554949	+	.	9	10	1292950_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1292950_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_16537501_16562501_57C;SPAN=19564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:17 GQ:2 PL:[38.3, 0.0, 2.0] SR:10 DR:9 LR:-40.1 LO:40.1);ALT=C[chr3:16554949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	17914057	+	chr10	71993020	+	.	53	14	1294793_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=TGAGGAAGACTCGGTACTCCAGGGAGAAGGG;MAPQ=42;MATEID=1294793_2;MATENM=0;NM=9;NUMPARTS=2;SCTG=c_3_17909501_17934501_217C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:32 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:14 DR:53 LR:-188.1 LO:188.1);ALT=G[chr10:71993020[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	18419819	+	chr3	18427888	+	.	5	5	1295442_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=1295442_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_18399501_18424501_92C;SPAN=8069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:5 DR:5 LR:-20.77 LO:21.8);ALT=T[chr3:18427888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	23244754	+	chr3	23250182	+	.	0	19	1301601_1	46.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=1301601_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_23226001_23251001_129C;SPAN=5428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:62 GQ:46.1 PL:[46.1, 0.0, 102.2] SR:19 DR:0 LR:-45.92 LO:47.18);ALT=G[chr3:23250182[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	23847580	+	chr3	23848726	+	.	41	4	1302368_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1302368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_23838501_23863501_262C;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:41 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:4 DR:41 LR:-125.4 LO:125.4);ALT=G[chr3:23848726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	23848912	+	chr3	23929055	+	AATTCAGAAGGAGCTGGCGGACATCACTTTAGACCCTCCACCTAATTG	3	22	1302374_1	82.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AATTCAGAAGGAGCTGGCGGACATCACTTTAGACCCTCCACCTAATTG;MAPQ=60;MATEID=1302374_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_23838501_23863501_230C;SPAN=80143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:22 DR:3 LR:-82.01 LO:82.01);ALT=G[chr3:23929055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	23848912	+	chr3	23852949	+	.	2	19	1302373_1	51.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=1302373_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_3_23838501_23863501_230C;SPAN=4037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:53 GQ:51.8 PL:[51.8, 0.0, 74.9] SR:19 DR:2 LR:-51.66 LO:51.93);ALT=G[chr3:23852949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	29831222	+	chr3	23971993	+	.	8	0	3230680_1	18.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3230680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:23971993(-)-7:29831222(+)__7_29816501_29841501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:0 DR:8 LR:-18.55 LO:19.42);ALT=]chr7:29831222]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	31624726	+	chr3	31627038	-	.	2	3	1335604_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCAAT;MAPQ=60;MATEID=1335604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_31605001_31630001_365C;SPAN=2312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:101 GQ:13.8 PL:[0.0, 13.8, 270.6] SR:3 DR:2 LR:14.16 LO:6.098);ALT=T]chr3:31627038];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	31670903	+	chr3	31674422	+	.	4	3	1335775_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGCAG;MAPQ=60;MATEID=1335775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_31654001_31679001_159C;SPAN=3519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:83 GQ:5.7 PL:[0.0, 5.7, 211.2] SR:3 DR:4 LR:5.982 LO:8.55);ALT=G[chr3:31674422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32102052	+	chr3	32107884	+	.	0	99	1337455_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1337455_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_32095001_32120001_84C;SPAN=5832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:54 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:99 DR:0 LR:-293.8 LO:293.8);ALT=C[chr3:32107884[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32163315	+	chr22	21309767	+	.	9	0	7224165_1	26.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=7224165_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:32163315(+)-22:21309767(-)__22_21290501_21315501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:9 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=T[chr22:21309767[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	32433557	+	chr3	32444523	+	.	0	10	1338863_1	17.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1338863_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32438001_32463001_376C;SPAN=10966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:10 DR:0 LR:-17.57 LO:22.03);ALT=G[chr3:32444523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32433559	+	chr3	32483331	+	.	31	38	1338760_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1338760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32462501_32487501_398C;SPAN=49772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:67 GQ:8.3 PL:[153.5, 0.0, 8.3] SR:38 DR:31 LR:-161.2 LO:161.2);ALT=T[chr3:32483331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32529529	+	chr3	32533201	+	.	3	4	1339013_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1339013_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32511501_32536501_372C;SPAN=3672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:98 GQ:9.9 PL:[0.0, 9.9, 257.4] SR:4 DR:3 LR:10.05 LO:8.181);ALT=C[chr3:32533201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32533379	+	chr3	32544100	+	.	30	36	1339260_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1339260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32536001_32561001_85C;SPAN=10721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:75 GQ:26 PL:[154.7, 0.0, 26.0] SR:36 DR:30 LR:-159.7 LO:159.7);ALT=C[chr3:32544100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32568402	+	chr3	32569937	+	.	0	11	1339189_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1339189_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32560501_32585501_274C;SPAN=1535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:106 GQ:7.7 PL:[7.7, 0.0, 248.6] SR:11 DR:0 LR:-7.593 LO:21.52);ALT=T[chr3:32569937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32587458	+	chr3	32612115	+	CAGCAGTAGCACGTTCTTCCCCGCAGGGAGCTTGGAGCGCGAGCGGGTGGAGACCTCGCTGAGGATGCAGG	6	30	1339486_1	91.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=CAGCAGTAGCACGTTCTTCCCCGCAGGGAGCTTGGAGCGCGAGCGGGTGGAGACCTCGCTGAGGATGCAGG;MAPQ=60;MATEID=1339486_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_32609501_32634501_201C;SPAN=24657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:54 GQ:38.3 PL:[91.1, 0.0, 38.3] SR:30 DR:6 LR:-92.08 LO:92.08);ALT=C[chr3:32612115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32716395	-	chr7	32117278	+	.	13	47	1340470_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GGTTCAAGC;MAPQ=51;MATEID=1340470_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_3_32707501_32732501_345C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:42 GQ:15 PL:[165.0, 15.0, 0.0] SR:47 DR:13 LR:-165.0 LO:165.0);ALT=[chr7:32117278[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	32726974	+	chr3	32745355	+	.	0	7	1340530_1	9.0	.	EVDNC=ASSMB;HOMSEQ=TGCAG;MAPQ=60;MATEID=1340530_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_32707501_32732501_430C;SPAN=18381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=G[chr3:32745355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	32806763	+	chr3	32808062	+	.	50	18	1340216_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=TTGCAGTGAGCCAAGAT;MAPQ=60;MATEID=1340216_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_32805501_32830501_315C;SPAN=1299;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:78 GQ:15.2 PL:[173.6, 0.0, 15.2] SR:18 DR:50 LR:-181.4 LO:181.4);ALT=T[chr3:32808062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	33114235	+	chr3	33138540	+	.	17	0	1341933_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1341933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:33114235(+)-3:33138540(-)__3_33124001_33149001D;SPAN=24305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:40 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:0 DR:17 LR:-45.28 LO:45.31);ALT=A[chr3:33138540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	33175758	+	chr3	33183885	+	.	3	5	1342145_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1342145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_33173001_33198001_255C;SPAN=8127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:93 GQ:5.1 PL:[0.0, 5.1, 234.3] SR:5 DR:3 LR:5.39 LO:10.44);ALT=G[chr3:33183885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	37019918	+	chr3	37020968	-	.	8	0	1353919_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1353919_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:37019918(+)-3:37020968(+)__3_37019501_37044501D;SPAN=1050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:120 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.103 LO:14.04);ALT=C]chr3:37020968];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	37133030	+	chr3	37136282	+	.	0	7	1354356_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1354356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37117501_37142501_79C;SPAN=3252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:107 GQ:5.7 PL:[0.0, 5.7, 270.6] SR:7 DR:0 LR:5.882 LO:12.23);ALT=C[chr3:37136282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	37190531	+	chr3	37216029	+	.	0	8	1354778_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1354778_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37166501_37191501_300C;SPAN=25498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:8 DR:0 LR:-13.67 LO:17.51);ALT=T[chr3:37216029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	37216099	+	chr3	37217551	+	.	0	28	1354886_1	65.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=1354886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37215501_37240501_280C;SPAN=1452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:101 GQ:65.3 PL:[65.3, 0.0, 177.5] SR:28 DR:0 LR:-65.07 LO:68.06);ALT=G[chr3:37217551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	37449928	+	chr3	39676077	-	.	36	42	1356067_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGTGAGCCAAGATCATGCCACTACACTCCAGCCTG;MAPQ=60;MATEID=1356067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37436001_37461001_212C;SPAN=2226149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:44 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:42 DR:36 LR:-221.2 LO:221.2);ALT=G]chr3:39676077];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	37450057	-	chr3	39675868	+	.	46	0	1356068_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=1356068_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:37450057(-)-3:39675868(-)__3_37436001_37461001D;SPAN=2225811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:60 GQ:10.1 PL:[135.5, 0.0, 10.1] SR:0 DR:46 LR:-142.0 LO:142.0);ALT=[chr3:39675868[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	37876187	-	chr3	37877290	+	.	3	3	1357327_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1357327_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_37877001_37902001_40C;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:54 GQ:1.2 PL:[0.0, 1.2, 132.0] SR:3 DR:3 LR:1.426 LO:7.211);ALT=[chr3:37877290[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	38164615	+	chr3	38167055	+	.	2	2	1357970_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1357970_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_38146501_38171501_86C;SPAN=2440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:110 GQ:16.5 PL:[0.0, 16.5, 300.3] SR:2 DR:2 LR:16.6 LO:5.948);ALT=T[chr3:38167055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	38173498	+	chr3	38178082	+	CAGAAACTGGGCGATTCGGGCCATGATTGCCCCGGCCCCAGGCTGCAGCACATTT	0	11	1358101_1	0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CAGAAACTGGGCGATTCGGGCCATGATTGCCCCGGCCCCAGGCTGCAGCACATTT;MAPQ=60;MATEID=1358101_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_38171001_38196001_222C;SPAN=4584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:135 GQ:0 PL:[0.0, 0.0, 326.7] SR:11 DR:0 LR:0.2638 LO:20.3);ALT=T[chr3:38178082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	38627164	+	chr3	149162142	-	.	7	83	1360381_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GATGGTGTGTGTGTG;MAPQ=60;MATEID=1360381_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_38612001_38637001_360C;SPAN=110534978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:93 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:83 DR:7 LR:-274.0 LO:274.0);ALT=G]chr3:149162142];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	39188216	+	chr3	39194928	+	.	0	10	1361867_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=1361867_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_39175501_39200501_258C;SPAN=6712;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:10 DR:0 LR:-4.834 LO:19.21);ALT=G[chr3:39194928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	40498968	+	chr12	63359104	+	.	92	9	5220782_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5220782_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_63357001_63382001_5C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:101 DP:1279 GQ:12.8 PL:[0.0, 12.8, 3132.0] SR:9 DR:92 LR:13.11 LO:185.0);ALT=G[chr12:63359104[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	41818076	+	chr3	41821494	+	.	43	24	1370814_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAGGTACAAAATG;MAPQ=60;MATEID=1370814_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_41821501_41846501_79C;SPAN=3418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:27 GQ:15 PL:[165.0, 15.0, 0.0] SR:24 DR:43 LR:-165.0 LO:165.0);ALT=G[chr3:41821494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	41996326	+	chr3	42003503	+	.	14	0	1371558_1	20.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1371558_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:41996326(+)-3:42003503(-)__3_41993001_42018001D;SPAN=7177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:95 GQ:20.6 PL:[20.6, 0.0, 208.7] SR:0 DR:14 LR:-20.48 LO:29.67);ALT=A[chr3:42003503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42610600	+	chr3	42623389	+	.	11	0	1373872_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1373872_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:42610600(+)-3:42623389(-)__3_42605501_42630501D;SPAN=12789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:0 DR:11 LR:-7.051 LO:21.42);ALT=C[chr3:42623389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42633146	+	chr3	42635913	+	.	40	0	1374140_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1374140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:42633146(+)-3:42635913(-)__3_42630001_42655001D;SPAN=2767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:110 GQ:99 PL:[102.2, 0.0, 164.9] SR:0 DR:40 LR:-102.2 LO:103.0);ALT=G[chr3:42635913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	35164256	+	chr3	42635913	+	.	12	0	4571479_1	31.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4571479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:42635913(-)-10:35164256(+)__10_35157501_35182501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:30 GQ:31.4 PL:[31.4, 0.0, 41.3] SR:0 DR:12 LR:-31.48 LO:31.56);ALT=]chr10:35164256]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	42659137	+	chr3	42660509	+	.	0	9	1374261_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=1374261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_42654501_42679501_266C;SPAN=1372;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:9 DR:0 LR:-3.429 LO:17.14);ALT=G[chr3:42660509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42676860	+	chr3	42678360	+	.	0	8	1374316_1	0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=1374316_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_42654501_42679501_191C;SPAN=1500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:8 DR:0 LR:3.394 LO:14.36);ALT=T[chr3:42678360[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	42838373	+	chr3	42840811	+	.	107	53	1374684_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGAATCTTATAACTTCC;MAPQ=60;MATEID=1374684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_42826001_42851001_299C;SPAN=2438;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:40 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:53 DR:107 LR:-452.2 LO:452.2);ALT=C[chr3:42840811[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	43586022	-	chr3	43587026	+	.	8	0	1377277_1	0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1377277_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:43586022(-)-3:43587026(-)__3_43585501_43610501D;SPAN=1004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:123 GQ:6.6 PL:[0.0, 6.6, 310.2] SR:0 DR:8 LR:6.916 LO:13.95);ALT=[chr3:43587026[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	43732533	+	chr3	43740766	+	.	6	4	1377576_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1377576_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_43732501_43757501_386C;SPAN=8233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:4 DR:6 LR:-3.971 LO:17.23);ALT=T[chr3:43740766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	44380346	+	chr3	44399230	+	.	8	0	1379796_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1379796_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:44380346(+)-3:44399230(-)__3_44394001_44419001D;SPAN=18884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=G[chr3:44399230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	44548451	+	chr3	44552040	+	.	26	0	1380505_1	52.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1380505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:44548451(+)-3:44552040(-)__3_44541001_44566001D;SPAN=3589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:124 GQ:52.4 PL:[52.4, 0.0, 247.1] SR:0 DR:26 LR:-52.23 LO:59.53);ALT=C[chr3:44552040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	44740991	-	chr3	44742263	+	.	78	81	1381228_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCACTTTGGGA;MAPQ=60;MATEID=1381228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_251C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:101 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:81 DR:78 LR:-429.1 LO:429.1);ALT=[chr3:44742263[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	44741013	+	chr3	44742285	-	.	61	63	1381229_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TCCCAAAGTGCTGGGATTACAGG;MAPQ=60;MATEID=1381229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44737001_44762001_127C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:105 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:63 DR:61 LR:-326.8 LO:326.8);ALT=A]chr3:44742285];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	45000953	+	chr3	45017425	+	.	0	9	1382048_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1382048_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_44982001_45007001_332C;SPAN=16472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:9 DR:0 LR:-14.54 LO:19.45);ALT=C[chr3:45017425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	45017842	+	chr3	45030630	+	.	10	0	1381938_1	4.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1381938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:45017842(+)-3:45030630(-)__3_45006501_45031501D;SPAN=12788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:0 DR:10 LR:-4.292 LO:19.12);ALT=G[chr3:45030630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	45017842	+	chr3	45031039	+	.	16	0	1382069_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1382069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:45017842(+)-3:45031039(-)__3_45031001_45056001D;SPAN=13197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:58 GQ:37.1 PL:[37.1, 0.0, 103.1] SR:0 DR:16 LR:-37.1 LO:38.85);ALT=G[chr3:45031039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	45031136	+	chr3	45038578	+	.	0	10	1382072_1	1.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1382072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_45031001_45056001_94C;SPAN=7442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:116 GQ:1.7 PL:[1.7, 0.0, 278.9] SR:10 DR:0 LR:-1.583 LO:18.71);ALT=G[chr3:45038578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	45049067	+	chr3	45052725	+	.	0	7	1382126_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1382126_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_45031001_45056001_250C;SPAN=3658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:126 GQ:10.8 PL:[0.0, 10.8, 326.7] SR:7 DR:0 LR:11.03 LO:11.72);ALT=G[chr3:45052725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	33049630	+	chr3	46610892	+	.	0	10	1387672_1	18.0	.	EVDNC=ASSMB;HOMSEQ=TTCCA;MAPQ=60;MATEID=1387672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_46599001_46624001_152C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:10 DR:0 LR:-18.11 LO:22.2);ALT=]chr15:33049630]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	46963803	+	chr3	46966946	+	AGTCAGGCTTCCGAGGAGCGAGGTTGGCCAGGTCCACCTCCTCGATGACGGGCTCGGGCTTGGCGGCCTCCAGCTGCTCCTTCACCTTCTCCTCCA	0	21	1389122_1	42.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AGTCAGGCTTCCGAGGAGCGAGGTTGGCCAGGTCCACCTCCTCGATGACGGGCTCGGGCTTGGCGGCCTCCAGCTGCTCCTTCACCTTCTCCTCCA;MAPQ=60;MATEID=1389122_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_46942001_46967001_405C;SPAN=3143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:101 GQ:42.2 PL:[42.2, 0.0, 200.6] SR:21 DR:0 LR:-41.96 LO:47.99);ALT=C[chr3:46966946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	46967028	+	chr3	47018126	+	TGCTTCTCGCCTTCTTCCTCCTCTTCTCTGAGATGCTTGGTCTTTGGCTCCCCATCTTCCTTGT	12	18	1389329_1	60.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TGCTTCTCGCCTTCTTCCTCCTCTTCTCTGAGATGCTTGGTCTTTGGCTCCCCATCTTCCTTGT;MAPQ=60;MATEID=1389329_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_47015501_47040501_310C;SPAN=51098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:71 GQ:60.2 PL:[60.2, 0.0, 109.7] SR:18 DR:12 LR:-59.99 LO:60.86);ALT=G[chr3:47018126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	46982557	+	chr3	47018126	+	.	6	4	1389330_1	4.0	.	DISC_MAPQ=48;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1389330_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GCGC;SCTG=c_3_47015501_47040501_310C;SPAN=35569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:71 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:4 DR:6 LR:-3.871 LO:13.53);ALT=T[chr3:47018126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47166040	+	chr3	47205344	+	CATTTTCTTCTTCT	5	3	1389932_1	11.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=CATTTTCTTCTTCT;MAPQ=60;MATEID=1389932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47187001_47212001_67C;SPAN=39304;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:32 GQ:11.3 PL:[11.3, 0.0, 64.1] SR:3 DR:5 LR:-11.14 LO:13.41);ALT=T[chr3:47205344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47206088	+	chr3	47210657	+	.	3	2	1390013_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1390013_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47187001_47212001_194C;SPAN=4569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:93 GQ:11.7 PL:[0.0, 11.7, 247.5] SR:2 DR:3 LR:11.99 LO:6.243);ALT=G[chr3:47210657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47316980	+	chr3	47318772	+	.	0	8	1390197_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1390197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47309501_47334501_93C;SPAN=1792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:8 DR:0 LR:-0.9411 LO:14.92);ALT=T[chr3:47318772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47324525	+	chr3	47328707	+	.	9	0	1390235_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1390235_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:47324525(+)-3:47328707(-)__3_47309501_47334501D;SPAN=4182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:0 DR:9 LR:-2.075 LO:16.94);ALT=G[chr3:47328707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47490669	+	chr3	47493441	+	.	78	40	1391327_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=1391327_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47481001_47506001_157C;SPAN=2772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:73 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:40 DR:78 LR:-283.9 LO:283.9);ALT=C[chr3:47493441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47551794	+	chr3	47555108	+	.	8	0	1392072_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1392072_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:47551794(+)-3:47555108(-)__3_47530001_47555001D;SPAN=3314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:52 GQ:12.5 PL:[12.5, 0.0, 111.5] SR:0 DR:8 LR:-12.32 LO:17.12);ALT=C[chr3:47555108[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47552718	+	chr3	47555026	+	.	0	11	1392078_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1392078_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_47530001_47555001_113C;SPAN=2308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:105 GQ:8 PL:[8.0, 0.0, 245.6] SR:11 DR:0 LR:-7.864 LO:21.56);ALT=T[chr3:47555026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47742893	+	chr3	47747899	+	.	4	8	1392721_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1392721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47726001_47751001_338C;SPAN=5006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:104 GQ:8.3 PL:[8.3, 0.0, 242.6] SR:8 DR:4 LR:-8.135 LO:21.61);ALT=C[chr3:47747899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47748022	+	chr3	47752173	+	.	2	5	1392747_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1392747_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_47726001_47751001_183C;SPAN=4151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:66 GQ:2 PL:[2.0, 0.0, 157.1] SR:5 DR:2 LR:-1.925 LO:11.37);ALT=T[chr3:47752173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	47844744	+	chr3	47852116	+	.	9	0	1393301_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1393301_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:47844744(+)-3:47852116(-)__3_47824001_47849001D;SPAN=7372;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:52 GQ:15.8 PL:[15.8, 0.0, 108.2] SR:0 DR:9 LR:-15.62 LO:19.77);ALT=G[chr3:47852116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48040413	+	chr3	48130267	+	.	22	0	1394287_1	61.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1394287_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48040413(+)-3:48130267(-)__3_48118001_48143001D;SPAN=89854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:41 GQ:35.3 PL:[61.7, 0.0, 35.3] SR:0 DR:22 LR:-61.81 LO:61.81);ALT=A[chr3:48130267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48155423	-	chr3	48156847	+	.	8	0	1394742_1	1.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=1394742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48155423(-)-3:48156847(-)__3_48142501_48167501D;SPAN=1424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=[chr3:48156847[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	48223008	-	chr14	92587989	+	.	9	0	5844808_1	5.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=5844808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48223008(-)-14:92587989(-)__14_92585501_92610501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.326 LO:17.45);ALT=[chr14:92587989[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	48338321	+	chr3	48339916	+	.	0	7	1395245_1	7.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1395245_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_48338501_48363501_321C;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:58 GQ:7.4 PL:[7.4, 0.0, 132.8] SR:7 DR:0 LR:-7.393 LO:14.18);ALT=T[chr3:48339916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48338356	+	chr3	48342797	+	.	8	0	1395246_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1395246_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48338356(+)-3:48342797(-)__3_48338501_48363501D;SPAN=4441;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=G[chr3:48342797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48511243	+	chr3	48514417	+	.	53	10	1396355_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=28;MATEID=1396355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48510001_48535001_18C;SPAN=3174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:130 GQ:99 PL:[162.8, 0.0, 152.9] SR:10 DR:53 LR:-162.9 LO:162.9);ALT=C[chr3:48514417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48642258	+	chr3	48647003	+	.	15	0	1396657_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1396657_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48642258(+)-3:48647003(-)__3_48632501_48657501D;SPAN=4745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:116 GQ:18.2 PL:[18.2, 0.0, 262.4] SR:0 DR:15 LR:-18.09 LO:30.87);ALT=C[chr3:48647003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48643290	+	chr3	48646592	+	.	3	97	1396661_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=1396661_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48632501_48657501_442C;SPAN=3302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:164 GQ:99 PL:[285.8, 0.0, 110.9] SR:97 DR:3 LR:-289.8 LO:289.8);ALT=C[chr3:48646592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48643336	+	chr3	48647003	+	.	63	0	1396662_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1396662_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48643336(+)-3:48647003(-)__3_48632501_48657501D;SPAN=3667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:107 GQ:80 PL:[179.0, 0.0, 80.0] SR:0 DR:63 LR:-181.0 LO:181.0);ALT=G[chr3:48647003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48732895	+	chr3	48754588	+	.	22	0	1397076_1	34.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1397076_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48732895(+)-3:48754588(-)__3_48730501_48755501D;SPAN=21693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:143 GQ:34.1 PL:[34.1, 0.0, 311.3] SR:0 DR:22 LR:-33.88 LO:47.08);ALT=C[chr3:48754588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48929507	+	chr3	48936121	+	.	0	10	1398219_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=1398219_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48926501_48951501_7C;SPAN=6614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:124 GQ:0.3 PL:[0.0, 0.3, 300.3] SR:10 DR:0 LR:0.5846 LO:18.41);ALT=T[chr3:48936121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48956401	+	chr3	48964892	+	.	13	0	1398087_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1398087_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:48956401(+)-3:48964892(-)__3_48951001_48976001D;SPAN=8491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:115 GQ:11.9 PL:[11.9, 0.0, 266.0] SR:0 DR:13 LR:-11.76 LO:25.94);ALT=G[chr3:48964892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48956431	+	chr3	48960180	+	.	10	14	1398088_1	37.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1398088_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48951001_48976001_348C;SPAN=3749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:81 GQ:37.7 PL:[37.7, 0.0, 156.5] SR:14 DR:10 LR:-37.47 LO:41.73);ALT=G[chr3:48960180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48956431	+	chr3	48962150	+	.	17	3	1398089_1	31.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1398089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48951001_48976001_115C;SPAN=5719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:93 GQ:31.1 PL:[31.1, 0.0, 192.8] SR:3 DR:17 LR:-30.92 LO:37.78);ALT=G[chr3:48962150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48960244	+	chr3	48962148	+	.	0	12	1398111_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1398111_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48951001_48976001_164C;SPAN=1904;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:94 GQ:14.3 PL:[14.3, 0.0, 212.3] SR:12 DR:0 LR:-14.15 LO:24.62);ALT=G[chr3:48962148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48960244	+	chr3	48964893	+	.	0	10	1398112_1	3.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1398112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48951001_48976001_338C;SPAN=4649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:108 GQ:3.8 PL:[3.8, 0.0, 257.9] SR:10 DR:0 LR:-3.75 LO:19.04);ALT=G[chr3:48964893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	48962272	+	chr3	48964893	+	.	0	10	1398132_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1398132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_48951001_48976001_397C;SPAN=2621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:107 GQ:4.1 PL:[4.1, 0.0, 254.9] SR:10 DR:0 LR:-4.021 LO:19.08);ALT=G[chr3:48964893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49058004	+	chr3	49059779	+	.	13	7	1398613_1	31.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1398613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49049001_49074001_322C;SPAN=1775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:81 GQ:31.1 PL:[31.1, 0.0, 163.1] SR:7 DR:13 LR:-30.87 LO:36.16);ALT=G[chr3:49059779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49133514	+	chr3	49135425	+	.	0	45	1399420_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1399420_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49122501_49147501_108C;SPAN=1911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:124 GQ:99 PL:[115.1, 0.0, 184.4] SR:45 DR:0 LR:-115.0 LO:115.9);ALT=T[chr3:49135425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49365251	+	chr3	49372902	+	.	0	13	1400240_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1400240_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49367501_49392501_239C;SPAN=7651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:13 DR:0 LR:-28.55 LO:30.78);ALT=T[chr3:49372902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49365293	+	chr3	49377400	+	.	11	0	1400241_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1400241_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:49365293(+)-3:49377400(-)__3_49367501_49392501D;SPAN=12107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=G[chr3:49377400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49373030	+	chr3	49377355	+	.	22	7	1400280_1	49.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1400280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49367501_49392501_312C;SPAN=4325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:109 GQ:49.7 PL:[49.7, 0.0, 214.7] SR:7 DR:22 LR:-49.69 LO:55.53);ALT=C[chr3:49377355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49397817	+	chr3	49399928	+	.	33	46	1400882_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1400882_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_49392001_49417001_2C;SPAN=2111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:120 GQ:89.6 PL:[201.8, 0.0, 89.6] SR:46 DR:33 LR:-204.2 LO:204.2);ALT=T[chr3:49399928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49397817	+	chr3	49412865	+	GCTTCATCTTGGCTAGCTCCCGCCTTGTGTGCTCATCATTCCGAAGATCCTTCTTATTCCCAACCAGGATGATGGGCACGTTGGGACAGAAATGCTTGACTTCTGGGGTCCACTTTTCTGGGATGTTTTCTAAACTATCAGGGCTGTCGATGGAAAAACACATCAGTATAACATCGGTATCTGGGTAGGAGAGGGGCCTCAGGCGATCATAATCTTCCTGCCCAGCTGTGTCCCACAAAGCCAACTCT	0	144	1400883_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=GCTTCATCTTGGCTAGCTCCCGCCTTGTGTGCTCATCATTCCGAAGATCCTTCTTATTCCCAACCAGGATGATGGGCACGTTGGGACAGAAATGCTTGACTTCTGGGGTCCACTTTTCTGGGATGTTTTCTAAACTATCAGGGCTGTCGATGGAAAAACACATCAGTATAACATCGGTATCTGGGTAGGAGAGGGGCCTCAGGCGATCATAATCTTCCTGCCCAGCTGTGTCCCACAAAGCCAACTCT;MAPQ=60;MATEID=1400883_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_49392001_49417001_2C;SPAN=15048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:144 DP:203 GQ:70.6 PL:[420.5, 0.0, 70.6] SR:144 DR:0 LR:-434.4 LO:434.4);ALT=T[chr3:49412865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49397862	+	chr3	49405859	+	.	26	0	1400885_1	56.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1400885_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:49397862(+)-3:49405859(-)__3_49392001_49417001D;SPAN=7997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:111 GQ:56 PL:[56.0, 0.0, 211.1] SR:0 DR:26 LR:-55.75 LO:60.96);ALT=C[chr3:49405859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49400061	+	chr3	49405861	+	.	27	18	1400901_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1400901_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AA;SCTG=c_3_49392001_49417001_2C;SPAN=5800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:120 GQ:99 PL:[99.5, 0.0, 191.9] SR:18 DR:27 LR:-99.53 LO:101.1);ALT=T[chr3:49405861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49400105	+	chr3	49412864	+	.	13	0	1400903_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=1400903_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:49400105(+)-3:49412864(-)__3_49392001_49417001D;SPAN=12759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:13 DP:177 GQ:4.9 PL:[0.0, 4.9, 439.0] SR:0 DR:13 LR:5.041 LO:23.39);ALT=T[chr3:49412864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49405984	+	chr3	49412865	+	.	0	94	1400942_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=ACCTG;MAPQ=60;MATEID=1400942_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TTT;SCTG=c_3_49392001_49417001_2C;SPAN=6881;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:224 GQ:99 PL:[249.8, 0.0, 292.7] SR:94 DR:0 LR:-249.6 LO:249.8);ALT=G[chr3:49412865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49413026	+	chr3	49449253	+	.	134	51	1400982_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1400982_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_49392001_49417001_476C;SPAN=36227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:142 DP:181 GQ:17.2 PL:[419.9, 0.0, 17.2] SR:51 DR:134 LR:-441.6 LO:441.6);ALT=T[chr3:49449253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	49712054	+	chr3	49713127	+	AGTGGACCCAGAGGGACCTGGAACGCATGGAGAACATTCGATTCTGCCGCCAATACCTGGTGTTCCATGACGGGGACTCAGTGGTGTTTGCAGGACCTGCAGGCAACAGTGTGGAGACCCGGGGGGA	5	25	1402123_1	61.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AGTGGACCCAGAGGGACCTGGAACGCATGGAGAACATTCGATTCTGCCGCCAATACCTGGTGTTCCATGACGGGGACTCAGTGGTGTTTGCAGGACCTGCAGGCAACAGTGTGGAGACCCGGGGGGA;MAPQ=60;MATEID=1402123_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_49710501_49735501_263C;SPAN=1073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:78 GQ:61.4 PL:[61.4, 0.0, 127.4] SR:25 DR:5 LR:-61.39 LO:62.68);ALT=G[chr3:49713127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50107985	+	chr3	50112631	+	.	2	3	1404129_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1404129_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50102501_50127501_86C;SPAN=4646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:85 GQ:6.3 PL:[0.0, 6.3, 217.8] SR:3 DR:2 LR:6.524 LO:8.497);ALT=G[chr3:50112631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50273741	+	chr3	50289530	+	.	10	0	1404474_1	16.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1404474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:50273741(+)-3:50289530(-)__3_50274001_50299001D;SPAN=15789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:63 GQ:16.1 PL:[16.1, 0.0, 134.9] SR:0 DR:10 LR:-15.94 LO:21.55);ALT=G[chr3:50289530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50273888	+	chr3	50289829	+	CTGGGGAGTCAGGGAAGAGCACCATCGTCAAGCAGATGAA	15	38	1404476_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTGGGGAGTCAGGGAAGAGCACCATCGTCAAGCAGATGAA;MAPQ=60;MATEID=1404476_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_50274001_50299001_278C;SPAN=15941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:51 GQ:10.2 PL:[141.9, 10.2, 0.0] SR:38 DR:15 LR:-141.8 LO:141.8);ALT=G[chr3:50289829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50289971	+	chr3	50293624	+	ACGACGCCAGGCAGCTATTTGCACTGTCCTGCACCGCCGAGGAGCAAGGCGTGCTCCCTGATGACCTGTCCGGCGTCATCCGGAGGCTCTGGGCTGACCATGGTGTGCAGGCCTGCTTTGGCCGCTCAAGGGAATACCAGCTCAACGACTCAGCTGCCTA	3	19	1404520_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ACGACGCCAGGCAGCTATTTGCACTGTCCTGCACCGCCGAGGAGCAAGGCGTGCTCCCTGATGACCTGTCCGGCGTCATCCGGAGGCTCTGGGCTGACCATGGTGTGCAGGCCTGCTTTGGCCGCTCAAGGGAATACCAGCTCAACGACTCAGCTGCCTA;MAPQ=60;MATEID=1404520_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_50274001_50299001_50C;SPAN=3653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:91 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:19 DR:3 LR:-38.07 LO:43.46);ALT=G[chr3:50293624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50290616	+	chr3	50293624	+	.	11	11	1404523_1	39.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=1404523_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_50274001_50299001_50C;SPAN=3008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:86 GQ:39.5 PL:[39.5, 0.0, 168.2] SR:11 DR:11 LR:-39.42 LO:43.99);ALT=A[chr3:50293624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50328112	+	chr3	50329645	+	.	18	16	1404891_1	58.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=1404891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50323001_50348001_345C;SPAN=1533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:115 GQ:58.1 PL:[58.1, 0.0, 219.8] SR:16 DR:18 LR:-57.97 LO:63.34);ALT=T[chr3:50329645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50363909	+	chr3	50365385	+	.	0	11	1405024_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1405024_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50347501_50372501_170C;SPAN=1476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:114 GQ:5.6 PL:[5.6, 0.0, 269.6] SR:11 DR:0 LR:-5.426 LO:21.15);ALT=C[chr3:50365385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50369586	+	chr3	50375335	+	.	4	7	1405047_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1405047_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50347501_50372501_353C;SPAN=5749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:7 DR:4 LR:-21.63 LO:23.53);ALT=C[chr3:50375335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50375442	+	chr3	50377987	+	.	0	11	1404643_1	9.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1404643_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50372001_50397001_204C;SPAN=2545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:98 GQ:9.8 PL:[9.8, 0.0, 227.6] SR:11 DR:0 LR:-9.76 LO:21.91);ALT=T[chr3:50377987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50375492	+	chr3	50378198	+	.	8	0	1404644_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1404644_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:50375492(+)-3:50378198(-)__3_50372001_50397001D;SPAN=2706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=G[chr3:50378198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50646025	+	chr3	50649062	+	.	15	5	1405846_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1405846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50641501_50666501_65C;SPAN=3037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:106 GQ:27.5 PL:[27.5, 0.0, 228.8] SR:5 DR:15 LR:-27.4 LO:36.71);ALT=C[chr3:50649062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	50655215	+	chr3	50677795	+	.	11	14	1405887_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1405887_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_50641501_50666501_115C;SPAN=22580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:14 DR:11 LR:-52.2 LO:52.37);ALT=G[chr3:50677795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51422879	+	chr3	51425166	+	.	13	0	1408553_1	10.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=1408553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:51422879(+)-3:51425166(-)__3_51401001_51426001D;SPAN=2287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:120 GQ:10.4 PL:[10.4, 0.0, 281.0] SR:0 DR:13 LR:-10.4 LO:25.69);ALT=G[chr3:51425166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51423766	+	chr3	51425167	+	.	2	19	1408556_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1408556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51401001_51426001_5C;SPAN=1401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:113 GQ:38.9 PL:[38.9, 0.0, 233.6] SR:19 DR:2 LR:-38.71 LO:46.84);ALT=G[chr3:51425167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51425309	+	chr3	51426335	+	.	0	5	1408571_1	1.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1408571_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51425501_51450501_236C;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:5 DR:0 LR:-1.062 LO:9.396);ALT=G[chr3:51426335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51705945	+	chr3	51708283	+	.	21	0	1409683_1	44.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1409683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:51705945(+)-3:51708283(-)__3_51695001_51720001D;SPAN=2338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:90 GQ:44.9 PL:[44.9, 0.0, 173.6] SR:0 DR:21 LR:-44.94 LO:49.2);ALT=C[chr3:51708283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51972222	+	chr3	51975425	+	.	0	8	1410549_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1410549_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51964501_51989501_352C;SPAN=3203;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:8 DR:0 LR:-4.192 LO:15.42);ALT=T[chr3:51975425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	51972266	+	chr3	51975842	+	.	11	0	1410550_1	6.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1410550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:51972266(+)-3:51975842(-)__3_51964501_51989501D;SPAN=3576;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:112 GQ:6.2 PL:[6.2, 0.0, 263.6] SR:0 DR:11 LR:-5.968 LO:21.24);ALT=C[chr3:51975842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52004203	+	chr3	52005474	+	.	0	16	1410896_1	19.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=1410896_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51989001_52014001_29C;SPAN=1271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:125 GQ:19.1 PL:[19.1, 0.0, 283.1] SR:16 DR:0 LR:-18.95 LO:32.85);ALT=G[chr3:52005474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52004251	+	chr3	52007977	+	.	28	0	1410897_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1410897_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52004251(+)-3:52007977(-)__3_51989001_52014001D;SPAN=3726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:128 GQ:57.8 PL:[57.8, 0.0, 252.5] SR:0 DR:28 LR:-57.75 LO:64.7);ALT=A[chr3:52007977[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52005866	+	chr3	52007978	+	.	97	0	1410901_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1410901_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52005866(+)-3:52007978(-)__3_51989001_52014001D;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:118 GQ:2.1 PL:[290.4, 2.1, 0.0] SR:0 DR:97 LR:-306.6 LO:306.6);ALT=G[chr3:52007978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52009220	+	chr3	52011886	+	.	42	12	1410917_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1410917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_51989001_52014001_151C;SPAN=2666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:112 GQ:99 PL:[118.4, 0.0, 151.4] SR:12 DR:42 LR:-118.2 LO:118.5);ALT=G[chr3:52011886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52018175	+	chr3	52019222	+	.	0	9	1411261_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=1411261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_52013501_52038501_214C;SPAN=1047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:101 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:9 DR:0 LR:-2.346 LO:16.98);ALT=G[chr3:52019222[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52184040	+	chr3	52188368	+	.	9	0	1411542_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1411542_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52184040(+)-3:52188368(-)__3_52185001_52210001D;SPAN=4328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:0 DR:9 LR:-14.0 LO:19.3);ALT=A[chr3:52188368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52266139	+	chr3	52269045	+	.	2	84	1411871_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1411871_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_52258501_52283501_34C;SPAN=2906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:149 GQ:99 PL:[240.2, 0.0, 121.4] SR:84 DR:2 LR:-242.3 LO:242.3);ALT=C[chr3:52269045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52266194	+	chr3	52273015	+	.	105	0	1411874_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1411874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52266194(+)-3:52273015(-)__3_52258501_52283501D;SPAN=6821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:103 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:0 DR:105 LR:-310.3 LO:310.3);ALT=G[chr3:52273015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52269123	+	chr3	52273008	+	.	51	35	1411885_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1411885_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_52258501_52283501_34C;SPAN=3885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:94 GQ:67.1 PL:[159.5, 0.0, 67.1] SR:35 DR:51 LR:-161.3 LO:161.3);ALT=C[chr3:52273008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52489752	+	chr3	52491858	+	.	4	4	1412690_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1412690_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_52479001_52504001_64C;SPAN=2106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:103 GQ:11.1 PL:[0.0, 11.1, 270.6] SR:4 DR:4 LR:11.4 LO:8.071);ALT=T[chr3:52491858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52570789	+	chr3	52574437	+	.	6	7	1412902_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1412902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_52552501_52577501_108C;SPAN=3648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:124 GQ:2.9 PL:[2.9, 0.0, 296.6] SR:7 DR:6 LR:-2.716 LO:20.73);ALT=G[chr3:52574437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52713743	+	chr3	52719765	+	.	0	7	1413597_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1413597_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_52699501_52724501_129C;SPAN=6022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:7 DR:0 LR:0.4634 LO:12.88);ALT=C[chr3:52719765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52720121	+	chr3	52721260	+	AGTTAAAGAAAGCAAGTAAACGCATGACCTGCCATAAGCGGTATAAAATCCAAAAAA	17	15	1413616_1	67.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=AGTTAAAGAAAGCAAGTAAACGCATGACCTGCCATAAGCGGTATAAAATCCAAAAAA;MAPQ=60;MATEID=1413616_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_52699501_52724501_147C;SPAN=1139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:82 GQ:67.1 PL:[67.1, 0.0, 129.8] SR:15 DR:17 LR:-66.91 LO:68.08);ALT=A[chr3:52721260[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	52740305	+	chr3	52741701	+	.	11	0	1413700_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1413700_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:52740305(+)-3:52741701(-)__3_52724001_52749001D;SPAN=1396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:156 GQ:5.8 PL:[0.0, 5.8, 389.4] SR:0 DR:11 LR:5.953 LO:19.59);ALT=G[chr3:52741701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53260896	+	chr3	53262072	+	.	4	18	1415715_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1415715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53238501_53263501_270C;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:119 GQ:40.4 PL:[40.4, 0.0, 248.3] SR:18 DR:4 LR:-40.38 LO:49.02);ALT=T[chr3:53262072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53260937	+	chr3	53262289	+	.	13	0	1415716_1	13.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1415716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53260937(+)-3:53262289(-)__3_53238501_53263501D;SPAN=1352;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:110 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:0 DR:13 LR:-13.11 LO:26.21);ALT=C[chr3:53262289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53263453	+	chr3	53264471	+	.	0	13	1415733_1	13.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=1415733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53263001_53288001_97C;SPAN=1018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:111 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:13 DR:0 LR:-12.84 LO:26.15);ALT=C[chr3:53264471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53264639	+	chr3	53267171	+	TGTCCCCAACTTTGTAGCTGGGCAGGCTGGGCATGCGGATGTTGGCAATGTCCACTGAGGGTGCGTCCTCCTGTGGAGGGGTTGCCAGGATCTTCTTTTTGCTCTGGATCTGGCTGTAGATCTCCTGGATGATCTGCTCAGCCATGTTTTTGGGGAGGGGCTTCCCATGCCAAGACTCCTTATCTTCTACC	2	33	1415739_1	76.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGTCCCCAACTTTGTAGCTGGGCAGGCTGGGCATGCGGATGTTGGCAATGTCCACTGAGGGTGCGTCCTCCTGTGGAGGGGTTGCCAGGATCTTCTTTTTGCTCTGGATCTGGCTGTAGATCTCCTGGATGATCTGCTCAGCCATGTTTTTGGGGAGGGGCTTCCCATGCCAAGACTCCTTATCTTCTACC;MAPQ=60;MATEID=1415739_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_53263001_53288001_464C;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:122 GQ:76.1 PL:[76.1, 0.0, 218.0] SR:33 DR:2 LR:-75.88 LO:79.79);ALT=T[chr3:53267171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53265567	+	chr3	53267171	+	.	6	24	1415743_1	58.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=1415743_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCCC;SCTG=c_3_53263001_53288001_464C;SPAN=1604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:126 GQ:58.4 PL:[58.4, 0.0, 246.5] SR:24 DR:6 LR:-58.29 LO:64.92);ALT=C[chr3:53267171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53265601	+	chr3	53268998	+	.	8	0	1415744_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1415744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53265601(+)-3:53268998(-)__3_53263001_53288001D;SPAN=3397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:104 GQ:1.5 PL:[0.0, 1.5, 254.1] SR:0 DR:8 LR:1.768 LO:14.56);ALT=T[chr3:53268998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53267291	+	chr3	53268999	+	.	16	12	1415748_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1415748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53263001_53288001_384C;SPAN=1708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:113 GQ:48.8 PL:[48.8, 0.0, 223.7] SR:12 DR:16 LR:-48.61 LO:55.1);ALT=C[chr3:53268999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53275312	+	chr3	53289851	+	.	76	0	1416153_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1416153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53275312(+)-3:53289851(-)__3_53287501_53312501D;SPAN=14539;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:87 GQ:16.8 PL:[244.2, 16.8, 0.0] SR:0 DR:76 LR:-246.4 LO:246.4);ALT=T[chr3:53289851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53312247	+	chr3	53315559	+	.	41	37	1416276_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AAGTGATC;MAPQ=27;MATEID=1416276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53287501_53312501_18C;SPAN=3312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:29 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:37 DR:41 LR:-188.1 LO:188.1);ALT=C[chr3:53315559[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53902891	+	chr3	53904008	+	.	0	6	1418076_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1418076_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_53900001_53925001_45C;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:123 GQ:13.2 PL:[0.0, 13.2, 323.4] SR:6 DR:0 LR:13.52 LO:9.698);ALT=T[chr3:53904008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53919590	+	chr3	53925796	+	TCCTCATCCACCAGCCATTGGAGGGGGACTAGGGCCACGCAGATGATTGATTCTACCCATTCTTCGGGGAGGGTTTCCTGGTGGCCCTCTTCCATCATCATATCTGGAATCAGATGAGTTTCCATAGCTTCTTCTTTTTTTCACATCTTGCTGAAGCAGAGTTTTGAAAAACAAAACCACAAACTCAGCTATTCCCCAGAAGAAATCTGTTATCAAAGATAATCTCCATGGAGACTGACTCCGGCTGTCCAACACTTGT	0	21	1418226_1	53.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCGTTCGAGATGTAAACCATCTTG;INSERTION=TCCTCATCCACCAGCCATTGGAGGGGGACTAGGGCCACGCAGATGATTGATTCTACCCATTCTTCGGGGAGGGTTTCCTGGTGGCCCTCTTCCATCATCATATCTGGAATCAGATGAGTTTCCATAGCTTCTTCTTTTTTTCACATCTTGCTGAAGCAGAGTTTTGAAAAACAAAACCACAAACTCAGCTATTCCCCAGAAGAAATCTGTTATCAAAGATAATCTCCATGGAGACTGACTCCGGCTGTCCAACACTTGT;MAPQ=60;MATEID=1418226_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_53924501_53949501_423C;SPAN=6206;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:61 GQ:53 PL:[53.0, 0.0, 92.6] SR:21 DR:0 LR:-52.8 LO:53.46);ALT=T[chr3:53925796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53919981	+	chr3	53925795	+	.	19	0	1418228_1	46.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=1418228_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53919981(+)-3:53925795(-)__3_53924501_53949501D;SPAN=5814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:60 GQ:46.4 PL:[46.4, 0.0, 99.2] SR:0 DR:19 LR:-46.46 LO:47.51);ALT=A[chr3:53925795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	53920979	+	chr3	53925794	+	.	29	0	1418229_1	79.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=1418229_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:53920979(+)-3:53925794(-)__3_53924501_53949501D;SPAN=4815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:60 GQ:66.2 PL:[79.4, 0.0, 66.2] SR:0 DR:29 LR:-79.54 LO:79.54);ALT=A[chr3:53925794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38184469	+	chr3	53925796	+	CTCTTCCATCATCATATCTGG	20	12	1418236_1	79.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCGTTCGAGATGTAAACCATCTTG;INSERTION=CTCTTCCATCATCATATCTGG;MAPQ=60;MATEID=1418236_2;MATENM=6;NM=0;NUMPARTS=4;SCTG=c_3_53924501_53949501_423C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:61 GQ:66.2 PL:[79.4, 0.0, 66.2] SR:12 DR:20 LR:-79.24 LO:79.24);ALT=]chr19:38184469]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	28226455	+	chr3	54428356	+	.	13	0	5136534_1	31.0	.	DISC_MAPQ=9;EVDNC=DSCRD;IMPRECISE;MAPQ=9;MATEID=5136534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:54428356(-)-12:28226455(+)__12_28224001_28249001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:42 GQ:31.7 PL:[31.7, 0.0, 68.0] SR:0 DR:13 LR:-31.53 LO:32.35);ALT=]chr12:28226455]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	54512690	-	chr9	118004803	+	.	7	22	1419998_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATATATATATATA;MAPQ=60;MATEID=1419998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_54488001_54513001_374C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:29 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:22 DR:7 LR:-85.54 LO:85.54);ALT=[chr9:118004803[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	54512706	+	chr9	118004854	-	ATAGCAATAT	8	17	1420001_1	54.0	.	DISC_MAPQ=36;EVDNC=TSI_G;HOMSEQ=ATATATATATAT;INSERTION=ATAGCAATAT;MAPQ=56;MATEID=1420001_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_3_54488001_54513001_111C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:29 GQ:15.2 PL:[54.8, 0.0, 15.2] SR:17 DR:8 LR:-56.08 LO:56.08);ALT=T]chr9:118004854];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	56517988	+	chr15	91701885	-	.	10	0	6032864_1	20.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=6032864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:56517988(+)-15:91701885(+)__15_91679001_91704001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:0 DR:10 LR:-20.55 LO:23.07);ALT=A]chr15:91701885];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	57261965	+	chr3	57269591	+	.	27	16	1429405_1	86.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1429405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57256501_57281501_250C;SPAN=7626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:95 GQ:86.6 PL:[86.6, 0.0, 142.7] SR:16 DR:27 LR:-86.5 LO:87.28);ALT=G[chr3:57269591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57261984	+	chr3	57271517	+	.	12	0	1429406_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1429406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:57261984(+)-3:57271517(-)__3_57256501_57281501D;SPAN=9533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:88 GQ:15.8 PL:[15.8, 0.0, 197.3] SR:0 DR:12 LR:-15.77 LO:24.99);ALT=T[chr3:57271517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57269692	+	chr3	57272070	+	AATGAATTAAGTGCAGCAACACACCTGACCTCAAAACTTTTAAAAGAATATGAAAAA	0	38	1429441_1	94.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AATGAATTAAGTGCAGCAACACACCTGACCTCAAAACTTTTAAAAGAATATGAAAAA;MAPQ=60;MATEID=1429441_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_57256501_57281501_101C;SPAN=2378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:115 GQ:94.4 PL:[94.4, 0.0, 183.5] SR:38 DR:0 LR:-94.28 LO:95.89);ALT=G[chr3:57272070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57272144	+	chr3	57276127	+	CTTAGCTCTTGTCATGCAGTGCTTTCAACTCAACTTGCTGATGCCATGATGTTCCCCATTACCCAGTTTAAAGAAAGAGATCTGAA	0	13	1429455_1	15.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTTAGCTCTTGTCATGCAGTGCTTTCAACTCAACTTGCTGATGCCATGATGTTCCCCATTACCCAGTTTAAAGAAAGAGATCTGAA;MAPQ=60;MATEID=1429455_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_57256501_57281501_184C;SPAN=3983;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:101 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:13 DR:0 LR:-15.55 LO:26.73);ALT=G[chr3:57276127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57280250	+	chr3	57281420	+	.	0	4	1429476_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1429476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57256501_57281501_396C;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:4 DR:0 LR:13.62 LO:6.133);ALT=G[chr3:57281420[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	57505598	+	chr3	141457288	-	.	56	0	1691813_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=1691813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:57505598(+)-3:141457288(+)__3_141438501_141463501D;SPAN=83951690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:76 GQ:19.1 PL:[164.3, 0.0, 19.1] SR:0 DR:56 LR:-170.8 LO:170.8);ALT=C]chr3:141457288];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	57524041	+	chr3	57522647	+	CTATGATTAGTGA	16	24	1430533_1	77.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=CTATGATTAGTGA;MAPQ=60;MATEID=1430533_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57501501_57526501_100C;SPAN=1394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:91 GQ:77.9 PL:[77.9, 0.0, 140.6] SR:24 DR:16 LR:-77.68 LO:78.74);ALT=]chr3:57524041]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	57570192	+	chr3	57582801	+	.	0	14	1431040_1	32.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1431040_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_57550501_57575501_251C;SPAN=12609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:51 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:14 DR:0 LR:-32.4 LO:33.96);ALT=C[chr3:57582801[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	58318760	+	chr3	58351599	+	.	9	0	1434041_1	18.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1434041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:58318760(+)-3:58351599(-)__3_58310001_58335001D;SPAN=32839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:43 GQ:18.2 PL:[18.2, 0.0, 84.2] SR:0 DR:9 LR:-18.06 LO:20.6);ALT=C[chr3:58351599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	58318818	+	chr3	58368239	+	AATATATTATTCGAGTGCAAAGAGGAATTTCTGTGGAAAACAGCTGGCAGATTGTTAGAAGATACAGTGACTTTGATTTGCTTAACAACAGCTTAC	0	26	1434044_1	75.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AATATATTATTCGAGTGCAAAGAGGAATTTCTGTGGAAAACAGCTGGCAGATTGTTAGAAGATACAGTGACTTTGATTTGCTTAACAACAGCTTAC;MAPQ=60;MATEID=1434044_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_58310001_58335001_76C;SPAN=49421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:37 GQ:13.1 PL:[75.8, 0.0, 13.1] SR:26 DR:0 LR:-78.22 LO:78.22);ALT=G[chr3:58368239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	58383449	+	chr3	58394649	+	TGGCCGTGTTGGAGTCTACGCTGTCTTGTGAAGCCTGTAAAAATGGCATGCCTACCATCTCCCGGCTCTTACAGATGCCATTATTCAGCGATGTTTTACTAACCACTTCTGAAAAACCACAGTTTA	0	13	1433784_1	21.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGGCCGTGTTGGAGTCTACGCTGTCTTGTGAAGCCTGTAAAAATGGCATGCCTACCATCTCCCGGCTCTTACAGATGCCATTATTCAGCGATGTTTTACTAACCACTTCTGAAAAACCACAGTTTA;MAPQ=60;MATEID=1433784_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_58383501_58408501_289C;SPAN=11200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:79 GQ:21.5 PL:[21.5, 0.0, 170.0] SR:13 DR:0 LR:-21.51 LO:28.24);ALT=G[chr3:58394649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	58417729	+	chr3	58419488	+	.	13	0	1434278_1	12.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1434278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:58417729(+)-3:58419488(-)__3_58408001_58433001D;SPAN=1759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:113 GQ:12.5 PL:[12.5, 0.0, 260.0] SR:0 DR:13 LR:-12.3 LO:26.05);ALT=A[chr3:58419488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	66271554	+	chr3	66286967	+	.	15	5	1459832_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1459832_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_66272501_66297501_9C;SPAN=15413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:57 GQ:44 PL:[44.0, 0.0, 93.5] SR:5 DR:15 LR:-43.98 LO:44.99);ALT=G[chr3:66286967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	66777004	-	chr3	66778062	+	.	8	0	1461680_1	0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=1461680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:66777004(-)-3:66778062(-)__3_66762501_66787501D;SPAN=1058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:0 DR:8 LR:2.581 LO:14.46);ALT=[chr3:66778062[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	67493708	+	chr3	67496800	+	.	47	25	1463988_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAATTAGATCTC;MAPQ=60;MATEID=1463988_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_67473001_67498001_289C;SPAN=3092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:58 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:25 DR:47 LR:-178.2 LO:178.2);ALT=C[chr3:67496800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	67660013	+	chr3	67704960	+	.	12	0	1464464_1	25.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1464464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:67660013(+)-3:67704960(-)__3_67693501_67718501D;SPAN=44947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:54 GQ:25.1 PL:[25.1, 0.0, 104.3] SR:0 DR:12 LR:-24.98 LO:27.82);ALT=T[chr3:67704960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69127063	+	chr3	69129483	+	.	10	0	1469140_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1469140_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:69127063(+)-3:69129483(-)__3_69114501_69139501D;SPAN=2420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.918 LO:19.39);ALT=A[chr3:69129483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69134376	+	chr3	69153615	+	TTCTGAGTCCCTTCAACATGATCCTGGGAGGAATCGTGGTGGTGCTGGTGTTCACAGGGTTTGTGTGGGCAGCCCACAATAAAGACGTCCTTCGCCGGATGAAGAAGCGCTACCCCACGACGTTCGTTATGGTGGTCATGTTGGCGAGCTATTTCCTTATCTCCATGTTTGGAGGAGTCATGGTCTTTGTGTTTGGCATTACTTTTCCTTTGCTGT	2	97	1469161_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=TTCTGAGTCCCTTCAACATGATCCTGGGAGGAATCGTGGTGGTGCTGGTGTTCACAGGGTTTGTGTGGGCAGCCCACAATAAAGACGTCCTTCGCCGGATGAAGAAGCGCTACCCCACGACGTTCGTTATGGTGGTCATGTTGGCGAGCTATTTCCTTATCTCCATGTTTGGAGGAGTCATGGTCTTTGTGTTTGGCATTACTTTTCCTTTGCTGT;MAPQ=60;MATEID=1469161_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_69114501_69139501_192C;SPAN=19239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:87 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:97 DR:2 LR:-293.8 LO:293.8);ALT=T[chr3:69153615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69134376	+	chr3	69150989	+	.	68	91	1469160_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=1469160_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_69114501_69139501_192C;SPAN=16613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:87 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:91 DR:68 LR:-406.0 LO:406.0);ALT=T[chr3:69150989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69151207	+	chr3	69153615	+	.	6	9	1469257_1	7.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=1469257_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_69139001_69164001_151C;SPAN=2408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:107 GQ:7.4 PL:[7.4, 0.0, 251.6] SR:9 DR:6 LR:-7.322 LO:21.47);ALT=T[chr3:69153615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	69383619	+	chr3	69402695	+	.	25	11	1470146_1	80.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1470146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_69359501_69384501_170C;SPAN=19076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:57 GQ:57.2 PL:[80.3, 0.0, 57.2] SR:11 DR:25 LR:-80.48 LO:80.48);ALT=T[chr3:69402695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	9666569	+	chr3	75606411	+	.	10	0	1491480_1	20.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=1491480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:75606411(-)-4:9666569(+)__3_75582501_75607501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=]chr4:9666569]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	94226377	+	chr7	102715698	-	.	10	0	3496225_1	20.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3496225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:94226377(+)-7:102715698(+)__7_102704001_102729001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:0 DR:10 LR:-20.55 LO:23.07);ALT=C]chr7:102715698];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	95214730	-	chr3	95216336	+	.	12	0	1539890_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1539890_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:95214730(-)-3:95216336(-)__3_95207001_95232001D;SPAN=1606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:128 GQ:5 PL:[5.0, 0.0, 305.3] SR:0 DR:12 LR:-4.934 LO:22.91);ALT=[chr3:95216336[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	95465768	+	chr3	95470764	+	.	53	45	1540653_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CAAG;MAPQ=60;MATEID=1540653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_95C;SPAN=4996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:104 GQ:8.1 PL:[267.3, 8.1, 0.0] SR:45 DR:53 LR:-276.8 LO:276.8);ALT=G[chr3:95470764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	95471000	+	chr3	95468117	+	TGCATAGGG	43	35	1540655_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGCATAGGG;MAPQ=60;MATEID=1540655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_95452001_95477001_267C;SPAN=2883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:97 GQ:72.8 PL:[161.9, 0.0, 72.8] SR:35 DR:43 LR:-163.7 LO:163.7);ALT=]chr3:95471000]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	97921336	+	chr3	97882020	+	.	16	0	1548009_1	43.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=1548009_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:97882020(-)-3:97921336(+)__3_97902001_97927001D;SPAN=39316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:34 GQ:37.1 PL:[43.7, 0.0, 37.1] SR:0 DR:16 LR:-43.62 LO:43.62);ALT=]chr3:97921336]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	98240187	+	chr3	98241691	+	.	9	0	1548481_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1548481_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:98240187(+)-3:98241691(-)__3_98220501_98245501D;SPAN=1504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:127 GQ:4.5 PL:[0.0, 4.5, 316.8] SR:0 DR:9 LR:4.698 LO:16.05);ALT=C[chr3:98241691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	98899063	+	chr3	98902390	+	.	43	29	1550958_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=1550958_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_98882001_98907001_475C;SPAN=3327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:57 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:29 DR:43 LR:-168.3 LO:168.3);ALT=T[chr3:98902390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	98899160	-	chr5	54764402	+	CACCTCA	6	52	1550966_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=CACCTCA;MAPQ=60;MATEID=1550966_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_3_98882001_98907001_145C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:15 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:52 DR:6 LR:-168.3 LO:168.3);ALT=[chr5:54764402[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	99536887	+	chr3	99865815	+	.	0	26	1553553_1	70.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1553553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_99862001_99887001_56C;SPAN=328928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:58 GQ:70.1 PL:[70.1, 0.0, 70.1] SR:26 DR:0 LR:-70.11 LO:70.11);ALT=G[chr3:99865815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	100053684	+	chr3	100057936	+	.	18	0	1554360_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1554360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:100053684(+)-3:100057936(-)__3_100058001_100083001D;SPAN=4252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:13 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=C[chr3:100057936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	100053691	+	chr3	100058657	+	.	42	0	1554362_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1554362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:100053691(+)-3:100058657(-)__3_100058001_100083001D;SPAN=4966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:58 GQ:17.3 PL:[122.9, 0.0, 17.3] SR:0 DR:42 LR:-127.4 LO:127.4);ALT=G[chr3:100058657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	100071347	+	chr3	100074019	+	GGGGAGGTTCTAGCCAAAGCTGGCACAGAAGAAGCAATCGTGTATTCAGACAT	0	70	1554435_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GGGGAGGTTCTAGCCAAAGCTGGCACAGAAGAAGCAATCGTGTATTCAGACAT;MAPQ=60;MATEID=1554435_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_100058001_100083001_101C;SPAN=2672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:124 GQ:99 PL:[197.6, 0.0, 101.9] SR:70 DR:0 LR:-199.1 LO:199.1);ALT=G[chr3:100074019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	100384270	+	chr14	54955636	+	.	8	0	5748626_1	13.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=5748626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:100384270(+)-14:54955636(-)__14_54953501_54978501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=G[chr14:54955636[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	101280848	+	chr3	101283613	+	.	15	8	1558261_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1558261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_101283001_101308001_395C;SPAN=2765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:57 GQ:44 PL:[44.0, 0.0, 93.5] SR:8 DR:15 LR:-43.98 LO:44.99);ALT=G[chr3:101283613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	101293131	+	chr3	101298430	+	.	59	0	1558296_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1558296_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101293131(+)-3:101298430(-)__3_101283001_101308001D;SPAN=5299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:105 GQ:87.2 PL:[166.4, 0.0, 87.2] SR:0 DR:59 LR:-167.6 LO:167.6);ALT=C[chr3:101298430[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	101293152	+	chr13	48902558	-	.	41	0	5490003_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5490003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101293152(+)-13:48902558(+)__13_48877501_48902501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:18 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=C]chr13:48902558];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	42924510	+	chr3	101405405	+	.	38	0	2819974_1	67.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2819974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:101405405(-)-6:42924510(+)__6_42899501_42924501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:213 GQ:67.9 PL:[67.9, 0.0, 447.5] SR:0 DR:38 LR:-67.73 LO:84.01);ALT=]chr6:42924510]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	101576303	+	chr3	101578159	+	.	4	7	1559554_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1559554_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_101577001_101602001_286C;SPAN=1856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:69 GQ:14.3 PL:[14.3, 0.0, 152.9] SR:7 DR:4 LR:-14.32 LO:21.12);ALT=G[chr3:101578159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	105586450	+	chr3	105587738	+	.	14	0	1571105_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1571105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:105586450(+)-3:105587738(-)__3_105570501_105595501D;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:108 GQ:17 PL:[17.0, 0.0, 244.7] SR:0 DR:14 LR:-16.95 LO:28.83);ALT=T[chr3:105587738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141379675	+	chr3	105828855	+	.	21	0	2599308_1	59.0	.	DISC_MAPQ=9;EVDNC=DSCRD;IMPRECISE;MAPQ=9;MATEID=2599308_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:105828855(-)-5:141379675(+)__5_141365001_141390001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:21 DP:20 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:21 LR:-59.41 LO:59.41);ALT=]chr5:141379675]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	119396187	-	chr13	47065110	+	.	9	0	1614989_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1614989_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:119396187(-)-13:47065110(-)__3_119388501_119413501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:0 DR:9 LR:-10.2 LO:18.38);ALT=[chr13:47065110[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	119431705	+	chr21	30382812	+	.	14	44	7151769_1	99.0	.	DISC_MAPQ=8;EVDNC=ASDIS;HOMSEQ=TCCCAGCTACTTGGGAGGCTGAG;MAPQ=30;MATEID=7151769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_30380001_30405001_72C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:40 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:44 DR:14 LR:-145.2 LO:145.2);ALT=G[chr21:30382812[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	120315279	+	chr4	43901106	+	.	23	0	1952936_1	65.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1952936_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:120315279(+)-4:43901106(-)__4_43879501_43904501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:0 DR:23 LR:-65.7 LO:65.7);ALT=A[chr4:43901106[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	120315385	+	chr3	120319956	+	.	36	0	1618392_1	86.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1618392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:120315385(+)-3:120319956(-)__3_120295001_120320001D;SPAN=4571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:121 GQ:86.3 PL:[86.3, 0.0, 205.1] SR:0 DR:36 LR:-86.05 LO:88.83);ALT=T[chr3:120319956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121352020	+	chr3	121353053	+	.	8	11	1621334_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1621334_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121348501_121373501_399C;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:111 GQ:19.7 PL:[19.7, 0.0, 247.4] SR:11 DR:8 LR:-19.44 LO:31.18);ALT=T[chr3:121353053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121353266	+	chr3	121355281	+	AGCTTCTATGGGCGTCGTCTTCTTATAAGCTGTGGTCGGGGCCTCCATTTCATTGAAGCCGACAGCGCT	3	36	1621342_1	84.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AGCTTCTATGGGCGTCGTCTTCTTATAAGCTGTGGTCGGGGCCTCCATTTCATTGAAGCCGACAGCGCT;MAPQ=60;MATEID=1621342_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_3_121348501_121373501_48C;SPAN=2015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:140 GQ:84.2 PL:[84.2, 0.0, 255.8] SR:36 DR:3 LR:-84.21 LO:89.02);ALT=C[chr3:121355281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121353266	+	chr3	121354584	+	A	2	34	1621341_1	77.0	.	DISC_MAPQ=41;EVDNC=TSI_L;INSERTION=A;MAPQ=60;MATEID=1621341_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_3_121348501_121373501_48C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:142 GQ:77.3 PL:[77.3, 0.0, 265.4] SR:34 DR:2 LR:-77.06 LO:82.96);ALT=C[chr3:121354584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121353307	+	chr3	121355992	+	.	9	0	1621344_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1621344_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121353307(+)-3:121355992(-)__3_121348501_121373501D;SPAN=2685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:111 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.3636 LO:16.59);ALT=G[chr3:121355992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121356105	+	chr3	121366166	+	TTCTGAGATGTGTGCTTCTCCACTTCTCCTTTATAATCAAAGCCGACTGCTGACTTGTCTGCCCTGTCCCTCTCAACTCCGTACTTGCCCCCAAAGCCTTTGGCAGCATCCGTCTGAGAAGAGTGCTTCTCCACCTCGGCAACATACTCATGGCCCACTGCACT	0	36	1621361_1	83.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTCTGAGATGTGTGCTTCTCCACTTCTCCTTTATAATCAAAGCCGACTGCTGACTTGTCTGCCCTGTCCCTCTCAACTCCGTACTTGCCCCCAAAGCCTTTGGCAGCATCCGTCTGAGAAGAGTGCTTCTCCACCTCGGCAACATACTCATGGCCCACTGCACT;MAPQ=60;MATEID=1621361_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_121348501_121373501_53C;SPAN=10061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:130 GQ:83.6 PL:[83.6, 0.0, 232.1] SR:36 DR:0 LR:-83.62 LO:87.48);ALT=T[chr3:121366166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121363777	+	chr3	121366166	+	.	4	15	1621403_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1621403_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TCTC;SCTG=c_3_121348501_121373501_53C;SPAN=2389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:121 GQ:30.2 PL:[30.2, 0.0, 261.2] SR:15 DR:4 LR:-29.94 LO:40.84);ALT=T[chr3:121366166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121366295	+	chr3	121376126	+	.	0	64	1621518_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1621518_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121373001_121398001_425C;SPAN=9831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:77 GQ:4.2 PL:[194.7, 4.2, 0.0] SR:64 DR:0 LR:-203.1 LO:203.1);ALT=G[chr3:121376126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121366339	+	chr3	121379674	+	.	36	0	1621519_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1621519_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121366339(+)-3:121379674(-)__3_121373001_121398001D;SPAN=13335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:62 GQ:46.1 PL:[102.2, 0.0, 46.1] SR:0 DR:36 LR:-103.1 LO:103.1);ALT=T[chr3:121379674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121376246	+	chr3	121379670	+	.	63	0	1621541_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1621541_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121376246(+)-3:121379670(-)__3_121373001_121398001D;SPAN=3424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:115 GQ:99 PL:[176.9, 0.0, 101.0] SR:0 DR:63 LR:-177.9 LO:177.9);ALT=A[chr3:121379670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121377196	+	chr3	121379667	+	.	34	13	1621548_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1621548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121373001_121398001_176C;SPAN=2471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:127 GQ:84.5 PL:[84.5, 0.0, 223.1] SR:13 DR:34 LR:-84.43 LO:87.92);ALT=T[chr3:121379667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121547820	+	chr3	121553235	+	.	0	10	1622073_1	4.0	.	EVDNC=ASSMB;HOMSEQ=TACC;MAPQ=60;MATEID=1622073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121544501_121569501_152C;SPAN=5415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:10 DR:0 LR:-4.292 LO:19.12);ALT=C[chr3:121553235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121547863	+	chr3	121553817	+	.	8	0	1622075_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1622075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121547863(+)-3:121553817(-)__3_121544501_121569501D;SPAN=5954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:0 DR:8 LR:2.581 LO:14.46);ALT=A[chr3:121553817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121554238	+	chr3	121563300	+	.	39	39	1622097_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=1622097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121544501_121569501_65C;SPAN=9062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:110 GQ:99 PL:[148.4, 0.0, 118.7] SR:39 DR:39 LR:-148.6 LO:148.6);ALT=T[chr3:121563300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121563394	+	chr3	121575858	+	.	0	11	1622229_1	20.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1622229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121569001_121594001_202C;SPAN=12464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:61 GQ:20 PL:[20.0, 0.0, 125.6] SR:11 DR:0 LR:-19.78 LO:24.38);ALT=A[chr3:121575858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121563395	+	chr3	121573534	+	.	0	13	1622230_1	31.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1622230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121569001_121594001_418C;SPAN=10139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:43 GQ:31.4 PL:[31.4, 0.0, 71.0] SR:13 DR:0 LR:-31.26 LO:32.19);ALT=G[chr3:121573534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121774300	+	chr3	121822357	+	.	12	0	1622848_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1622848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121774300(+)-3:121822357(-)__3_121814001_121839001D;SPAN=48057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:49 GQ:26.3 PL:[26.3, 0.0, 92.3] SR:0 DR:12 LR:-26.34 LO:28.41);ALT=C[chr3:121822357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121796824	+	chr3	121822357	+	.	9	0	1622849_1	16.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1622849_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:121796824(+)-3:121822357(-)__3_121814001_121839001D;SPAN=25533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=T[chr3:121822357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	121825347	+	chr3	121828109	+	.	3	11	1622878_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAG;MAPQ=60;MATEID=1622878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_121814001_121839001_301C;SPAN=2762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:107 GQ:10.7 PL:[10.7, 0.0, 248.3] SR:11 DR:3 LR:-10.62 LO:23.9);ALT=G[chr3:121828109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122044207	+	chr3	122056392	+	.	33	30	1623628_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1623628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122034501_122059501_147C;SPAN=12185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:113 GQ:99 PL:[134.6, 0.0, 137.9] SR:30 DR:33 LR:-134.4 LO:134.4);ALT=T[chr3:122056392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122044235	+	chr3	122060281	+	.	71	0	1623683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1623683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:122044235(+)-3:122060281(-)__3_122059001_122084001D;SPAN=16046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:55 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=G[chr3:122060281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122056497	+	chr3	122060284	+	.	2	28	1623667_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1623667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122034501_122059501_141C;SPAN=3787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:61 GQ:62.9 PL:[82.7, 0.0, 62.9] SR:28 DR:2 LR:-82.61 LO:82.61);ALT=T[chr3:122060284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122103147	+	chr3	122121605	+	.	53	10	1623847_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1623847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122108001_122133001_270C;SPAN=18458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:56 GQ:15 PL:[165.0, 15.0, 0.0] SR:10 DR:53 LR:-165.0 LO:165.0);ALT=G[chr3:122121605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122103185	+	chr3	122123104	+	.	32	0	1623849_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1623849_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:122103185(+)-3:122123104(-)__3_122108001_122133001D;SPAN=19919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:51 GQ:29.3 PL:[92.0, 0.0, 29.3] SR:0 DR:32 LR:-93.4 LO:93.4);ALT=G[chr3:122123104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122121730	+	chr3	122123105	+	.	3	45	1623909_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1623909_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122108001_122133001_122C;SPAN=1375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:119 GQ:99 PL:[126.2, 0.0, 162.5] SR:45 DR:3 LR:-126.2 LO:126.5);ALT=G[chr3:122123105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122123212	+	chr3	122126128	+	.	0	27	1623914_1	62.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=1623914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122108001_122133001_75C;SPAN=2916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:99 GQ:62.3 PL:[62.3, 0.0, 177.8] SR:27 DR:0 LR:-62.31 LO:65.4);ALT=T[chr3:122126128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122126237	+	chr3	122128584	+	.	0	30	1623925_1	70.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1623925_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122108001_122133001_136C;SPAN=2347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:107 GQ:70.1 PL:[70.1, 0.0, 188.9] SR:30 DR:0 LR:-70.04 LO:73.1);ALT=G[chr3:122128584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122215418	+	chr3	122233604	+	.	0	7	1624318_1	13.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1624318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122230501_122255501_406C;SPAN=18186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:35 GQ:13.7 PL:[13.7, 0.0, 69.8] SR:7 DR:0 LR:-13.62 LO:15.86);ALT=C[chr3:122233604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122296700	+	chr3	122324782	+	.	0	8	1624593_1	12.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1624593_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122304001_122329001_423C;SPAN=28082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:8 DR:0 LR:-12.05 LO:17.05);ALT=G[chr3:122324782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122786056	+	chr3	122808014	+	.	5	3	1626325_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=1626325_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122794001_122819001_147C;SPAN=21958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:3 DR:5 LR:-10.37 LO:14.87);ALT=G[chr3:122808014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	122861362	-	chr3	122862666	+	CTGTCCAGAGGAGGAG	4	8	1626476_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGTCCAGAGGAGGAG;MAPQ=60;MATEID=1626476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_122843001_122868001_81C;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:127 GQ:1.2 PL:[0.0, 1.2, 310.2] SR:8 DR:4 LR:1.397 LO:18.3);ALT=[chr3:122862666[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	123675651	+	chr3	123679997	+	.	11	0	1629414_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1629414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:123675651(+)-3:123679997(-)__3_123676001_123701001D;SPAN=4346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:71 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:0 DR:11 LR:-17.08 LO:23.58);ALT=T[chr3:123679997[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	133382791	+	chr3	124470194	+	.	0	21	4463301_1	54.0	.	EVDNC=ASSMB;HOMSEQ=GAGAGGGAGAGGGA;MAPQ=60;MATEID=4463301_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_133378001_133403001_439C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:56 GQ:54.2 PL:[54.2, 0.0, 80.6] SR:21 DR:0 LR:-54.15 LO:54.46);ALT=]chr9:133382791]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	125050083	+	chr3	125093945	+	.	0	7	1634502_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1634502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_125072501_125097501_232C;SPAN=43862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:52 GQ:9.2 PL:[9.2, 0.0, 114.8] SR:7 DR:0 LR:-9.019 LO:14.54);ALT=C[chr3:125093945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	125438323	+	chr3	125416084	+	.	8	0	1635974_1	0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=1635974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:125416084(-)-3:125438323(+)__3_125415501_125440501D;SPAN=22239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:0 DR:8 LR:0.4135 LO:14.74);ALT=]chr3:125438323]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	125462253	+	chr3	125439593	+	.	25	0	1636769_1	62.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=1636769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:125439593(-)-3:125462253(+)__3_125440001_125465001D;SPAN=22660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:76 GQ:62 PL:[62.0, 0.0, 121.4] SR:0 DR:25 LR:-61.94 LO:63.03);ALT=]chr3:125462253]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	126423191	+	chr3	126445919	+	.	10	0	1639900_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1639900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:126423191(+)-3:126445919(-)__3_126444501_126469501D;SPAN=22728;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=G[chr3:126445919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127318391	+	chr3	127323449	+	.	0	7	1642647_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1642647_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127302001_127327001_264C;SPAN=5058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=G[chr3:127323449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127391926	+	chr3	127394812	+	ACCTGCTGGAGCAGCGAGACGTGGAGGTACTATGCCTGCTTGTGTGGGCACGAGGAGCTGGTACTCTACCTTCTGGCCAAT	16	16	1643012_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ACCTGCTGGAGCAGCGAGACGTGGAGGTACTATGCCTGCTTGTGTGGGCACGAGGAGCTGGTACTCTACCTTCTGGCCAAT;MAPQ=60;MATEID=1643012_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_127375501_127400501_340C;SPAN=2886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:92 GQ:57.8 PL:[57.8, 0.0, 163.4] SR:16 DR:16 LR:-57.6 LO:60.51);ALT=T[chr3:127394812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127411168	+	chr3	127413818	+	.	0	14	1643089_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1643089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127400001_127425001_17C;SPAN=2650;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:14 DR:0 LR:-18.58 LO:29.2);ALT=T[chr3:127413818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127500738	+	chr3	127540536	+	.	0	15	1643463_1	33.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1643463_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127522501_127547501_363C;SPAN=39798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:61 GQ:33.2 PL:[33.2, 0.0, 112.4] SR:15 DR:0 LR:-32.99 LO:35.54);ALT=C[chr3:127540536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127500785	+	chr3	127541964	+	.	14	0	1643464_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1643464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:127500785(+)-3:127541964(-)__3_127522501_127547501D;SPAN=41179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:29 GQ:31.7 PL:[38.3, 0.0, 31.7] SR:0 DR:14 LR:-38.39 LO:38.39);ALT=T[chr3:127541964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127540682	+	chr3	127541926	+	.	43	21	1643512_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1643512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127522501_127547501_87C;SPAN=1244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:113 GQ:99 PL:[131.3, 0.0, 141.2] SR:21 DR:43 LR:-131.1 LO:131.2);ALT=C[chr3:127541926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127831865	+	chr3	127838171	+	.	0	10	1644443_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1644443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127816501_127841501_325C;SPAN=6306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:117 GQ:1.4 PL:[1.4, 0.0, 281.9] SR:10 DR:0 LR:-1.312 LO:18.67);ALT=T[chr3:127838171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	127838259	+	chr3	127842426	+	.	0	19	1644654_1	44.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1644654_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_127841001_127866001_20C;SPAN=4167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:66 GQ:44.9 PL:[44.9, 0.0, 114.2] SR:19 DR:0 LR:-44.84 LO:46.56);ALT=T[chr3:127842426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	64220892	+	chr3	128306019	+	.	8	0	6470752_1	18.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6470752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:128306019(-)-17:64220892(+)__17_64214501_64239501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=]chr17:64220892]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	128341254	+	chr3	128344376	+	.	4	2	1646090_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1646090_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128331001_128356001_401C;SPAN=3122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:117 GQ:15 PL:[0.0, 15.0, 313.5] SR:2 DR:4 LR:15.19 LO:7.789);ALT=T[chr3:128344376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128351003	+	chr3	128356641	+	.	4	3	1646793_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=1646793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128355501_128380501_195C;SPAN=5638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:3 DR:4 LR:-10.37 LO:14.87);ALT=G[chr3:128356641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128356950	+	chr3	128363762	+	.	4	8	1646799_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1646799_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128355501_128380501_500C;SPAN=6812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:111 GQ:6.5 PL:[6.5, 0.0, 260.6] SR:8 DR:4 LR:-6.238 LO:21.28);ALT=T[chr3:128363762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128363828	+	chr3	128369381	+	.	0	27	1646835_1	60.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=1646835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128355501_128380501_443C;SPAN=5553;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:106 GQ:60.5 PL:[60.5, 0.0, 195.8] SR:27 DR:0 LR:-60.41 LO:64.45);ALT=T[chr3:128369381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128445118	+	chr3	128514201	+	.	49	0	1646917_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1646917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:128445118(+)-3:128514201(-)__3_128502501_128527501D;SPAN=69083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:66 GQ:15.2 PL:[143.9, 0.0, 15.2] SR:0 DR:49 LR:-149.8 LO:149.8);ALT=C[chr3:128514201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128445193	+	chr3	128516784	+	.	25	0	1646918_1	63.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1646918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:128445193(+)-3:128516784(-)__3_128502501_128527501D;SPAN=71591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:72 GQ:63.2 PL:[63.2, 0.0, 109.4] SR:0 DR:25 LR:-63.02 LO:63.76);ALT=A[chr3:128516784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128445202	+	chr3	128525212	+	TTTGAAGGATGACCTCTAGGAAGAAAGTGTTGCTGAAGGTTATCATCCTGGGAGATTCTGGAGTCGGGAAGACATCACTCATGAACCAGTATGTGAATAAGAAATTCAGCAATCAGTACAAAGCCACAATAGGAGCTGACTTTCTGACCAAGGAGGTGATGGTGGATGACAGGCTAGTCACAATG	0	72	1646920_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=TTTGAAGGATGACCTCTAGGAAGAAAGTGTTGCTGAAGGTTATCATCCTGGGAGATTCTGGAGTCGGGAAGACATCACTCATGAACCAGTATGTGAATAAGAAATTCAGCAATCAGTACAAAGCCACAATAGGAGCTGACTTTCTGACCAAGGAGGTGATGGTGGATGACAGGCTAGTCACAATG;MAPQ=60;MATEID=1646920_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_3_128502501_128527501_323C;SPAN=80010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:49 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:72 DR:0 LR:-211.3 LO:211.3);ALT=G[chr3:128525212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128526515	+	chr3	128532167	+	.	6	5	1647108_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=1647108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128527001_128552001_126C;SPAN=5652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:5 DR:6 LR:-15.67 LO:21.47);ALT=G[chr3:128532167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128853797	+	chr3	128859211	+	.	0	8	1648403_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1648403_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128845501_128870501_342C;SPAN=5414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:108 GQ:2.7 PL:[0.0, 2.7, 267.3] SR:8 DR:0 LR:2.852 LO:14.42);ALT=G[chr3:128859211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128859328	+	chr3	128864604	+	.	0	7	1648440_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1648440_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128845501_128870501_244C;SPAN=5276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:106 GQ:5.4 PL:[0.0, 5.4, 267.3] SR:7 DR:0 LR:5.611 LO:12.26);ALT=T[chr3:128864604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128864717	+	chr3	128875698	+	ATTCTGAATCTGAGCCACTTTTTTAGAGATCTCTCCAATGAT	0	25	1648520_1	62.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ATTCTGAATCTGAGCCACTTTTTTAGAGATCTCTCCAATGAT;MAPQ=60;MATEID=1648520_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_128870001_128895001_130C;SPAN=10981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:74 GQ:62.6 PL:[62.6, 0.0, 115.4] SR:25 DR:0 LR:-62.48 LO:63.39);ALT=C[chr3:128875698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128875765	+	chr3	128879815	+	TCACTTTTCCCTCTTCCAGCTGAGCCTGGCGAAATCTTGCTAAGGCCGTCATGGCCTTTTCTGCATTTCGGG	23	27	1648545_1	83.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TCACTTTTCCCTCTTCCAGCTGAGCCTGGCGAAATCTTGCTAAGGCCGTCATGGCCTTTTCTGCATTTCGGG;MAPQ=60;MATEID=1648545_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_128870001_128895001_194C;SPAN=4050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:94 GQ:83.6 PL:[83.6, 0.0, 143.0] SR:27 DR:23 LR:-83.47 LO:84.37);ALT=T[chr3:128879815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	128890617	+	chr3	128902619	+	.	255	26	1648624_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=1648624_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_128870001_128895001_315C;SPAN=12002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:258 DP:72 GQ:69.7 PL:[765.7, 69.7, 0.0] SR:26 DR:255 LR:-765.8 LO:765.8);ALT=T[chr3:128902619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	129115984	+	chr3	129117850	+	.	0	15	1649608_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1649608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_129115001_129140001_318C;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:115 GQ:18.5 PL:[18.5, 0.0, 259.4] SR:15 DR:0 LR:-18.36 LO:30.93);ALT=C[chr3:129117850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	129156794	+	chr3	129158573	+	.	0	8	1649580_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1649580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_129139501_129164501_243C;SPAN=1779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:115 GQ:4.5 PL:[0.0, 4.5, 287.1] SR:8 DR:0 LR:4.748 LO:14.2);ALT=C[chr3:129158573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	129763382	+	chr3	129806746	+	.	64	34	1652305_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=1652305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_129801001_129826001_158C;SPAN=43364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:39 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:34 DR:64 LR:-237.7 LO:237.7);ALT=C[chr3:129806746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	129886026	+	chr12	8460446	+	.	9	0	1653105_1	29.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=1653105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:129886026(+)-12:8460446(-)__3_129874501_129899501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:11 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:9 LR:-28.4 LO:28.4);ALT=G[chr12:8460446[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	130569773	+	chr3	130574722	+	.	0	7	1655025_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=1655025_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_130560501_130585501_219C;SPAN=4949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:98 GQ:3.3 PL:[0.0, 3.3, 244.2] SR:7 DR:0 LR:3.444 LO:12.5);ALT=G[chr3:130574722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140236164	+	chr3	130705716	+	.	17	23	2235525_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=AGTTTAGTTTAG;MAPQ=47;MATEID=2235525_2;MATENM=0;NM=11;NUMPARTS=2;SCTG=c_4_140213501_140238501_393C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:54 GQ:21.8 PL:[107.6, 0.0, 21.8] SR:23 DR:17 LR:-110.5 LO:110.5);ALT=]chr4:140236164]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	130717233	+	chr3	130718359	+	.	2	4	1655516_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1655516_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_130707501_130732501_207C;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:4 DR:2 LR:5.711 LO:8.577);ALT=G[chr3:130718359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	131220589	+	chr3	131221623	+	.	14	0	1657083_1	16.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=1657083_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:131220589(+)-3:131221623(-)__3_131197501_131222501D;SPAN=1034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:110 GQ:16.4 PL:[16.4, 0.0, 250.7] SR:0 DR:14 LR:-16.41 LO:28.71);ALT=A[chr3:131221623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50169357	+	chr3	131245418	+	.	11	0	6849925_1	25.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6849925_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:131245418(-)-19:50169357(+)__19_50151501_50176501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:42 GQ:25.1 PL:[25.1, 0.0, 74.6] SR:0 DR:11 LR:-24.93 LO:26.41);ALT=]chr19:50169357]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	140660937	+	chr3	140675368	+	.	10	23	1689142_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1689142_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_140654501_140679501_233C;SPAN=14431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:108 GQ:63.2 PL:[63.2, 0.0, 198.5] SR:23 DR:10 LR:-63.17 LO:67.09);ALT=G[chr3:140675368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	140675534	+	chr3	140678305	+	.	2	12	1689200_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1689200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_140654501_140679501_127C;SPAN=2771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:109 GQ:13.4 PL:[13.4, 0.0, 251.0] SR:12 DR:2 LR:-13.38 LO:26.26);ALT=G[chr3:140678305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	140692847	+	chr3	140695101	+	.	2	5	1689250_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1689250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_140679001_140704001_375C;SPAN=2254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:99 GQ:6.9 PL:[0.0, 6.9, 254.1] SR:5 DR:2 LR:7.016 LO:10.28);ALT=G[chr3:140695101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	141385018	-	chr19	30401093	+	.	4	11	1691702_1	39.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=AAGGAAGGAAGGAAGGAAGGAAGGAAGGAAGGA;MAPQ=60;MATEID=1691702_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_141365001_141390001_186C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:6 GQ:3.6 PL:[39.6, 3.6, 0.0] SR:11 DR:4 LR:-39.61 LO:39.61);ALT=[chr19:30401093[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	141457264	+	chr3	141463999	+	.	18	0	1692209_1	42.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=1692209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:141457264(+)-3:141463999(-)__3_141463001_141488001D;SPAN=6735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:63 GQ:42.5 PL:[42.5, 0.0, 108.5] SR:0 DR:18 LR:-42.35 LO:44.03);ALT=C[chr3:141463999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	141622591	+	chr3	141626007	+	.	2	5	1692648_1	0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1692648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_141610001_141635001_393C;SPAN=3416;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:110 GQ:9.9 PL:[0.0, 9.9, 287.1] SR:5 DR:2 LR:9.996 LO:9.995);ALT=G[chr3:141626007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	141713984	+	chr3	141724283	+	.	0	23	1693326_1	45.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1693326_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_141708001_141733001_327C;SPAN=10299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:112 GQ:45.8 PL:[45.8, 0.0, 224.0] SR:23 DR:0 LR:-45.58 LO:52.42);ALT=C[chr3:141724283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	141714032	+	chr3	141747418	+	.	24	0	1693328_1	62.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1693328_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:141714032(+)-3:141747418(-)__3_141708001_141733001D;SPAN=33386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:60 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:0 DR:24 LR:-62.97 LO:63.12);ALT=G[chr3:141747418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	141724441	+	chr3	141747419	+	.	15	0	1693361_1	37.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1693361_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:141724441(+)-3:141747419(-)__3_141708001_141733001D;SPAN=22978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:45 GQ:37.4 PL:[37.4, 0.0, 70.4] SR:0 DR:15 LR:-37.32 LO:37.92);ALT=T[chr3:141747419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142151739	+	chr3	142166712	+	.	15	7	1694621_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGA;MAPQ=60;MATEID=1694621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142149001_142174001_94C;SPAN=14973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:109 GQ:33.2 PL:[33.2, 0.0, 231.2] SR:7 DR:15 LR:-33.19 LO:41.79);ALT=A[chr3:142166712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142285139	+	chr3	142297504	+	.	8	0	1695173_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1695173_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:142285139(+)-3:142297504(-)__3_142296001_142321001D;SPAN=12365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.443 LO:16.0);ALT=A[chr3:142297504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142286998	+	chr3	142297488	+	.	2	3	1695135_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1695135_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142271501_142296501_1C;SPAN=10490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:32 GQ:8 PL:[8.0, 0.0, 67.4] SR:3 DR:2 LR:-7.835 LO:10.74);ALT=T[chr3:142297488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142720539	+	chr3	142731061	+	.	24	0	1696514_1	50.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1696514_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:142720539(+)-3:142731061(-)__3_142712501_142737501D;SPAN=10522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:107 GQ:50.3 PL:[50.3, 0.0, 208.7] SR:0 DR:24 LR:-50.24 LO:55.75);ALT=A[chr3:142731061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142731195	+	chr3	142733153	+	.	0	20	1696560_1	41.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1696560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142712501_142737501_36C;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:91 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:20 DR:0 LR:-41.37 LO:46.26);ALT=A[chr3:142733153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142733252	+	chr3	142735097	+	.	0	14	1696566_1	18.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1696566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142712501_142737501_170C;SPAN=1845;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:14 DR:0 LR:-18.58 LO:29.2);ALT=G[chr3:142735097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142754947	+	chr3	142756019	+	.	4	5	1696386_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1696386_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142737001_142762001_316C;SPAN=1072;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:5 DR:4 LR:-1.212 LO:14.96);ALT=G[chr3:142756019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142772637	+	chr3	142773783	+	.	7	2	1696657_1	0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1696657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142761501_142786501_140C;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:114 GQ:4.2 PL:[0.0, 4.2, 283.8] SR:2 DR:7 LR:4.477 LO:14.23);ALT=G[chr3:142773783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142772650	+	chr3	142775151	+	.	8	0	1696658_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1696658_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:142772650(+)-3:142775151(-)__3_142761501_142786501D;SPAN=2501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=C[chr3:142775151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	142773961	+	chr3	142775152	+	.	0	6	1696662_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1696662_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_142761501_142786501_361C;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:114 GQ:10.8 PL:[0.0, 10.8, 297.0] SR:6 DR:0 LR:11.08 LO:9.9);ALT=G[chr3:142775152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	143219592	+	chr3	143221217	+	.	40	35	1698113_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATGTTA;MAPQ=60;MATEID=1698113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_143202501_143227501_296C;SPAN=1625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:56 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:35 DR:40 LR:-181.5 LO:181.5);ALT=A[chr3:143221217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	84250213	+	chr3	143592939	+	.	12	0	1699626_1	23.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1699626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:143592939(-)-13:84250213(+)__3_143570001_143595001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:0 DR:12 LR:-23.36 LO:27.2);ALT=]chr13:84250213]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	148281440	+	chr3	148285420	+	.	27	26	1713272_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GTCCTG;MAPQ=60;MATEID=1713272_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148274001_148299001_210C;SPAN=3980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:61 GQ:3.5 PL:[142.1, 0.0, 3.5] SR:26 DR:27 LR:-149.4 LO:149.4);ALT=G[chr3:148285420[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	148709431	+	chr3	148714086	+	.	9	0	1714639_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1714639_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:148709431(+)-3:148714086(-)__3_148690501_148715501D;SPAN=4655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:0 DR:9 LR:-3.971 LO:17.23);ALT=A[chr3:148714086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	148709434	+	chr3	148711927	+	.	32	12	1714640_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1714640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148690501_148715501_306C;SPAN=2493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:112 GQ:92 PL:[92.0, 0.0, 177.8] SR:12 DR:32 LR:-91.79 LO:93.37);ALT=G[chr3:148711927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	148712064	+	chr3	148714087	+	.	0	26	1714648_1	55.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1714648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148690501_148715501_343C;SPAN=2023;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:113 GQ:55.4 PL:[55.4, 0.0, 217.1] SR:26 DR:0 LR:-55.21 LO:60.73);ALT=G[chr3:148714087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	148802678	+	chr3	148804103	+	.	0	6	1714984_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1714984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_148788501_148813501_243C;SPAN=1425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:85 GQ:3 PL:[0.0, 3.0, 211.2] SR:6 DR:0 LR:3.223 LO:10.69);ALT=T[chr3:148804103[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	149468639	+	chr3	149469996	+	ATGAGCTTTGAGCTCTCAGTGAGGAGATACGTTAATCCTTCCACACCATGCTGGACAGTGTCACTACTCACATTGAGTTTT	0	14	1717421_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATGAGCTTTGAGCTCTCAGTGAGGAGATACGTTAATCCTTCCACACCATGCTGGACAGTGTCACTACTCACATTGAGTTTT;MAPQ=60;MATEID=1717421_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_149450001_149475001_410C;SPAN=1357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:112 GQ:16.1 PL:[16.1, 0.0, 253.7] SR:14 DR:0 LR:-15.87 LO:28.59);ALT=C[chr3:149469996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	149531142	+	chr3	149563796	+	.	2	2	1717632_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1717632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_149548001_149573001_317C;SPAN=32654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:54 GQ:1.2 PL:[0.0, 1.2, 132.0] SR:2 DR:2 LR:1.426 LO:7.211);ALT=T[chr3:149563796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150262286	+	chr3	150263490	+	.	0	54	1720097_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1720097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_150258501_150283501_127C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:126 GQ:99 PL:[144.2, 0.0, 160.7] SR:54 DR:0 LR:-144.1 LO:144.2);ALT=C[chr3:150263490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150262316	+	chr3	150263838	+	.	9	0	1720098_1	1.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1720098_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150262316(+)-3:150263838(-)__3_150258501_150283501D;SPAN=1522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:106 GQ:1.1 PL:[1.1, 0.0, 255.2] SR:0 DR:9 LR:-0.991 LO:16.78);ALT=A[chr3:150263838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150264663	+	chr3	150281301	+	.	8	0	1720104_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1720104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150264663(+)-3:150281301(-)__3_150258501_150283501D;SPAN=16638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:0 DR:8 LR:-3.109 LO:15.25);ALT=C[chr3:150281301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150264663	+	chr3	150276172	+	.	16	0	1720103_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1720103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150264663(+)-3:150276172(-)__3_150258501_150283501D;SPAN=11509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:95 GQ:27.2 PL:[27.2, 0.0, 202.1] SR:0 DR:16 LR:-27.08 LO:34.93);ALT=C[chr3:150276172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150264665	+	chr3	150280328	+	.	45	0	1720105_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1720105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150264665(+)-3:150280328(-)__3_150258501_150283501D;SPAN=15663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:93 GQ:99 PL:[123.5, 0.0, 100.4] SR:0 DR:45 LR:-123.5 LO:123.5);ALT=T[chr3:150280328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150290316	+	chr3	150293435	+	.	0	7	1720212_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1720212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_150283001_150308001_229C;SPAN=3119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:93 GQ:1.8 PL:[0.0, 1.8, 227.7] SR:7 DR:0 LR:2.089 LO:12.67);ALT=G[chr3:150293435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	150321202	+	chr9	6278666	+	.	9	0	4131708_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4131708_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150321202(+)-9:6278666(-)__9_6272001_6297001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=A[chr9:6278666[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	150321204	+	chr3	150340169	+	.	28	0	1720509_1	79.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1720509_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:150321204(+)-3:150340169(-)__3_150332001_150357001D;SPAN=18965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:49 GQ:39.5 PL:[79.1, 0.0, 39.5] SR:0 DR:28 LR:-79.86 LO:79.86);ALT=G[chr3:150340169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	151148544	-	chr5	39787751	+	.	22	47	2458236_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=2458236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_39763501_39788501_137C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:42 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:47 DR:22 LR:-184.8 LO:184.8);ALT=[chr5:39787751[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	151591540	+	chr3	151598345	+	.	24	0	1724661_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1724661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:151591540(+)-3:151598345(-)__3_151581501_151606501D;SPAN=6805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:98 GQ:52.7 PL:[52.7, 0.0, 184.7] SR:0 DR:24 LR:-52.67 LO:56.81);ALT=C[chr3:151598345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	151962215	+	chr3	152017192	+	TAAAGCATAG	54	7	1726448_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TAAAGCATAG;MAPQ=60;MATEID=1726448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_151998001_152023001_33C;SPAN=54977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:80 GQ:24.5 PL:[169.7, 0.0, 24.5] SR:7 DR:54 LR:-176.0 LO:176.0);ALT=T[chr3:152017192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	152018156	+	chr3	152019708	+	.	9	5	1726529_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1726529_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_151998001_152023001_349C;SPAN=1552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:118 GQ:11 PL:[11.0, 0.0, 275.0] SR:5 DR:9 LR:-10.94 LO:25.79);ALT=A[chr3:152019708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	152311738	+	chr3	152313156	+	.	75	42	1727140_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAGGTCACTGTTT;MAPQ=60;MATEID=1727140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_152292001_152317001_39C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:96 DP:235 GQ:99 PL:[253.4, 0.0, 316.1] SR:42 DR:75 LR:-253.2 LO:253.6);ALT=T[chr3:152313156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	152810869	+	chr7	87740201	-	.	12	0	3440945_1	30.0	.	DISC_MAPQ=10;EVDNC=DSCRD;IMPRECISE;MAPQ=10;MATEID=3440945_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:152810869(+)-7:87740201(+)__7_87734501_87759501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:0 DR:12 LR:-30.4 LO:30.71);ALT=G]chr7:87740201];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	153153198	-	chr3	153154605	+	.	10	0	1730455_1	11.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=1730455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:153153198(-)-3:153154605(-)__3_153149501_153174501D;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.34 LO:20.42);ALT=[chr3:153154605[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	154033954	+	chr3	154041963	+	.	0	9	1732959_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1732959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_154031501_154056501_339C;SPAN=8009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:9 DR:0 LR:-1.533 LO:16.86);ALT=T[chr3:154041963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101730148	+	chr3	155027227	+	.	17	0	1735932_1	45.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1735932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:155027227(-)-8:101730148(+)__3_155011501_155036501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:40 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:0 DR:17 LR:-45.28 LO:45.31);ALT=]chr8:101730148]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	155215996	-	chr3	155217435	+	.	8	0	1736814_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1736814_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:155215996(-)-3:155217435(-)__3_155207501_155232501D;SPAN=1439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=[chr3:155217435[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	155290513	-	chr3	155292821	+	.	8	0	1736443_1	0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=1736443_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:155290513(-)-3:155292821(-)__3_155281001_155306001D;SPAN=2308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=[chr3:155292821[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	155588686	+	chr3	155611305	+	.	0	27	1737888_1	75.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1737888_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_155575001_155600001_228C;SPAN=22619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:52 GQ:48.8 PL:[75.2, 0.0, 48.8] SR:27 DR:0 LR:-75.28 LO:75.28);ALT=G[chr3:155611305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	155633982	+	chr3	155637020	+	.	2	3	1737970_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=1737970_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGAGGA;SCTG=c_3_155624001_155649001_125C;SPAN=3038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:102 GQ:14.2 PL:[0.0, 14.2, 210.6] SR:3 DR:2 LR:14.62 LO:4.667);ALT=G[chr3:155637020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131451934	+	chr3	155705203	+	.	27	11	1738500_1	89.0	.	DISC_MAPQ=4;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1738500_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_3_155697501_155722501_174C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:74 GQ:89 PL:[89.0, 0.0, 89.0] SR:11 DR:27 LR:-88.89 LO:88.89);ALT=]chr9:131451934]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	156261058	+	chr3	156262096	+	.	4	21	1740042_1	52.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=G;MAPQ=15;MATEID=1740042_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_156261001_156286001_214C;SPAN=1038;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:99 GQ:52.4 PL:[52.4, 0.0, 187.7] SR:21 DR:4 LR:-52.4 LO:56.69);ALT=C[chr3:156262096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	156271570	+	chr3	156272745	+	.	29	54	1740076_1	99.0	.	DISC_MAPQ=29;EVDNC=ASDIS;HOMSEQ=C;MAPQ=18;MATEID=1740076_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_156261001_156286001_30C;SPAN=1175;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:127 GQ:81.2 PL:[226.4, 0.0, 81.2] SR:54 DR:29 LR:-230.1 LO:230.1);ALT=C[chr3:156272745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	156392586	+	chr3	156395444	+	.	17	12	1740487_1	41.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1740487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_156383501_156408501_176C;SPAN=2858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:93 GQ:41 PL:[41.0, 0.0, 182.9] SR:12 DR:17 LR:-40.82 LO:46.04);ALT=G[chr3:156395444[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	157828000	+	chr3	157839890	+	.	30	7	1745094_1	94.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1745094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_157829001_157854001_44C;SPAN=11890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:55 GQ:38 PL:[94.1, 0.0, 38.0] SR:7 DR:30 LR:-95.25 LO:95.25);ALT=G[chr3:157839890[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	157840087	+	chr3	157841653	+	.	4	23	1745145_1	55.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1745145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_157829001_157854001_372C;SPAN=1566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:89 GQ:55.1 PL:[55.1, 0.0, 160.7] SR:23 DR:4 LR:-55.11 LO:57.99);ALT=G[chr3:157841653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	157841782	+	chr3	157920859	+	.	0	18	1745148_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=1745148_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_157829001_157854001_65C;SPAN=79077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:35 GQ:33.5 PL:[50.0, 0.0, 33.5] SR:18 DR:0 LR:-50.08 LO:50.08);ALT=T[chr3:157920859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	158350740	+	chr3	158351912	+	.	60	35	1746939_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1746939_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_158343501_158368501_258C;SPAN=1172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:68 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:35 DR:60 LR:-217.9 LO:217.9);ALT=C[chr3:158351912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	158520016	+	chr3	158522106	+	.	22	0	1747155_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1747155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:158520016(+)-3:158522106(-)__3_158515001_158540001D;SPAN=2090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:127 GQ:38.3 PL:[38.3, 0.0, 269.3] SR:0 DR:22 LR:-38.21 LO:48.32);ALT=C[chr3:158522106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	158520134	+	chr3	158523150	+	.	21	0	1747160_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1747160_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:158520134(+)-3:158523150(-)__3_158515001_158540001D;SPAN=3016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:116 GQ:38 PL:[38.0, 0.0, 242.6] SR:0 DR:21 LR:-37.89 LO:46.57);ALT=C[chr3:158523150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	159431108	+	chr21	31260473	-	.	8	0	7153285_1	23.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7153285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:159431108(+)-21:31260473(+)__21_31237501_31262501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:11 GQ:0.5 PL:[23.6, 0.0, 0.5] SR:0 DR:8 LR:-24.3 LO:24.3);ALT=T]chr21:31260473];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	159558004	+	chr3	159583950	+	.	18	22	1750309_1	87.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1750309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_159544001_159569001_171C;SPAN=25946;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:68 GQ:77.3 PL:[87.2, 0.0, 77.3] SR:22 DR:18 LR:-87.24 LO:87.24);ALT=G[chr3:159583950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	160156979	+	chr3	160167470	+	.	8	0	1752411_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1752411_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:160156979(+)-3:160167470(-)__3_160156501_160181501D;SPAN=10491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:0 DR:8 LR:3.123 LO:14.39);ALT=C[chr3:160167470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	160170211	-	chr11	62389375	+	.	14	0	1752453_1	32.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=1752453_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:160170211(-)-11:62389375(-)__3_160156501_160181501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:51 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:0 DR:14 LR:-32.4 LO:33.96);ALT=[chr11:62389375[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	160939233	+	chr3	160942717	+	.	11	0	1754793_1	18.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1754793_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:160939233(+)-3:160942717(-)__3_160916001_160941001D;SPAN=3484;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:0 DR:11 LR:-18.43 LO:23.96);ALT=G[chr3:160942717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	160939845	+	chr3	160942718	+	.	2	6	1754796_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1754796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_160916001_160941001_84C;SPAN=2873;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:41 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:6 DR:2 LR:-12.0 LO:15.33);ALT=T[chr3:160942718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	163919285	+	chr10	36760446	+	.	50	39	4574086_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=4574086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_36750001_36775001_210C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:38 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:39 DR:50 LR:-201.3 LO:201.3);ALT=A[chr10:36760446[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	169684647	+	chr3	169693393	+	.	15	12	1781868_1	72.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=1781868_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_169687001_169712001_353C;SPAN=8746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:48 GQ:43.1 PL:[72.8, 0.0, 43.1] SR:12 DR:15 LR:-73.21 LO:73.21);ALT=G[chr3:169693393[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	169684685	+	chr3	169694728	+	.	35	0	1781870_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1781870_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:169684685(+)-3:169694728(-)__3_169687001_169712001D;SPAN=10043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:57 GQ:37.4 PL:[100.1, 0.0, 37.4] SR:0 DR:35 LR:-101.6 LO:101.6);ALT=C[chr3:169694728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	169693504	+	chr3	169694733	+	.	0	35	1781889_1	85.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1781889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_169687001_169712001_227C;SPAN=1229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:110 GQ:85.7 PL:[85.7, 0.0, 181.4] SR:35 DR:0 LR:-85.73 LO:87.61);ALT=G[chr3:169694733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	169694840	+	chr3	169700493	+	.	0	34	1781892_1	79.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=1781892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_169687001_169712001_528C;SPAN=5653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:123 GQ:79.1 PL:[79.1, 0.0, 217.7] SR:34 DR:0 LR:-78.91 LO:82.59);ALT=G[chr3:169700493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	146184521	+	chr3	170395035	+	.	2	6	4121126_1	10.0	.	DISC_MAPQ=1;EVDNC=TSI_L;HOMSEQ=GGTTGGGGTACTTGCCCCTCCCCTAGAAAAGCAGGACTTGCC;MAPQ=60;MATEID=4121126_2;MATENM=0;NM=5;NUMPARTS=3;REPSEQ=GG;SCTG=c_8_146167001_146192001_268C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:6 DR:2 LR:-10.42 LO:16.64);ALT=]chr8:146184521]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	170395175	+	chr8	146184452	+	TCCCAGAAAAGTG	11	17	4121127_1	72.0	.	DISC_MAPQ=0;EVDNC=TSI_L;HOMSEQ=GGTTGGGGTACTTGCCCCTCCCCTAGAAAAGCAGGACTTGCC;INSERTION=TCCCAGAAAAGTG;MAPQ=60;MATEID=4121127_2;MATENM=1;NM=5;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_8_146167001_146192001_268C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:50 GQ:49.1 PL:[72.2, 0.0, 49.1] SR:17 DR:11 LR:-72.52 LO:72.52);ALT=C[chr8:146184452[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	170584319	+	chr3	170585800	+	.	0	163	1784520_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCTTTTA;MAPQ=60;MATEID=1784520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_170569001_170594001_386C;SPAN=1481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:163 DP:105 GQ:43.9 PL:[481.9, 43.9, 0.0] SR:163 DR:0 LR:-481.9 LO:481.9);ALT=A[chr3:170585800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	170584372	+	chr3	170587947	+	.	30	0	1784521_1	60.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1784521_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:170584372(+)-3:170587947(-)__3_170569001_170594001D;SPAN=3575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:142 GQ:60.8 PL:[60.8, 0.0, 281.9] SR:0 DR:30 LR:-60.56 LO:68.8);ALT=T[chr3:170587947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	170586204	+	chr3	170587947	+	.	54	0	1784532_1	99.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1784532_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:170586204(+)-3:170587947(-)__3_170569001_170594001D;SPAN=1743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:149 GQ:99 PL:[137.9, 0.0, 223.7] SR:0 DR:54 LR:-137.9 LO:139.0);ALT=T[chr3:170587947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	170587947	-	chr4	55087355	+	.	8	0	1971635_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1971635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:170587947(-)-4:55087355(-)__4_55076001_55101001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=[chr4:55087355[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	179065603	+	chr3	179066639	+	.	9	0	1812182_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1812182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:179065603(+)-3:179066639(-)__3_179046001_179071001D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:0 DR:9 LR:-1.533 LO:16.86);ALT=G[chr3:179066639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179137295	+	chr3	179143931	+	GAACAAGCGTTGCATCATTACATGCTTTCCGAGCAT	0	9	1812464_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTGAA;INSERTION=GAACAAGCGTTGCATCATTACATGCTTTCCGAGCAT;MAPQ=60;MATEID=1812464_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_179119501_179144501_367C;SPAN=6636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-7.764 LO:17.89);ALT=T[chr3:179143931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179137344	+	chr3	179169138	+	.	8	0	1812591_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1812591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:179137344(+)-3:179169138(-)__3_179168501_179193501D;SPAN=31794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=G[chr3:179169138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179144033	+	chr3	179169134	+	.	8	7	1812592_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=1812592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179168501_179193501_248C;SPAN=25101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:34 GQ:23.9 PL:[23.9, 0.0, 56.9] SR:7 DR:8 LR:-23.8 LO:24.62);ALT=G[chr3:179169134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179306785	+	chr3	179310432	+	.	0	26	1813191_1	53.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1813191_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179291001_179316001_287C;SPAN=3647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:120 GQ:53.3 PL:[53.3, 0.0, 238.1] SR:26 DR:0 LR:-53.32 LO:59.95);ALT=T[chr3:179310432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179310528	+	chr3	179311552	+	.	0	13	1813212_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1813212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179291001_179316001_152C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:119 GQ:10.7 PL:[10.7, 0.0, 278.0] SR:13 DR:0 LR:-10.67 LO:25.74);ALT=C[chr3:179311552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179316560	+	chr3	179320439	+	AAAGTTTGTGTAAATCTTCATTACTTTTGTTCCTTAGTTGCTGACAGGTCCATGCTGCT	0	30	1813228_1	68.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AAAGTTTGTGTAAATCTTCATTACTTTTGTTCCTTAGTTGCTGACAGGTCCATGCTGCT;MAPQ=60;MATEID=1813228_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_179315501_179340501_247C;SPAN=3879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:114 GQ:68.3 PL:[68.3, 0.0, 206.9] SR:30 DR:0 LR:-68.15 LO:72.11);ALT=C[chr3:179320439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179319621	+	chr3	179322365	+	.	8	0	1813242_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1813242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:179319621(+)-3:179322365(-)__3_179315501_179340501D;SPAN=2744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:113 GQ:3.9 PL:[0.0, 3.9, 280.5] SR:0 DR:8 LR:4.207 LO:14.26);ALT=G[chr3:179322365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179320586	+	chr3	179322313	+	.	39	9	1813245_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1813245_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179315501_179340501_263C;SPAN=1727;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:109 GQ:99 PL:[102.5, 0.0, 161.9] SR:9 DR:39 LR:-102.5 LO:103.2);ALT=C[chr3:179322313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179322727	+	chr3	179332758	+	.	58	44	1813256_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=1813256_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GTCGTC;SCTG=c_3_179315501_179340501_325C;SPAN=10031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:103 DP:136 GQ:12.8 PL:[231.3, 0.0, 12.8] SR:44 DR:58 LR:-244.7 LO:244.7);ALT=G[chr3:179332758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179322729	+	chr3	179334770	+	.	12	7	1813258_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=1813258_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_3_179315501_179340501_321C;SPAN=12041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:126 GQ:18.8 PL:[18.8, 0.0, 286.1] SR:7 DR:12 LR:-18.68 LO:32.79);ALT=T[chr3:179334770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179322729	+	chr3	179336201	+	CAAGCTGAACTAGCAGAAATTCCAGAAGGCTATGTCCCAGAACACTGGGAATATTATA	6	20	1813259_1	46.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAAGCTGAACTAGCAGAAATTCCAGAAGGCTATGTCCCAGAACACTGGGAATATTATA;MAPQ=60;MATEID=1813259_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_179315501_179340501_321C;SPAN=13472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:135 GQ:46.1 PL:[46.1, 0.0, 280.4] SR:20 DR:6 LR:-45.95 LO:55.72);ALT=T[chr3:179336201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179334832	+	chr3	179336201	+	.	0	23	1813301_1	46.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1813301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179315501_179340501_445C;SPAN=1369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:109 GQ:46.4 PL:[46.4, 0.0, 218.0] SR:23 DR:0 LR:-46.39 LO:52.73);ALT=G[chr3:179336201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	179336310	+	chr3	179341707	+	.	10	14	1813334_1	60.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1813334_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_179340001_179365001_22C;SPAN=5397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:46 GQ:50.3 PL:[60.2, 0.0, 50.3] SR:14 DR:10 LR:-60.19 LO:60.19);ALT=G[chr3:179341707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	180630553	+	chr3	180651119	+	.	15	0	1817635_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1817635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:180630553(+)-3:180651119(-)__3_180614001_180639001D;SPAN=20566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:56 GQ:34.4 PL:[34.4, 0.0, 100.4] SR:0 DR:15 LR:-34.34 LO:36.19);ALT=T[chr3:180651119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	180630560	+	chr3	180632453	+	.	29	0	1817636_1	65.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1817636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:180630560(+)-3:180632453(-)__3_180614001_180639001D;SPAN=1893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:110 GQ:65.9 PL:[65.9, 0.0, 201.2] SR:0 DR:29 LR:-65.93 LO:69.74);ALT=G[chr3:180632453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	180707414	-	chr14	45759196	+	.	36	0	5726304_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5726304_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:180707414(-)-14:45759196(-)__14_45741501_45766501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:51 GQ:16.1 PL:[105.2, 0.0, 16.1] SR:0 DR:36 LR:-108.4 LO:108.4);ALT=[chr14:45759196[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	182511575	+	chr3	182538047	+	.	5	7	1823674_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1823674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_182525001_182550001_17C;SPAN=26472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:62 GQ:13.1 PL:[13.1, 0.0, 135.2] SR:7 DR:5 LR:-12.91 LO:19.01);ALT=G[chr3:182538047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	182810337	+	chr3	182817139	+	GGCTGTTGTGTACTTCATGGTTCTTTGCCTCCACACCCATGT	0	12	1824767_1	2.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GGCTGTTGTGTACTTCATGGTTCTTTGCCTCCACACCCATGT;MAPQ=60;MATEID=1824767_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_182794501_182819501_25C;SPAN=6802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:136 GQ:2.9 PL:[2.9, 0.0, 326.3] SR:12 DR:0 LR:-2.766 LO:22.58);ALT=T[chr3:182817139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183415781	+	chr3	183432931	+	.	3	3	1827139_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1827139_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183407001_183432001_203C;SPAN=17150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:29 GQ:8.6 PL:[8.6, 0.0, 61.4] SR:3 DR:3 LR:-8.648 LO:10.97);ALT=G[chr3:183432931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183547497	+	chr3	183551280	+	.	0	11	1827590_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1827590_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183529501_183554501_2C;SPAN=3783;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:129 GQ:1.4 PL:[1.4, 0.0, 311.6] SR:11 DR:0 LR:-1.362 LO:20.53);ALT=T[chr3:183551280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183585850	+	chr3	183595938	+	.	6	2	1828388_1	0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=1828388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183578501_183603501_268C;SPAN=10088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:126 GQ:14.1 PL:[0.0, 14.1, 333.3] SR:2 DR:6 LR:14.33 LO:9.634);ALT=T[chr3:183595938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183585850	+	chr3	183602508	+	.	52	27	1828389_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=1828389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183578501_183603501_240C;SPAN=16658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:130 GQ:99 PL:[176.0, 0.0, 139.7] SR:27 DR:52 LR:-176.3 LO:176.3);ALT=T[chr3:183602508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183732233	+	chr3	183735616	+	.	8	0	1828280_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1828280_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:183732233(+)-3:183735616(-)__3_183725501_183750501D;SPAN=3383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=T[chr3:183735616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183853370	+	chr3	183854399	+	.	0	14	1828961_1	12.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=1828961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183848001_183873001_346C;SPAN=1029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:126 GQ:12.2 PL:[12.2, 0.0, 292.7] SR:14 DR:0 LR:-12.08 LO:27.83);ALT=T[chr3:183854399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183892749	+	chr3	183894737	+	.	60	13	1828920_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=1828920_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183872501_183897501_12C;SPAN=1988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:136 GQ:99 PL:[177.8, 0.0, 151.4] SR:13 DR:60 LR:-177.8 LO:177.8);ALT=T[chr3:183894737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183892781	+	chr3	183896641	+	.	60	0	1828921_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1828921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:183892781(+)-3:183896641(-)__3_183872501_183897501D;SPAN=3860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:128 GQ:99 PL:[163.4, 0.0, 146.9] SR:0 DR:60 LR:-163.4 LO:163.4);ALT=A[chr3:183896641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183894856	+	chr3	183896644	+	.	0	81	1828926_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=1828926_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183872501_183897501_92C;SPAN=1788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:161 GQ:99 PL:[224.0, 0.0, 164.6] SR:81 DR:0 LR:-224.2 LO:224.2);ALT=G[chr3:183896644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183896910	+	chr3	183897956	+	.	9	13	1828931_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1828931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183872501_183897501_261C;SPAN=1046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:13 DR:9 LR:-31.91 LO:35.06);ALT=G[chr3:183897956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183963602	+	chr3	183966570	+	.	25	3	1829196_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1829196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_183946001_183971001_403C;SPAN=2968;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:113 GQ:52.1 PL:[52.1, 0.0, 220.4] SR:3 DR:25 LR:-51.91 LO:57.9);ALT=T[chr3:183966570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	183967680	+	chr3	183975259	+	.	0	10	1829375_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=1829375_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_183970501_183995501_69C;SPAN=7579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=T[chr3:183975259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184034006	+	chr3	184035106	+	.	0	7	1829634_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1829634_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_184019501_184044501_310C;SPAN=1100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:104 GQ:4.8 PL:[0.0, 4.8, 260.7] SR:7 DR:0 LR:5.069 LO:12.32);ALT=G[chr3:184035106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184081353	+	chr3	184082752	+	.	43	20	1829901_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1829901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_184068501_184093501_123C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:118 GQ:99 PL:[133.1, 0.0, 152.9] SR:20 DR:43 LR:-133.1 LO:133.2);ALT=G[chr3:184082752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184083015	+	chr3	184085965	+	GCTGACCAGTTTGAGTATGTAATGTATGGAAAAGTGTACAGGATTGAGGGAGATGAAACTTCTACTGAAGCAGCAACACGCCT	0	17	1829911_1	28.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=GCTGACCAGTTTGAGTATGTAATGTATGGAAAAGTGTACAGGATTGAGGGAGATGAAACTTCTACTGAAGCAGCAACACGCCT;MAPQ=60;MATEID=1829911_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_184068501_184093501_463C;SPAN=2950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:102 GQ:28.7 PL:[28.7, 0.0, 216.8] SR:17 DR:0 LR:-28.48 LO:37.03);ALT=G[chr3:184085965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184084588	+	chr3	184085965	+	.	2	7	1829922_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=1829922_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_184068501_184093501_463C;SPAN=1377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:7 DR:2 LR:0.6845 LO:14.7);ALT=T[chr3:184085965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	184264648	+	chr3	184265715	-	.	9	0	1830709_1	15.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1830709_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:184264648(+)-3:184265715(+)__3_184240001_184265001D;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:0 DR:9 LR:-15.35 LO:19.68);ALT=G]chr3:184265715];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	185000867	+	chr3	185009397	+	.	18	0	1833303_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1833303_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185000867(+)-3:185009397(-)__3_184999501_185024501D;SPAN=8530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:134 GQ:23.3 PL:[23.3, 0.0, 300.5] SR:0 DR:18 LR:-23.11 LO:37.37);ALT=T[chr3:185009397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185258342	-	chr3	185259354	+	.	8	0	1834339_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=1834339_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185258342(-)-3:185259354(-)__3_185244501_185269501D;SPAN=1012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr3:185259354[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	185304302	+	chr3	185307899	+	.	5	4	1834622_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=1834622_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185293501_185318501_242C;SPAN=3597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:112 GQ:13.5 PL:[0.0, 13.5, 297.0] SR:4 DR:5 LR:13.84 LO:7.886);ALT=G[chr3:185307899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185404980	+	chr3	185407142	+	.	0	16	1835100_1	25.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1835100_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185391501_185416501_245C;SPAN=2162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:102 GQ:25.4 PL:[25.4, 0.0, 220.1] SR:16 DR:0 LR:-25.18 LO:34.39);ALT=C[chr3:185407142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185709137	+	chr3	185628707	+	.	9	0	1836298_1	18.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1836298_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185628707(-)-3:185709137(+)__3_185685501_185710501D;SPAN=80430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=]chr3:185709137]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	185635526	+	chr3	185637224	+	.	10	0	1836032_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1836032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185635526(+)-3:185637224(-)__3_185612001_185637001D;SPAN=1698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=G[chr3:185637224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185636233	+	chr3	185638892	+	TCTGATCCCTGTCTTGGGCAGCTCTCCATCCTCCTCCTCCTCCACCTCCTCCT	6	19	1836037_1	56.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=CTGT;INSERTION=TCTGATCCCTGTCTTGGGCAGCTCTCCATCCTCCTCCTCCTCCACCTCCTCCT;MAPQ=60;MATEID=1836037_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_185612001_185637001_35C;SPAN=2659;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:61 GQ:56.3 PL:[56.3, 0.0, 89.3] SR:19 DR:6 LR:-56.1 LO:56.57);ALT=A[chr3:185638892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185639020	+	chr3	185641582	+	.	12	0	1836198_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1836198_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185639020(+)-3:185641582(-)__3_185636501_185661501D;SPAN=2562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:136 GQ:2.9 PL:[2.9, 0.0, 326.3] SR:0 DR:12 LR:-2.766 LO:22.58);ALT=A[chr3:185641582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185641773	+	chr3	185643251	+	.	14	11	1836208_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1836208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185636501_185661501_68C;SPAN=1478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:127 GQ:41.6 PL:[41.6, 0.0, 266.0] SR:11 DR:14 LR:-41.52 LO:51.01);ALT=C[chr3:185643251[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185643449	+	chr3	185649363	+	.	17	0	1836216_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1836216_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:185643449(+)-3:185649363(-)__3_185636501_185661501D;SPAN=5914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:97 GQ:29.9 PL:[29.9, 0.0, 204.8] SR:0 DR:17 LR:-29.84 LO:37.44);ALT=A[chr3:185649363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185644522	+	chr3	185649364	+	.	28	11	1836223_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1836223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185636501_185661501_170C;SPAN=4842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:113 GQ:85.1 PL:[85.1, 0.0, 187.4] SR:11 DR:28 LR:-84.92 LO:87.11);ALT=C[chr3:185649364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185644523	+	chr3	185655612	+	.	24	14	1836224_1	52.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1836224_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185636501_185661501_322C;SPAN=11089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:161 GQ:52.4 PL:[52.4, 0.0, 336.2] SR:14 DR:24 LR:-52.11 LO:64.25);ALT=C[chr3:185655612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	185649641	+	chr3	185655611	+	.	27	72	1836245_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=1836245_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_185636501_185661501_192C;SPAN=5970;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:88 DP:217 GQ:99 PL:[231.8, 0.0, 294.5] SR:72 DR:27 LR:-231.7 LO:232.1);ALT=C[chr3:185655611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186288754	+	chr3	186289883	+	.	0	16	1838487_1	20.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1838487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_186273501_186298501_282C;SPAN=1129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:121 GQ:20.3 PL:[20.3, 0.0, 271.1] SR:16 DR:0 LR:-20.03 LO:33.1);ALT=G[chr3:186289883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7694765	+	chr3	186314753	+	.	19	0	1838693_1	37.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=1838693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186314753(-)-19:7694765(+)__3_186298001_186323001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:93 GQ:37.7 PL:[37.7, 0.0, 186.2] SR:0 DR:19 LR:-37.52 LO:43.26);ALT=]chr19:7694765]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	186442176	+	chr3	186513632	+	.	8	13	1839246_1	39.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1839246_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_186494001_186519001_222C;SPAN=71456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:50 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:13 DR:8 LR:-39.27 LO:40.1);ALT=T[chr3:186513632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186469052	-	chr8	64032515	+	.	21	8	1839231_1	80.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=TTGTATTTTTAGTAGAGACGGGGTTTCACCGTGTTAGCCAGGATGGTCTTGATCTCCTGA;MAPQ=60;MATEID=1839231_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_3_186445001_186470001_9C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:57 GQ:57.2 PL:[80.3, 0.0, 57.2] SR:8 DR:21 LR:-80.48 LO:80.48);ALT=[chr8:64032515[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	186501450	+	chrX	52862812	-	.	41	0	7424856_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7424856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186501450(+)-23:52862812(+)__23_52846501_52871501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:28 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=G]chrX:52862812];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	186501451	+	chr3	186503669	+	.	18	0	1839284_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1839284_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186501451(+)-3:186503669(-)__3_186494001_186519001D;SPAN=2218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:102 GQ:32 PL:[32.0, 0.0, 213.5] SR:0 DR:18 LR:-31.78 LO:39.7);ALT=C[chr3:186503669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186501451	+	chr3	186502747	+	.	10	0	1839283_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1839283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186501451(+)-3:186502747(-)__3_186494001_186519001D;SPAN=1296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=C[chr3:186502747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186502485	+	chr3	186503670	+	.	7	45	1839288_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1839288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_186494001_186519001_368C;SPAN=1185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:114 GQ:99 PL:[131.0, 0.0, 144.2] SR:45 DR:7 LR:-130.9 LO:130.9);ALT=G[chr3:186503670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186581033	+	chr3	186585285	+	.	75	42	1839808_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GAAAAATATTGCAAATAG;MAPQ=60;MATEID=1839808_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_186567501_186592501_262C;SPAN=4252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:85 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:42 DR:75 LR:-293.8 LO:293.8);ALT=G[chr3:186585285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	186585325	+	chr19	45118991	-	.	23	0	1839837_1	65.0	.	DISC_MAPQ=8;EVDNC=DSCRD;IMPRECISE;MAPQ=8;MATEID=1839837_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:186585325(+)-19:45118991(+)__3_186567501_186592501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:0 DR:23 LR:-65.7 LO:65.7);ALT=G]chr19:45118991];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	187085160	-	chr22	30993411	+	.	22	21	1841562_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=CACCAATCAGCACCCTGTGTCTAGCTCA;MAPQ=22;MATEID=1841562_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_187082001_187107001_168C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:63 GQ:39.2 PL:[111.8, 0.0, 39.2] SR:21 DR:22 LR:-113.4 LO:113.4);ALT=[chr22:30993411[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	187872080	+	chr3	187925985	+	.	13	0	1844323_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=1844323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:187872080(+)-3:187925985(-)__3_187915001_187940001D;SPAN=53905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:50 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:0 DR:13 LR:-29.37 LO:31.17);ALT=G[chr3:187925985[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	192875332	+	chr3	192885406	+	.	46	38	1860239_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TCT;MAPQ=60;MATEID=1860239_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_192864001_192889001_30C;SPAN=10074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:70 GQ:15.6 PL:[201.3, 15.6, 0.0] SR:38 DR:46 LR:-202.4 LO:202.4);ALT=T[chr3:192885406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	92116020	+	chr3	193258757	+	.	18	79	5843956_1	99.0	.	DISC_MAPQ=4;EVDNC=ASDIS;MAPQ=43;MATEID=5843956_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_92095501_92120501_270C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:36 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:79 DR:18 LR:-274.0 LO:274.0);ALT=]chr14:92116020]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr3	193311198	+	chr3	193332511	+	.	9	7	1861844_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1861844_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_193329501_193354501_223C;SPAN=21313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:78 GQ:21.8 PL:[21.8, 0.0, 167.0] SR:7 DR:9 LR:-21.78 LO:28.31);ALT=G[chr3:193332511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	193430615	+	chr15	71379741	-	.	5	19	1862286_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGCAA;MAPQ=60;MATEID=1862286_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_193427501_193452501_81C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:28 GQ:12.2 PL:[55.1, 0.0, 12.2] SR:19 DR:5 LR:-56.61 LO:56.61);ALT=T]chr15:71379741];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	193829745	+	chr9	130506502	-	.	10	0	1863681_1	23.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=1863681_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:193829745(+)-9:130506502(+)__3_193819501_193844501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:36 GQ:23.3 PL:[23.3, 0.0, 62.9] SR:0 DR:10 LR:-23.26 LO:24.32);ALT=T]chr9:130506502];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	194458297	+	chr3	194456950	+	.	27	0	1865933_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1865933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:194456950(-)-3:194458297(+)__3_194432001_194457001D;SPAN=1347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:42 GQ:21.8 PL:[77.9, 0.0, 21.8] SR:0 DR:27 LR:-79.3 LO:79.3);ALT=]chr3:194458297]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	194543294	+	chr3	194546257	+	.	0	78	1866317_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GGTG;MAPQ=60;MATEID=1866317_2;MATENM=0;NM=5;NUMPARTS=3;SCTG=c_3_194530001_194555001_108C;SPAN=2963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:88 GQ:20.4 PL:[254.1, 20.4, 0.0] SR:78 DR:0 LR:-254.8 LO:254.8);ALT=G[chr3:194546257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	194546431	+	chr3	194543310	+	.	78	92	1866318_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1866318_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_194530001_194555001_83C;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:99 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:92 DR:78 LR:-429.1 LO:429.1);ALT=]chr3:194546431]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	195053852	+	chr3	195063200	+	TGATTTTAGGATTTCTGATCTCCTTTTTGATTGAAGAACATTAAT	4	8	1867914_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTGA;INSERTION=TGATTTTAGGATTTCTGATCTCCTTTTTGATTGAAGAACATTAAT;MAPQ=60;MATEID=1867914_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_195044501_195069501_95C;SPAN=9348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:8 DR:4 LR:-5.326 LO:17.45);ALT=T[chr3:195063200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	195102800	+	chr3	195163589	+	.	22	0	1868410_1	56.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1868410_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195102800(+)-3:195163589(-)__3_195142501_195167501D;SPAN=60789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:59 GQ:56.6 PL:[56.6, 0.0, 86.3] SR:0 DR:22 LR:-56.64 LO:56.98);ALT=T[chr3:195163589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	195112925	+	chr3	195163657	+	.	21	0	1868412_1	55.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1868412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195112925(+)-3:195163657(-)__3_195142501_195167501D;SPAN=50732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:50 GQ:55.7 PL:[55.7, 0.0, 65.6] SR:0 DR:21 LR:-55.78 LO:55.82);ALT=A[chr3:195163657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	195400669	+	chr5	236627	+	.	11	0	1869848_1	11.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=1869848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195400669(+)-5:236627(-)__3_195387501_195412501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:93 GQ:11.3 PL:[11.3, 0.0, 212.6] SR:0 DR:11 LR:-11.12 LO:22.18);ALT=T[chr5:236627[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr3	195412855	-	chr5	1572306	+	.	10	0	1871043_1	8.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=1871043_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195412855(-)-5:1572306(-)__3_195412001_195437001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:0 DR:10 LR:-7.814 LO:19.72);ALT=[chr5:1572306[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	195671187	+	chr3	195668842	+	.	11	0	1871543_1	0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=1871543_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195668842(-)-3:195671187(+)__3_195657001_195682001D;SPAN=2345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:156 GQ:5.8 PL:[0.0, 5.8, 389.4] SR:0 DR:11 LR:5.953 LO:19.59);ALT=]chr3:195671187]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr3	195971910	+	chr3	196346529	-	.	8	0	1875013_1	16.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=1875013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:195971910(+)-3:196346529(+)__3_196343001_196368001D;SPAN=374619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:37 GQ:16.4 PL:[16.4, 0.0, 72.5] SR:0 DR:8 LR:-16.38 LO:18.44);ALT=A]chr3:196346529];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr3	196018245	+	chr3	196022876	+	.	0	7	1873452_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1873452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196000001_196025001_221C;SPAN=4631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:111 GQ:6.6 PL:[0.0, 6.6, 280.5] SR:7 DR:0 LR:6.966 LO:12.11);ALT=C[chr3:196022876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196043104	+	chr3	196044910	+	.	0	8	1873537_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=1873537_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196024501_196049501_209C;SPAN=1806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:8 DR:0 LR:5.29 LO:14.13);ALT=T[chr3:196044910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196366747	+	chr3	196381398	+	.	45	13	1875112_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1875112_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_3_196343001_196368001_446C;SPAN=14651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:48 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:13 DR:45 LR:-145.2 LO:145.2);ALT=G[chr3:196381398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196467029	+	chr3	196509496	+	.	50	58	1875735_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1875735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196465501_196490501_162C;SPAN=42467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:70 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:58 DR:50 LR:-250.9 LO:250.9);ALT=G[chr3:196509496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196664519	+	chr3	196666122	+	.	0	9	1876313_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1876313_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196661501_196686501_13C;SPAN=1603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:9 DR:0 LR:-1.262 LO:16.82);ALT=T[chr3:196666122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196666304	+	chr3	196669296	+	.	25	4	1876323_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1876323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196661501_196686501_169C;SPAN=2992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:101 GQ:65.3 PL:[65.3, 0.0, 177.5] SR:4 DR:25 LR:-65.07 LO:68.06);ALT=C[chr3:196669296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196678923	+	chr3	196695614	+	.	9	0	1876501_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1876501_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:196678923(+)-3:196695614(-)__3_196686001_196711001D;SPAN=16691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:20 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.29 LO:24.29);ALT=T[chr3:196695614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	196934573	+	chr3	196939256	+	CAGACT	56	38	1877108_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CAGACT;MAPQ=60;MATEID=1877108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_196931001_196956001_77C;SPAN=4683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:70 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:38 DR:56 LR:-217.9 LO:217.9);ALT=A[chr3:196939256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197273358	+	chr3	197282652	+	.	0	12	1878613_1	25.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1878613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_197249501_197274501_402C;SPAN=9294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:54 GQ:25.1 PL:[25.1, 0.0, 104.3] SR:12 DR:0 LR:-24.98 LO:27.82);ALT=C[chr3:197282652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197476945	+	chr3	197483296	+	.	13	9	1879051_1	33.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1879051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_197470001_197495001_51C;SPAN=6351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:96 GQ:33.5 PL:[33.5, 0.0, 198.5] SR:9 DR:13 LR:-33.41 LO:40.23);ALT=G[chr3:197483296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197483430	+	chr3	197495309	+	.	0	7	1879077_1	7.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=1879077_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_197470001_197495001_290C;SPAN=11879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:57 GQ:7.7 PL:[7.7, 0.0, 129.8] SR:7 DR:0 LR:-7.664 LO:14.24);ALT=T[chr3:197495309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197677850	+	chr3	197680874	+	CTGTGGTCCAAGGCCATTTTTGCTGGCTATAAGCGGGGTCTCCGGAACCAAAGGGAGCACACAGCTCTTCTTAAAATTGAAGGTGTTTACGCCCGAGATGAAACAGAATTCTATTTGGGCAAGAGATGCGCTTATGTATATAAAGCAAAGAA	2	161	1880776_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTGTGGTCCAAGGCCATTTTTGCTGGCTATAAGCGGGGTCTCCGGAACCAAAGGGAGCACACAGCTCTTCTTAAAATTGAAGGTGTTTACGCCCGAGATGAAACAGAATTCTATTTGGGCAAGAGATGCGCTTATGTATATAAAGCAAAGAA;MAPQ=60;MATEID=1880776_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_3_197666001_197691001_29C;SPAN=3024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:163 DP:454 GQ:99 PL:[415.3, 0.0, 685.9] SR:161 DR:2 LR:-415.1 LO:418.7);ALT=G[chr3:197680874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197681000	+	chr3	197682619	+	.	20	0	1880790_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1880790_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:197681000(+)-3:197682619(-)__3_197666001_197691001D;SPAN=1619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:20 DP:524 GQ:75.6 PL:[0.0, 75.6, 1423.0] SR:0 DR:20 LR:75.95 LO:30.16);ALT=T[chr3:197682619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	197843929	+	chr3	197850167	+	.	92	79	1881562_1	99.0	.	DISC_MAPQ=25;EVDNC=ASDIS;HOMSEQ=GGC;MAPQ=60;MATEID=1881562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_197837501_197862501_505C;SPAN=6238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:36 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:79 DR:92 LR:-425.8 LO:425.8);ALT=C[chr3:197850167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	86017	+	chr4	367143	+	.	10	23	1882552_1	91.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGGAGAGAAACCCTACAAATGTGAAAAATGTGGCAAAGC;MAPQ=60;MATEID=1882552_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_4_343001_368001_242C;SPAN=281126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:42 GQ:8.6 PL:[91.1, 0.0, 8.6] SR:23 DR:10 LR:-94.59 LO:94.59);ALT=C[chr4:367143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	666358	+	chr4	667998	+	.	48	0	1883237_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=1883237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:666358(+)-4:667998(-)__4_661501_686501D;SPAN=1640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:164 GQ:99 PL:[114.2, 0.0, 282.5] SR:0 DR:48 LR:-114.0 LO:118.0);ALT=T[chr4:667998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	926358	+	chr4	941523	+	.	13	0	1883857_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1883857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:926358(+)-4:941523(-)__4_906501_931501D;SPAN=15165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:19 GQ:8 PL:[37.7, 0.0, 8.0] SR:0 DR:13 LR:-38.82 LO:38.82);ALT=T[chr4:941523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1193884	+	chr4	1195116	+	.	9	0	1884657_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1884657_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1193884(+)-4:1195116(-)__4_1176001_1201001D;SPAN=1232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=G[chr4:1195116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1219356	+	chr4	1221986	+	.	3	2	1884743_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=1884743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1200501_1225501_218C;SPAN=2630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:47 GQ:0.5 PL:[0.5, 0.0, 112.7] SR:2 DR:3 LR:-0.4706 LO:7.462);ALT=T[chr4:1221986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1222133	+	chr4	1231969	+	.	0	7	1884748_1	16.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=1884748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1200501_1225501_34C;SPAN=9836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:26 GQ:16.1 PL:[16.1, 0.0, 45.8] SR:7 DR:0 LR:-16.06 LO:16.91);ALT=T[chr4:1231969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1267490	+	chr4	1266053	+	.	37	0	1885387_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=1885387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1266053(-)-4:1267490(+)__4_1249501_1274501D;SPAN=1437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:71 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.2 LO:103.2);ALT=]chr4:1267490]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	1283777	+	chr4	1305781	+	.	9	0	1885287_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1885287_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:1283777(+)-4:1305781(-)__4_1298501_1323501D;SPAN=22004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=G[chr4:1305781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1576273	+	chr4	1581885	+	.	2	3	1885614_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1885614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1568001_1593001_100C;SPAN=5612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:44 GQ:4.7 PL:[4.7, 0.0, 100.4] SR:3 DR:2 LR:-4.584 LO:9.99);ALT=T[chr4:1581885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1705429	+	chr4	1713601	+	.	0	20	1886112_1	50.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=1886112_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_1690501_1715501_260C;SPAN=8172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:59 GQ:50 PL:[50.0, 0.0, 92.9] SR:20 DR:0 LR:-50.04 LO:50.75);ALT=T[chr4:1713601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1725597	+	chr4	1729435	+	.	15	12	1886005_1	49.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1886005_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1715001_1740001_260C;SPAN=3838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:51 GQ:49.1 PL:[49.1, 0.0, 72.2] SR:12 DR:15 LR:-48.9 LO:49.2);ALT=A[chr4:1729435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1873269	+	chr4	1902351	+	.	7	4	1886367_1	23.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=1886367_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_1886501_1911501_142C;SPAN=29082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:4 DR:7 LR:-23.21 LO:23.34);ALT=G[chr4:1902351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	1993444	+	chr4	2010477	+	.	0	7	1886489_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1886489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2009001_2034001_195C;SPAN=17033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:40 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:7 DR:0 LR:-12.27 LO:15.41);ALT=T[chr4:2010477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2044551	+	chr4	2045587	+	.	0	59	1886589_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=1886589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2033501_2058501_225C;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:84 GQ:30.2 PL:[172.1, 0.0, 30.2] SR:59 DR:0 LR:-177.5 LO:177.5);ALT=G[chr4:2045587[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2845752	+	chr4	2877621	+	.	20	7	1888270_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=1888270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2842001_2867001_53C;SPAN=31869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:21 DP:8 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:7 DR:20 LR:-59.41 LO:59.41);ALT=G[chr4:2877621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2877838	+	chr4	2883625	+	.	2	5	1888231_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1888231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2866501_2891501_93C;SPAN=5787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:55 GQ:8.3 PL:[8.3, 0.0, 123.8] SR:5 DR:2 LR:-8.206 LO:14.35);ALT=G[chr4:2883625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2883789	+	chr4	2886242	+	.	2	3	1888240_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=1888240_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2866501_2891501_31C;SPAN=2453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:55 GQ:1.5 PL:[0.0, 1.5, 135.3] SR:3 DR:2 LR:1.697 LO:7.178);ALT=T[chr4:2886242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2901163	+	chr4	2906490	+	.	4	4	1888342_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=1888342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2891001_2916001_175C;SPAN=5327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:62 GQ:3.2 PL:[3.2, 0.0, 145.1] SR:4 DR:4 LR:-3.009 LO:11.54);ALT=G[chr4:2906490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	2959469	+	chr4	2964852	+	.	7	10	1888496_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1888496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_2940001_2965001_36C;SPAN=5383;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:10 DR:7 LR:-23.36 LO:27.2);ALT=T[chr4:2964852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	3364879	+	chr4	3363369	+	.	21	0	1889234_1	52.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1889234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3363369(-)-4:3364879(+)__4_3356501_3381501D;SPAN=1510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:64 GQ:52.1 PL:[52.1, 0.0, 101.6] SR:0 DR:21 LR:-51.98 LO:52.91);ALT=]chr4:3364879]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	3514786	+	chr4	3516475	+	.	9	0	1889532_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1889532_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3514786(+)-4:3516475(-)__4_3503501_3528501D;SPAN=1689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=A[chr4:3516475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	3517926	+	chr4	3519761	+	.	2	4	1889536_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=1889536_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_3503501_3528501_259C;SPAN=1835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:48 GQ:6.8 PL:[6.8, 0.0, 109.1] SR:4 DR:2 LR:-6.802 LO:12.25);ALT=C[chr4:3519761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	3520720	+	chr4	3521798	+	.	5	4	1889547_1	10.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=1889547_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_3503501_3528501_63C;SPAN=1078;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:4 DR:5 LR:-10.37 LO:14.87);ALT=T[chr4:3521798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	3526778	+	chr4	3533936	+	.	0	109	1890164_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=1890164_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_3528001_3553001_297C;SPAN=7158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:52 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:109 DR:0 LR:-323.5 LO:323.5);ALT=G[chr4:3533936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	3570224	+	chr4	3568952	+	.	22	0	1890338_1	42.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=1890338_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3568952(-)-4:3570224(+)__4_3552501_3577501D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:111 GQ:42.8 PL:[42.8, 0.0, 224.3] SR:0 DR:22 LR:-42.55 LO:49.76);ALT=]chr4:3570224]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	3575944	+	chr19	51378983	+	.	9	0	1890408_1	5.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=1890408_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3575944(+)-19:51378983(-)__4_3552501_3577501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:0 DR:9 LR:-5.597 LO:17.5);ALT=G[chr19:51378983[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr19	51379108	+	chr4	3576050	+	.	12	0	1890412_1	27.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=1890412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3576050(-)-19:51379108(+)__4_3552501_3577501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:44 GQ:27.8 PL:[27.8, 0.0, 77.3] SR:0 DR:12 LR:-27.69 LO:29.07);ALT=]chr19:51379108]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	4175792	+	chr4	3903140	+	.	15	0	1891016_1	44.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=1891016_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3903140(-)-4:4175792(+)__4_4165001_4190001D;SPAN=272652;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:19 GQ:1.4 PL:[44.3, 0.0, 1.4] SR:0 DR:15 LR:-46.75 LO:46.75);ALT=]chr4:4175792]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	3903331	+	chr4	4176050	+	.	16	0	1891017_1	52.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=1891017_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:3903331(+)-4:4176050(-)__4_4165001_4190001D;SPAN=272719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:18 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:16 LR:-52.35 LO:52.35);ALT=T[chr4:4176050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	4276496	+	chr4	4281173	+	.	0	7	1891389_1	9.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1891389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_4263001_4288001_235C;SPAN=4677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=C[chr4:4281173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	4285557	+	chr4	4291787	+	.	10	0	1891421_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1891421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:4285557(+)-4:4291787(-)__4_4287501_4312501D;SPAN=6230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:0 DR:10 LR:-26.78 LO:26.78);ALT=A[chr4:4291787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	4543524	-	chr17	28395777	+	.	8	4	6359037_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACTTCGCGGGCCCGGCTGGAGAAGTCGCCCTTGGGCC;MAPQ=60;MATEID=6359037_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_17_28395501_28420501_270C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:4 DR:8 LR:-24.12 LO:26.03);ALT=[chr17:28395777[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	5018691	+	chr4	5021019	+	GTGTATGTCCAGGTACAGCCTGGGCAGGTATCTCACACATGGCT	0	27	1892764_1	73.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GTGTATGTCCAGGTACAGCCTGGGCAGGTATCTCACACATGGCT;MAPQ=60;MATEID=1892764_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_4998001_5023001_164C;SPAN=2328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:58 GQ:66.8 PL:[73.4, 0.0, 66.8] SR:27 DR:0 LR:-73.43 LO:73.43);ALT=T[chr4:5021019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	5018961	+	chr4	5021096	+	.	23	0	1892766_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1892766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:5018961(+)-4:5021096(-)__4_4998001_5023001D;SPAN=2135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:62 GQ:59.3 PL:[59.3, 0.0, 89.0] SR:0 DR:23 LR:-59.13 LO:59.5);ALT=A[chr4:5021096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	6173251	+	chr17	54870116	-	.	8	0	6441813_1	20.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6441813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:6173251(+)-17:54870116(+)__17_54855501_54880501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:0 DR:8 LR:-19.91 LO:20.23);ALT=T]chr17:54870116];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	6651593	+	chr4	6652911	+	.	63	47	1895414_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CAGA;MAPQ=60;MATEID=1895414_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_6639501_6664501_271C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:24 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:47 DR:63 LR:-270.7 LO:270.7);ALT=A[chr4:6652911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	6784578	+	chr4	6825909	+	.	8	0	1895563_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1895563_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:6784578(+)-4:6825909(-)__4_6762001_6787001D;SPAN=41331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:8 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=G[chr4:6825909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	6897382	+	chr4	6900394	+	.	16	0	1895913_1	41.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=1895913_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:6897382(+)-4:6900394(-)__4_6884501_6909501D;SPAN=3012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:41 GQ:41.9 PL:[41.9, 0.0, 55.1] SR:0 DR:16 LR:-41.71 LO:41.85);ALT=T[chr4:6900394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	6911678	+	chr4	6925099	+	.	19	7	1895846_1	57.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=1895846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_6909001_6934001_149C;SPAN=13421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:43 GQ:44.6 PL:[57.8, 0.0, 44.6] SR:7 DR:19 LR:-57.73 LO:57.73);ALT=G[chr4:6925099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	7064194	+	chr4	7065787	+	.	0	7	1896138_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=1896138_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_7056001_7081001_172C;SPAN=1593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:41 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:7 DR:0 LR:-12.0 LO:15.33);ALT=C[chr4:7065787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	7065962	+	chr4	7069708	+	.	12	0	1896142_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1896142_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:7065962(+)-4:7069708(-)__4_7056001_7081001D;SPAN=3746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:51 GQ:26 PL:[26.0, 0.0, 95.3] SR:0 DR:12 LR:-25.8 LO:28.16);ALT=T[chr4:7069708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	7995809	+	chr4	7996894	+	.	63	32	1898035_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGGAAGCATTCTT;MAPQ=60;MATEID=1898035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_7987001_8012001_254C;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:104 GQ:8.3 PL:[242.6, 0.0, 8.3] SR:32 DR:63 LR:-255.4 LO:255.4);ALT=T[chr4:7996894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	8168999	+	chr4	8167984	+	.	19	0	1898236_1	42.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1898236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:8167984(-)-4:8168999(+)__4_8158501_8183501D;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:74 GQ:42.8 PL:[42.8, 0.0, 135.2] SR:0 DR:19 LR:-42.67 LO:45.43);ALT=]chr4:8168999]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	9457101	+	chr4	9481577	+	.	15	0	1901104_1	49.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=1901104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:9457101(+)-4:9481577(-)__4_9481501_9506501D;SPAN=24476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:17 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:15 LR:-48.87 LO:48.87);ALT=A[chr4:9481577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	9583341	+	chr12	8495209	-	.	8	0	5087171_1	14.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=5087171_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:9583341(+)-12:8495209(+)__12_8477001_8502001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=G]chr12:8495209];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	10077110	+	chr4	10078928	+	.	9	6	1902575_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1902575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_10069501_10094501_223C;SPAN=1818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:62 GQ:29.6 PL:[29.6, 0.0, 118.7] SR:6 DR:9 LR:-29.42 LO:32.57);ALT=T[chr4:10078928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	10100765	+	chr4	10118275	+	CCGGAGGCAATGTAGAATCCGCTGGGCGCATACTTGGCCACCACCACCTGATGGGCGTGCTCTGTGTAGATGTCAGCAAGGGCTGGGTTGTCGATGTTCCTTAGGATGACGCACTTTCCATTGGTGTACAGAAAATTGTTGCCCTTAGGGTCGCCGCCGATGATCTTGGAGACGCCCCTCTCCACCTGCGGGAGGCTGGCGAACACCTTCT	7	39	1902624_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCGGAGGCAATGTAGAATCCGCTGGGCGCATACTTGGCCACCACCACCTGATGGGCGTGCTCTGTGTAGATGTCAGCAAGGGCTGGGTTGTCGATGTTCCTTAGGATGACGCACTTTCCATTGGTGTACAGAAAATTGTTGCCCTTAGGGTCGCCGCCGATGATCTTGGAGACGCCCCTCTCCACCTGCGGGAGGCTGGCGAACACCTTCT;MAPQ=60;MATEID=1902624_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_4_10094001_10119001_182C;SPAN=17510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:34 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:39 DR:7 LR:-118.8 LO:118.8);ALT=T[chr4:10118275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	10105658	+	chr4	10118307	+	.	32	0	1902634_1	94.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=1902634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:10105658(+)-4:10118307(-)__4_10094001_10119001D;SPAN=12649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:42 GQ:5.3 PL:[94.4, 0.0, 5.3] SR:0 DR:32 LR:-98.59 LO:98.59);ALT=A[chr4:10118307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	10211267	+	chr4	10234568	+	.	65	49	1902852_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTTTCAA;MAPQ=60;MATEID=1902852_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_10192001_10217001_168C;SPAN=23301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:12 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:49 DR:65 LR:-267.4 LO:267.4);ALT=A[chr4:10234568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	17510987	+	chr4	17513573	+	.	0	7	1913226_1	4.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1913226_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_17493001_17518001_43C;SPAN=2586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:71 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:7 DR:0 LR:-3.871 LO:13.53);ALT=C[chr4:17513573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	17579208	+	chr6	36641580	+	.	43	0	1913378_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1913378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:17579208(+)-6:36641580(-)__4_17566501_17591501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:23 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=G[chr6:36641580[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	17616352	+	chr4	17623207	+	.	17	0	1913628_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1913628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:17616352(+)-4:17623207(-)__4_17615501_17640501D;SPAN=6855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:53 GQ:41.9 PL:[41.9, 0.0, 84.8] SR:0 DR:17 LR:-41.76 LO:42.63);ALT=C[chr4:17623207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	17616352	+	chr4	17621520	+	.	22	0	1913627_1	56.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1913627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:17616352(+)-4:17621520(-)__4_17615501_17640501D;SPAN=5168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:58 GQ:56.9 PL:[56.9, 0.0, 83.3] SR:0 DR:22 LR:-56.91 LO:57.19);ALT=C[chr4:17621520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	18371282	+	chr19	16096606	-	.	8	0	6747306_1	23.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6747306_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:18371282(+)-19:16096606(+)__19_16096501_16121501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:4 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=A]chr19:16096606];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	18419959	-	chr12	131712701	+	.	22	0	5397686_1	62.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=5397686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:18419959(-)-12:131712701(-)__12_131712001_131737001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:21 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:0 DR:22 LR:-62.72 LO:62.72);ALT=[chr12:131712701[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	18420151	+	chr12	131712545	-	.	33	0	5397687_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5397687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:18420151(+)-12:131712545(+)__12_131712001_131737001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:33 LR:-102.3 LO:102.3);ALT=G]chr12:131712545];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	19079465	+	chr4	19085551	+	.	17	12	1915948_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCACTGATTTGCTTT;MAPQ=60;MATEID=1915948_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_19061001_19086001_96C;SPAN=6086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:22 DP:2727 GQ:99 PL:[0.0, 665.5, 7955.0] SR:12 DR:17 LR:666.2 LO:18.58);ALT=T[chr4:19085551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39030219	+	chr4	39033846	+	.	15	16	1944220_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1944220_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_39028501_39053501_157C;SPAN=3627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:52 GQ:62 PL:[62.0, 0.0, 62.0] SR:16 DR:15 LR:-61.84 LO:61.84);ALT=T[chr4:39033846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39344090	+	chr4	39352966	+	AATCATAGATGATCCTCTTTTTCTTGCTTGGTTGCTTTTGTTTGAAGTCATCCTCTTTACGGGAGCTATTT	2	22	1944689_1	66.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=AATCATAGATGATCCTCTTTTTCTTGCTTGGTTGCTTTTGTTTGAAGTCATCCTCTTTACGGGAGCTATTT;MAPQ=60;MATEID=1944689_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_39347001_39372001_45C;SPAN=8876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:22 GQ:6 PL:[66.0, 6.0, 0.0] SR:22 DR:2 LR:-66.02 LO:66.02);ALT=G[chr4:39352966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39344090	+	chr4	39347021	+	.	3	11	1944688_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=1944688_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_39347001_39372001_45C;SPAN=2931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:24 GQ:20 PL:[36.5, 0.0, 20.0] SR:11 DR:3 LR:-36.61 LO:36.61);ALT=G[chr4:39347021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39347127	+	chr4	39367892	+	.	8	0	1944692_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=1944692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:39347127(+)-4:39367892(-)__4_39347001_39372001D;SPAN=20765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=A[chr4:39367892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39353097	+	chr4	39367858	+	.	16	6	1944701_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1944701_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_39347001_39372001_234C;SPAN=14761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:56 GQ:47.6 PL:[47.6, 0.0, 87.2] SR:6 DR:16 LR:-47.55 LO:48.22);ALT=C[chr4:39367858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39460784	+	chr4	39462409	+	.	6	2	1945038_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=1945038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_39445001_39470001_187C;SPAN=1625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:65 GQ:5.6 PL:[5.6, 0.0, 150.8] SR:2 DR:6 LR:-5.497 LO:13.81);ALT=T[chr4:39462409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39606801	+	chr4	39640359	+	.	13	8	1945344_1	40.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=1945344_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_39616501_39641501_92C;SPAN=33558;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:34 GQ:40.4 PL:[40.4, 0.0, 40.4] SR:8 DR:13 LR:-40.3 LO:40.31);ALT=C[chr4:39640359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39700010	+	chr4	39739038	+	.	0	12	1945891_1	31.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1945891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_39739001_39764001_83C;SPAN=39028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:30 GQ:31.4 PL:[31.4, 0.0, 41.3] SR:12 DR:0 LR:-31.48 LO:31.56);ALT=G[chr4:39739038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39814526	+	chr4	39815872	+	CTGGGTGTGTGGTTGTGATTGGGTGTGTGGTGTGGGTGTCTGAGTGTGGGTGTGTGGTTGTGATTGTGAGTGTGGGCGTGA	6	118	1946150_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;INSERTION=CTGGGTGTGTGGTTGTGATTGGGTGTGTGGTGTGGGTGTCTGAGTGTGGGTGTGTGGTTGTGATTGTGAGTGTGGGCGTGA;MAPQ=53;MATEID=1946150_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_39812501_39837501_122C;SPAN=1346;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:119 DP:219 GQ:99 PL:[333.5, 0.0, 198.2] SR:118 DR:6 LR:-335.3 LO:335.3);ALT=T[chr4:39815872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	39968868	-	chr4	39970061	+	.	9	0	1946316_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1946316_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:39968868(-)-4:39970061(-)__4_39959501_39984501D;SPAN=1193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:0 DR:9 LR:-14.0 LO:19.3);ALT=[chr4:39970061[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	101717277	+	chr4	39974899	+	.	8	0	3995857_1	13.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=3995857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:39974899(-)-8:101717277(+)__8_101699501_101724501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=]chr8:101717277]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	40011028	-	chr18	23771459	+	.	2	5	1946665_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=1946665_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_40008501_40033501_198C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:25 GQ:9.8 PL:[9.8, 0.0, 49.4] SR:5 DR:2 LR:-9.732 LO:11.33);ALT=[chr18:23771459[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	40024955	+	chr4	40026282	+	.	20	15	1946691_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GGCCGGGTGTGGTGGCTCACGCCTGTAATCCCAGCACTTT;MAPQ=60;MATEID=1946691_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_4_40008501_40033501_150C;SPAN=1327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:15 DR:20 LR:-99.02 LO:99.02);ALT=T[chr4:40026282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	40198920	+	chr4	40244331	+	.	0	10	1946971_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=1946971_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_40229001_40254001_301C;SPAN=45411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:26 GQ:26 PL:[26.0, 0.0, 35.9] SR:10 DR:0 LR:-25.97 LO:26.07);ALT=G[chr4:40244331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	40235027	-	chr4	40237059	+	.	28	17	1946983_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=1946983_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_4_40229001_40254001_68C;SPAN=2032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:41 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:17 DR:28 LR:-118.8 LO:118.8);ALT=[chr4:40237059[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	54319300	+	chr4	54325467	+	CGATGAAGAACGATACAGATACAGGGAATATGCAGAAAGAGGTTATGAGCGTCACAGAGCAAGTCGAGAAAAAGAAGAACGACATAGAGAAAGACGACACAGGGAGAAAGAGGAAACCAGACATAAGTCTTCTCGA	2	14	1969332_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CGATGAAGAACGATACAGATACAGGGAATATGCAGAAAGAGGTTATGAGCGTCACAGAGCAAGTCGAGAAAAAGAAGAACGACATAGAGAAAGACGACACAGGGAGAAAGAGGAAACCAGACATAAGTCTTCTCGA;MAPQ=60;MATEID=1969332_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_54316501_54341501_135C;SPAN=6167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:89 GQ:25.4 PL:[25.4, 0.0, 190.4] SR:14 DR:2 LR:-25.4 LO:32.75);ALT=G[chr4:54325467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	54319300	+	chr4	54324817	+	.	3	8	1969331_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=1969331_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_54316501_54341501_135C;SPAN=5517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:91 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:8 DR:3 LR:-8.356 LO:19.82);ALT=G[chr4:54324817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	64563186	+	chr9	135361784	-	.	2	19	2001515_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACACA;MAPQ=60;MATEID=2001515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_64557501_64582501_161C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:45 GQ:50.6 PL:[50.6, 0.0, 57.2] SR:19 DR:2 LR:-50.53 LO:50.56);ALT=G]chr9:135361784];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	67928939	+	chr4	66372379	+	.	16	0	2011642_1	39.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=2011642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:66372379(-)-4:67928939(+)__4_67914001_67939001D;SPAN=1556560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.0 LO:39.93);ALT=]chr4:67928939]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	68411083	-	chr12	89893844	+	.	17	0	5281783_1	44.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5281783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:68411083(-)-12:89893844(-)__12_89890501_89915501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:42 GQ:44.9 PL:[44.9, 0.0, 54.8] SR:0 DR:17 LR:-44.74 LO:44.82);ALT=[chr12:89893844[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	68547934	+	chr4	68562363	+	.	0	7	2013567_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CTA;MAPQ=60;MATEID=2013567_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_68551001_68576001_170C;SPAN=14429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:43 GQ:11.6 PL:[11.6, 0.0, 90.8] SR:7 DR:0 LR:-11.46 LO:15.17);ALT=A[chr4:68562363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	68547954	+	chr4	68566791	+	.	9	0	2013568_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2013568_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:68547954(+)-4:68566791(-)__4_68551001_68576001D;SPAN=18837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:0 DR:9 LR:-15.35 LO:19.68);ALT=A[chr4:68566791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	68855990	-	chr6	45256305	+	CACACAC	3	19	2014505_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TATATATATATATATA;INSERTION=CACACAC;MAPQ=60;MATEID=2014505_2;MATENM=0;NM=7;NUMPARTS=3;REPSEQ=TATATATATATA;SCTG=c_4_68845001_68870001_33C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:32 GQ:1.7 PL:[21.0, 0.0, 1.7] SR:19 DR:3 LR:-21.82 LO:21.82);ALT=[chr6:45256305[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	68957530	-	chr8	141428790	+	.	8	0	2015303_1	16.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2015303_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:68957530(-)-8:141428790(-)__4_68943001_68968001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:0 DR:8 LR:-16.11 LO:18.33);ALT=[chr8:141428790[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	69180041	+	chr4	69182032	+	.	4	4	2015515_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2015515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_69163501_69188501_38C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:97 GQ:3 PL:[0.0, 3.0, 240.9] SR:4 DR:4 LR:3.173 LO:12.54);ALT=G[chr4:69182032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	69204104	+	chr4	69215444	+	.	0	11	2015613_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2015613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_69212501_69237501_3C;SPAN=11340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:58 GQ:20.6 PL:[20.6, 0.0, 119.6] SR:11 DR:0 LR:-20.6 LO:24.64);ALT=T[chr4:69215444[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56642594	+	chr4	69242035	+	.	29	0	6219218_1	85.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6219218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:69242035(-)-16:56642594(+)__16_56619501_56644501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:25 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=]chr16:56642594]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	69373781	+	chr4	69491144	+	.	10	0	2016300_1	23.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2016300_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:69373781(+)-4:69491144(-)__4_69482001_69507001D;SPAN=117363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:36 GQ:23.3 PL:[23.3, 0.0, 62.9] SR:0 DR:10 LR:-23.26 LO:24.32);ALT=A[chr4:69491144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	69505212	+	chr4	69506268	-	.	9	0	2016350_1	4.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=2016350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:69505212(+)-4:69506268(+)__4_69482001_69507001D;SPAN=1056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:0 DR:9 LR:-4.242 LO:17.27);ALT=T]chr4:69506268];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	70052508	+	chr4	70167672	-	.	11	0	2018080_1	23.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2018080_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70052508(+)-4:70167672(+)__4_70143501_70168501D;SPAN=115164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:47 GQ:23.6 PL:[23.6, 0.0, 89.6] SR:0 DR:11 LR:-23.58 LO:25.79);ALT=G]chr4:70167672];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	70053058	-	chr4	70167189	+	.	28	0	2017974_1	85.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=2017974_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70053058(-)-4:70167189(-)__4_70045501_70070501D;SPAN=114131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:29 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:28 LR:-85.82 LO:85.82);ALT=[chr4:70167189[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	70107417	-	chr4	70173859	+	.	9	0	2018245_1	17.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2018245_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:70107417(-)-4:70173859(-)__4_70094501_70119501D;SPAN=66442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=[chr4:70173859[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	71522256	+	chr4	71527809	+	AGGTCAGACAAATGGTACACAAATCTGGTTCTCAATGGTGAGGTGGGATCAGAGATATTCTCCCTGTTGTTCAGAGGAACA	6	146	2022422_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;INSERTION=AGGTCAGACAAATGGTACACAAATCTGGTTCTCAATGGTGAGGTGGGATCAGAGATATTCTCCCTGTTGTTCAGAGGAACA;MAPQ=60;MATEID=2022422_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_71515501_71540501_347C;SPAN=5553;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:131 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:146 DR:6 LR:-448.9 LO:448.9);ALT=G[chr4:71527809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71522293	+	chr4	71532143	+	.	16	0	2022423_1	23.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2022423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:71522293(+)-4:71532143(-)__4_71515501_71540501D;SPAN=9850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:108 GQ:23.6 PL:[23.6, 0.0, 238.1] SR:0 DR:16 LR:-23.56 LO:33.95);ALT=A[chr4:71532143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71523008	+	chr4	71527809	+	.	2	108	2022424_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=2022424_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_71515501_71540501_347C;SPAN=4801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:108 DP:146 GQ:36.5 PL:[317.0, 0.0, 36.5] SR:108 DR:2 LR:-329.8 LO:329.8);ALT=A[chr4:71527809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71523073	+	chr4	71532143	+	.	71	0	2022425_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=2022425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:71523073(+)-4:71532143(-)__4_71515501_71540501D;SPAN=9070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:98 GQ:29.6 PL:[207.8, 0.0, 29.6] SR:0 DR:71 LR:-215.5 LO:215.5);ALT=G[chr4:71532143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71527935	+	chr4	71532144	+	.	94	21	2022439_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=2022439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_71515501_71540501_247C;SPAN=4209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:112 GQ:30 PL:[330.0, 30.0, 0.0] SR:21 DR:94 LR:-330.1 LO:330.1);ALT=T[chr4:71532144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	71702031	+	chr4	71704944	+	.	5	2	2023320_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2023320_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_71687001_71712001_341C;SPAN=2913;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:2 DR:5 LR:3.764 LO:10.62);ALT=C[chr4:71704944[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	72167580	-	chr5	139946153	+	.	9	0	2596631_1	22.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=2596631_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:72167580(-)-5:139946153(-)__5_139944001_139969001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:0 DR:9 LR:-22.39 LO:22.75);ALT=[chr5:139946153[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	74606473	+	chr4	74607665	+	.	18	0	2032214_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2032214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:74606473(+)-4:74607665(-)__4_74602501_74627501D;SPAN=1192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:104 GQ:31.4 PL:[31.4, 0.0, 219.5] SR:0 DR:18 LR:-31.24 LO:39.53);ALT=T[chr4:74607665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	74719731	-	chr4	74847057	+	.	10	0	2032552_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2032552_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:74719731(-)-4:74847057(-)__4_74700501_74725501D;SPAN=127326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:43 GQ:21.5 PL:[21.5, 0.0, 80.9] SR:0 DR:10 LR:-21.36 LO:23.41);ALT=[chr4:74847057[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	75023999	+	chr4	75027495	+	ACCAGCAGAGAGAAGAGATTCCATCTTCCAG	17	27	2033313_1	87.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACCAGCAGAGAGAAGAGATTCCATCTTCCAG;MAPQ=60;MATEID=2033313_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_75019001_75044001_165C;SPAN=3496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:103 GQ:87.8 PL:[87.8, 0.0, 160.4] SR:27 DR:17 LR:-87.63 LO:88.85);ALT=G[chr4:75027495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	75023999	+	chr4	75025770	+	.	34	25	2033312_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2033312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_75019001_75044001_219C;SPAN=1771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:135 GQ:99 PL:[115.4, 0.0, 211.1] SR:25 DR:34 LR:-115.3 LO:116.8);ALT=G[chr4:75025770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	75144496	+	chr4	75195914	+	.	0	11	2033854_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2033854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_75190501_75215501_262C;SPAN=51418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:11 DR:0 LR:-24.12 LO:26.03);ALT=C[chr4:75195914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	75642738	+	chr4	75648840	+	.	21	0	2035366_1	50.0	.	DISC_MAPQ=11;EVDNC=DSCRD;IMPRECISE;MAPQ=11;MATEID=2035366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:75642738(+)-4:75648840(-)__4_75631501_75656501D;SPAN=6102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:72 GQ:50 PL:[50.0, 0.0, 122.6] SR:0 DR:21 LR:-49.81 LO:51.6);ALT=G[chr4:75648840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	76434508	+	chr4	76439406	+	.	8	5	2037246_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2037246_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_76415501_76440501_288C;SPAN=4898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:5 DR:8 LR:-0.7201 LO:16.74);ALT=T[chr4:76439406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	76582914	+	chr4	76587113	+	ATTTTGGCCATAAACAGCTTCCTGGGGCTTTCCACTAGCATCTACTCCACCATGAACATAGGAAGAATTCCTGCCATAAA	0	24	2037813_1	49.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=ATTTTGGCCATAAACAGCTTCCTGGGGCTTTCCACTAGCATCTACTCCACCATGAACATAGGAAGAATTCCTGCCATAAA;MAPQ=60;MATEID=2037813_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_76562501_76587501_171C;SPAN=4199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:110 GQ:49.4 PL:[49.4, 0.0, 217.7] SR:24 DR:0 LR:-49.42 LO:55.42);ALT=C[chr4:76587113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	76584111	+	chr4	76587113	+	.	0	19	2037895_1	48.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=2037895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_76587001_76612001_441C;SPAN=3002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:52 GQ:48.8 PL:[48.8, 0.0, 75.2] SR:19 DR:0 LR:-48.63 LO:48.99);ALT=G[chr4:76587113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	76587235	+	chr4	76598392	+	.	0	33	2037899_1	76.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2037899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_76587001_76612001_83C;SPAN=11157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:122 GQ:76.1 PL:[76.1, 0.0, 218.0] SR:33 DR:0 LR:-75.88 LO:79.79);ALT=T[chr4:76598392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	76903192	+	chr4	76911905	+	.	0	14	2039269_1	33.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2039269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_76881001_76906001_434C;SPAN=8713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:48 GQ:33.2 PL:[33.2, 0.0, 82.7] SR:14 DR:0 LR:-33.21 LO:34.4);ALT=T[chr4:76911905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77265746	-	chr20	17949054	+	.	9	0	6942896_1	11.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6942896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:77265746(-)-20:17949054(-)__20_17934001_17959001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=[chr20:17949054[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	77871083	+	chr4	77917578	+	.	19	17	2042830_1	69.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=2042830_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_77910001_77935001_357C;SPAN=46495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:60 GQ:69.5 PL:[69.5, 0.0, 76.1] SR:17 DR:19 LR:-69.57 LO:69.59);ALT=T[chr4:77917578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77917694	+	chr4	77926753	+	.	2	8	2042857_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2042857_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_77910001_77935001_95C;SPAN=9059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:119 GQ:0.8 PL:[0.8, 0.0, 287.9] SR:8 DR:2 LR:-0.77 LO:18.6);ALT=T[chr4:77926753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77933076	+	chr4	77936007	+	.	3	5	2042903_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2042903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_77910001_77935001_375C;SPAN=2931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:48 GQ:3.5 PL:[3.5, 0.0, 112.4] SR:5 DR:3 LR:-3.501 LO:9.789);ALT=T[chr4:77936007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77936172	+	chr4	77940318	+	.	0	9	2042759_1	0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=2042759_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_77934501_77959501_327C;SPAN=4146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:108 GQ:0.5 PL:[0.5, 0.0, 261.2] SR:9 DR:0 LR:-0.4492 LO:16.7);ALT=T[chr4:77940318[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77940414	+	chr4	77941654	+	.	2	16	2042776_1	24.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2042776_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_4_77934501_77959501_256C;SPAN=1240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:129 GQ:24.5 PL:[24.5, 0.0, 288.5] SR:16 DR:2 LR:-24.47 LO:37.69);ALT=G[chr4:77941654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77940414	+	chr4	77949780	+	TTGAGAATGAAAATCATTGCGATTTTGTGAAACTTCGAGAGATGCTGATCCGCGTGAACATGGAGGACTTGCGAGAGCAGACTCACACCCGCCACTATGAATTGTACCGACGCTGTAAGCTTGAAGAGATGGGGTTCAAGGACACTGACCCTGACAGCAAACCCTTC	0	26	2042777_1	52.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTGAGAATGAAAATCATTGCGATTTTGTGAAACTTCGAGAGATGCTGATCCGCGTGAACATGGAGGACTTGCGAGAGCAGACTCACACCCGCCACTATGAATTGTACCGACGCTGTAAGCTTGAAGAGATGGGGTTCAAGGACACTGACCCTGACAGCAAACCCTTC;MAPQ=60;MATEID=2042777_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_77934501_77959501_256C;SPAN=9366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:124 GQ:52.4 PL:[52.4, 0.0, 247.1] SR:26 DR:0 LR:-52.23 LO:59.53);ALT=G[chr4:77949780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77969818	+	chr4	77976303	+	.	17	19	2043206_1	76.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2043206_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_77959001_77984001_199C;SPAN=6485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:121 GQ:76.4 PL:[76.4, 0.0, 215.0] SR:19 DR:17 LR:-76.15 LO:79.93);ALT=G[chr4:77976303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77977257	+	chr4	77979659	+	CATCTTCCTCAACAGTCTTGGCAGCTAGGAAAAAACAGCTGATTGCAATACAACTCAAGTATTTTGGATGAG	3	14	2043228_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CATCTTCCTCAACAGTCTTGGCAGCTAGGAAAAAACAGCTGATTGCAATACAACTCAAGTATTTTGGATGAG;MAPQ=60;MATEID=2043228_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_77959001_77984001_188C;SPAN=2402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:99 GQ:29.3 PL:[29.3, 0.0, 210.8] SR:14 DR:3 LR:-29.3 LO:37.27);ALT=T[chr4:77979659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77979790	+	chr4	77987402	+	.	6	4	2043262_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2043262_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_77983501_78008501_381C;SPAN=7612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:4 DR:6 LR:-15.35 LO:19.68);ALT=T[chr4:77987402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	77987566	+	chr4	77996651	+	.	17	0	2043281_1	27.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2043281_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:77987566(+)-4:77996651(-)__4_77983501_78008501D;SPAN=9085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:105 GQ:27.8 PL:[27.8, 0.0, 225.8] SR:0 DR:17 LR:-27.67 LO:36.79);ALT=A[chr4:77996651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	78179079	-	chr4	79035861	+	.	13	0	2046744_1	26.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=2046744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:78179079(-)-4:79035861(-)__4_79012501_79037501D;SPAN=856782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:61 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.39 LO:29.87);ALT=[chr4:79035861[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	78695905	+	chr4	78740439	+	.	10	0	2045425_1	20.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2045425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:78695905(+)-4:78740439(-)__4_78694001_78719001D;SPAN=44534;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:0 DR:10 LR:-20.28 LO:22.97);ALT=C[chr4:78740439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	78784126	+	chr4	78804395	+	.	13	0	2045964_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2045964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:78784126(+)-4:78804395(-)__4_78767501_78792501D;SPAN=20269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:67 GQ:24.8 PL:[24.8, 0.0, 137.0] SR:0 DR:13 LR:-24.76 LO:29.27);ALT=A[chr4:78804395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	78793011	+	chr4	78804396	+	.	0	8	2045811_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=2045811_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_78792001_78817001_222C;SPAN=11385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-2.025 LO:15.08);ALT=T[chr4:78804396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	79269134	+	chr4	79275196	+	.	56	15	2047479_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAGCTTCAAGATA;MAPQ=60;MATEID=2047479_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_79257501_79282501_431C;SPAN=6062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:199 GQ:99 PL:[154.1, 0.0, 329.0] SR:15 DR:56 LR:-154.1 LO:157.5);ALT=A[chr4:79275196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	49282763	+	chr4	79750908	+	.	3	24	2048995_1	74.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=TCTTTTCTTTTCTTTTCTTTTCTTTT;MAPQ=0;MATEID=2048995_2;MATENM=6;NM=1;NUMPARTS=2;SCTG=c_4_79747501_79772501_344C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:41 GQ:22.1 PL:[74.9, 0.0, 22.1] SR:24 DR:3 LR:-76.1 LO:76.1);ALT=]chr20:49282763]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	83196114	-	chr12	51717804	+	.	54	4	2059126_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;HOMSEQ=ACCTTCTCCTGGGCCCTGCT;MAPQ=43;MATEID=2059126_2;MATENM=0;NM=7;NUMPARTS=2;SCTG=c_4_83177501_83202501_264C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:57 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:4 DR:54 LR:-171.6 LO:171.6);ALT=[chr12:51717804[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	83275310	+	chr4	83276455	+	.	11	16	2059441_1	68.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=44;MATEID=2059441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83251001_83276001_282C;SPAN=1145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:66 GQ:68 PL:[68.0, 0.0, 91.1] SR:16 DR:11 LR:-67.95 LO:68.15);ALT=G[chr4:83276455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83276554	+	chr4	83277690	+	.	2	9	2059458_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2059458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83275501_83300501_76C;SPAN=1136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:127 GQ:1.2 PL:[0.0, 1.2, 310.2] SR:9 DR:2 LR:1.397 LO:18.3);ALT=T[chr4:83277690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83276555	+	chr4	83277949	+	.	0	14	2059459_1	11.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2059459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83275501_83300501_108C;SPAN=1394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:127 GQ:11.9 PL:[11.9, 0.0, 295.7] SR:14 DR:0 LR:-11.81 LO:27.77);ALT=C[chr4:83277949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83280793	+	chr4	83292680	+	.	3	15	2059476_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=2059476_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTCTTC;SCTG=c_4_83275501_83300501_305C;SPAN=11887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:107 GQ:18 PL:[18.0, 0.0, 174.0] SR:15 DR:3 LR:-17.85 LO:26.76);ALT=C[chr4:83292680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83280793	+	chr4	83294599	+	ATTCTTCCCGCTGTGCCGTCGCTGCTTCAGAGTGTCGTGGGGAGGAGTTTGAATGG	0	28	2059477_1	57.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATTCTTCCCGCTGTGCCGTCGCTGCTTCAGAGTGTCGTGGGGAGGAGTTTGAATGG;MAPQ=60;MATEID=2059477_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_83275501_83300501_305C;SPAN=13806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:131 GQ:57.2 PL:[57.2, 0.0, 258.5] SR:28 DR:0 LR:-56.94 LO:64.37);ALT=C[chr4:83294599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83292738	+	chr4	83294599	+	.	7	13	2059532_1	32.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2059532_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_4_83275501_83300501_305C;SPAN=1861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:126 GQ:32 PL:[32.0, 0.0, 272.9] SR:13 DR:7 LR:-31.88 LO:43.09);ALT=C[chr4:83294599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83323608	+	chrX	69353870	-	.	8	0	7443254_1	19.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7443254_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:83323608(+)-23:69353870(+)__23_69335001_69360001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:27 GQ:19.1 PL:[19.1, 0.0, 45.5] SR:0 DR:8 LR:-19.09 LO:19.72);ALT=A]chrX:69353870];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	83352067	+	chr4	83369071	+	.	4	4	2059685_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2059685_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83349001_83374001_368C;SPAN=17004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:4 DR:4 LR:-0.6702 LO:14.89);ALT=G[chr4:83369071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83616163	+	chr5	134263298	+	AAC	33	18	2060658_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AAC;MAPQ=60;MATEID=2060658_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_83594001_83619001_229C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:58 GQ:0.8 PL:[139.4, 0.0, 0.8] SR:18 DR:33 LR:-147.8 LO:147.8);ALT=C[chr5:134263298[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	83740406	+	chr4	83742190	+	.	0	7	2061292_1	9.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2061292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83741001_83766001_395C;SPAN=1784;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:50 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:7 DR:0 LR:-9.561 LO:14.67);ALT=G[chr4:83742190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83800083	+	chr4	83801949	+	.	3	5	2061879_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TACCT;MAPQ=60;MATEID=2061879_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_83790001_83815001_14C;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:5 DR:3 LR:0.4135 LO:14.74);ALT=T[chr4:83801949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83800083	+	chr4	83803010	+	GTGAGAAGAGGAGAATGTGGCACAAGATTTCATATCCAAGGATGGATCAGAGAGGTCTAATTCAAATATCTCAAGGGAAGCATTCGTACTAAATGTTGCATCCAATTGCTGAGCAGATGTT	0	28	2061880_1	63.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GTGAGAAGAGGAGAATGTGGCACAAGATTTCATATCCAAGGATGGATCAGAGAGGTCTAATTCAAATATCTCAAGGGAAGCATTCGTACTAAATGTTGCATCCAATTGCTGAGCAGATGTT;MAPQ=60;MATEID=2061880_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_83790001_83815001_14C;SPAN=2927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:106 GQ:63.8 PL:[63.8, 0.0, 192.5] SR:28 DR:0 LR:-63.71 LO:67.36);ALT=T[chr4:83803010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83802115	+	chr4	83812239	+	.	13	0	2061892_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2061892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:83802115(+)-4:83812239(-)__4_83790001_83815001D;SPAN=10124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=T[chr4:83812239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83923136	-	chr17	7644589	+	T	4	19	2062014_1	58.0	.	DISC_MAPQ=47;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=2062014_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_83912501_83937501_7C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:27 GQ:5.9 PL:[58.7, 0.0, 5.9] SR:19 DR:4 LR:-61.09 LO:61.09);ALT=[chr17:7644589[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	83956452	+	chr4	83970316	+	.	15	0	2062496_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2062496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:83956452(+)-4:83970316(-)__4_83961501_83986501D;SPAN=13864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:56 GQ:34.4 PL:[34.4, 0.0, 100.4] SR:0 DR:15 LR:-34.34 LO:36.19);ALT=G[chr4:83970316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	83956453	+	chr4	83966779	+	.	12	4	2062497_1	35.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=2062497_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_83961501_83986501_145C;SPAN=10326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:41 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:4 DR:12 LR:-35.11 LO:35.58);ALT=T[chr4:83966779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84015944	+	chr4	84026048	+	.	3	64	2062180_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=C;MAPQ=18;MATEID=2062180_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_84010501_84035501_305C;SPAN=10104;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:126 GQ:99 PL:[183.8, 0.0, 121.1] SR:64 DR:3 LR:-184.4 LO:184.4);ALT=C[chr4:84026048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84015973	+	chr4	84035816	+	.	14	0	2062619_1	32.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=2062619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84015973(+)-4:84035816(-)__4_84035001_84060001D;SPAN=19843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:53 GQ:32 PL:[32.0, 0.0, 94.7] SR:0 DR:14 LR:-31.86 LO:33.68);ALT=T[chr4:84035816[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84026173	+	chr4	84028955	+	.	0	74	2062228_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=25;MATEID=2062228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_84010501_84035501_330C;SPAN=2782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:74 DP:115 GQ:64.7 PL:[213.2, 0.0, 64.7] SR:74 DR:0 LR:-217.4 LO:217.4);ALT=C[chr4:84028955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84026199	+	chr4	84035817	+	.	50	0	2062620_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=2062620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84026199(+)-4:84035817(-)__4_84035001_84060001D;SPAN=9618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:50 LR:-161.7 LO:161.7);ALT=T[chr4:84035817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84029103	+	chr4	84035819	+	.	84	10	2062621_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;MAPQ=60;MATEID=2062621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_84035001_84060001_125C;SPAN=6716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:61 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:10 DR:84 LR:-250.9 LO:250.9);ALT=A[chr4:84035819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	132611296	+	chr4	84035816	+	.	65	0	5400324_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5400324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84035816(-)-12:132611296(+)__12_132594001_132619001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:36 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=]chr12:132611296]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	84200268	+	chr4	84205664	+	.	0	8	2062953_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2062953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_84182001_84207001_261C;SPAN=5396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:126 GQ:7.5 PL:[0.0, 7.5, 320.1] SR:8 DR:0 LR:7.729 LO:13.87);ALT=C[chr4:84205664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	84377306	+	chrX	53852543	+	.	17	0	7426485_1	49.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=7426485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84377306(+)-23:53852543(-)__23_53851001_53876001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:26 GQ:12.8 PL:[49.1, 0.0, 12.8] SR:0 DR:17 LR:-50.15 LO:50.15);ALT=C[chrX:53852543[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	84377323	+	chr4	84379497	+	.	10	0	2063857_1	17.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=2063857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:84377323(+)-4:84379497(-)__4_84353501_84378501D;SPAN=2174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=T[chr4:84379497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	85719024	+	chr12	7830042	+	.	0	39	2068113_1	99.0	.	EVDNC=ASSMB;HOMSEQ=T;MAPQ=60;MATEID=2068113_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_85701001_85726001_290C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:59 GQ:30.2 PL:[112.7, 0.0, 30.2] SR:39 DR:0 LR:-115.4 LO:115.4);ALT=T[chr12:7830042[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	87854696	+	chr4	87857140	+	.	4	2	2074710_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2074710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_87832501_87857501_117C;SPAN=2444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:94 GQ:12 PL:[0.0, 12.0, 250.8] SR:2 DR:4 LR:12.26 LO:6.224);ALT=T[chr4:87857140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88258520	+	chr4	88261641	+	.	0	8	2076610_1	2.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2076610_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_4_88249001_88274001_337C;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:8 DR:0 LR:-2.567 LO:15.16);ALT=T[chr4:88261641[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88258520	+	chr4	88278431	+	TTCCAATGTTGTTAAAAAAGCTATAGAAGATGGAATAAAAATCATCTTCTGCTCAGTCAGAATCCCATGCATCAGCCTGTTTACCACTTCCTCAGGTTCCAGAGTGGGTCCCAAA	6	14	2076611_1	42.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTCCAATGTTGTTAAAAAAGCTATAGAAGATGGAATAAAAATCATCTTCTGCTCAGTCAGAATCCCATGCATCAGCCTGTTTACCACTTCCTCAGGTTCCAGAGTGGGTCCCAAA;MAPQ=60;MATEID=2076611_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_4_88249001_88274001_337C;SPAN=19911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:51 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:14 DR:6 LR:-42.3 LO:42.98);ALT=T[chr4:88278431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88261760	+	chr4	88278431	+	.	3	6	2076168_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2076168_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_88273501_88298501_240C;SPAN=16671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:6 DR:3 LR:-14.54 LO:19.45);ALT=T[chr4:88278431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88303516	+	chr4	88312013	+	.	35	67	2076300_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2076300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_88298001_88323001_247C;SPAN=8497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:127 GQ:87.8 PL:[219.8, 0.0, 87.8] SR:67 DR:35 LR:-222.8 LO:222.8);ALT=T[chr4:88312013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88483900	+	chr4	88486313	+	.	88	56	2077334_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAGTTACAAACAAC;MAPQ=60;MATEID=2077334_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_88469501_88494501_334C;SPAN=2413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:51 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:56 DR:88 LR:-340.0 LO:340.0);ALT=C[chr4:88486313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	88847164	-	chr4	88858700	+	A	115	69	2078496_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=2078496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_88837001_88862001_254C;SPAN=11536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:68 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:69 DR:115 LR:-458.8 LO:458.8);ALT=[chr4:88858700[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	89443200	+	chr4	89444795	+	.	17	0	2080374_1	25.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2080374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:89443200(+)-4:89444795(-)__4_89425001_89450001D;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:113 GQ:25.7 PL:[25.7, 0.0, 246.8] SR:0 DR:17 LR:-25.5 LO:36.2);ALT=A[chr4:89444795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	93570162	+	chr4	93567358	+	TTGAACAAGTTCAATTTAAAATATTTCATAAGCTTGTATGATATCATTGGGGCTAGAGTAGACGTGATACTAAATGTAGGAAATAAATGGAATAAACACTCAGAGAGGAACTATATGTTTTGTCTTAAAACTTCATTAAGTCTAAGAATTGATATTTTGTTGCTGGATGAATTGGTGGTTTGTGAGTTATAGTGAATATATCTCCCTGTTACATTCCTGTCGTTGTCCTATCCATTGTCCTATTGTTGGATGTTTCACTTGTATATCCCATGTTACATAATTTTATCATAGAGAGCAAAAGAATTTGACTACAGTAAACTTAATGCTTTGCCATGTACAGATGTATGACAAAGAACATGTTATTTTGAAAGTTTTTGCTCTTATATTTTCTTTGCAGTCTGACTTCTTAATATTTGCTTCATTTTCATGTATGTGTTTTTACAAAGCATTCTCTTGGTATCACTAACCAAATACCTGTTTAGAGAAACAAAAGGCCAACTGGGGATGAAAACAGTTTATTTACTTACTGCACAGTATG	2	147	2092253_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTGAACAAGTTCAATTTAAAATATTTCATAAGCTTGTATGATATCATTGGGGCTAGAGTAGACGTGATACTAAATGTAGGAAATAAATGGAATAAACACTCAGAGAGGAACTATATGTTTTGTCTTAAAACTTCATTAAGTCTAAGAATTGATATTTTGTTGCTGGATGAATTGGTGGTTTGTGAGTTATAGTGAATATATCTCCCTGTTACATTCCTGTCGTTGTCCTATCCATTGTCCTATTGTTGGATGTTTCACTTGTATATCCCATGTTACATAATTTTATCATAGAGAGCAAAAGAATTTGACTACAGTAAACTTAATGCTTTGCCATGTACAGATGTATGACAAAGAACATGTTATTTTGAAAGTTTTTGCTCTTATATTTTCTTTGCAGTCTGACTTCTTAATATTTGCTTCATTTTCATGTATGTGTTTTTACAAAGCATTCTCTTGGTATCACTAACCAAATACCTGTTTAGAGAAACAAAAGGCCAACTGGGGATGAAAACAGTTTATTTACTTACTGCACAGTATG;MAPQ=60;MATEID=2092253_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_93565501_93590501_297C;SPAN=2804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:148 DP:95 GQ:40 PL:[439.0, 40.0, 0.0] SR:147 DR:2 LR:-439.0 LO:439.0);ALT=]chr4:93570162]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	94559454	+	chr4	94565491	+	.	107	64	2094967_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAAAACTTGCATCTT;MAPQ=60;MATEID=2094967_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_94545501_94570501_233C;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:46 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:64 DR:107 LR:-399.4 LO:399.4);ALT=T[chr4:94565491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	95373180	+	chr4	95444874	+	.	8	0	2097562_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2097562_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:95373180(+)-4:95444874(-)__4_95427501_95452501D;SPAN=71694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=G[chr4:95444874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	95518746	+	chr7	46904659	+	.	95	84	3290388_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAGCC;MAPQ=60;MATEID=3290388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_46893001_46918001_396C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:45 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:84 DR:95 LR:-432.4 LO:432.4);ALT=C[chr7:46904659[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	99678413	-	chr4	99679873	+	.	8	0	2109815_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2109815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:99678413(-)-4:99679873(-)__4_99666001_99691001D;SPAN=1460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:104 GQ:1.5 PL:[0.0, 1.5, 254.1] SR:0 DR:8 LR:1.768 LO:14.56);ALT=[chr4:99679873[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	99917041	+	chr4	99955380	+	.	9	0	2110768_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2110768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:99917041(+)-4:99955380(-)__4_99911001_99936001D;SPAN=38339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:0 DR:9 LR:-21.04 LO:21.94);ALT=A[chr4:99955380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	100003277	+	chr4	100009837	+	.	10	0	2111367_1	18.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=2111367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:100003277(+)-4:100009837(-)__4_100009001_100034001D;SPAN=6560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:54 GQ:18.5 PL:[18.5, 0.0, 110.9] SR:0 DR:10 LR:-18.38 LO:22.29);ALT=C[chr4:100009837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	100806874	+	chr4	100815490	+	.	8	0	2113577_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=2113577_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:100806874(+)-4:100815490(-)__4_100793001_100818001D;SPAN=8616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:99 GQ:0.3 PL:[0.0, 0.3, 240.9] SR:0 DR:8 LR:0.4135 LO:14.74);ALT=A[chr4:100815490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	100870127	+	chr4	100871361	+	.	23	0	2113964_1	50.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2113964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:100870127(+)-4:100871361(-)__4_100866501_100891501D;SPAN=1234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:95 GQ:50.3 PL:[50.3, 0.0, 179.0] SR:0 DR:23 LR:-50.19 LO:54.31);ALT=C[chr4:100871361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	71016305	+	chr4	100871369	+	.	26	0	2113973_1	43.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2113973_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:100871369(-)-8:71016305(+)__4_100866501_100891501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:158 GQ:43.1 PL:[43.1, 0.0, 340.1] SR:0 DR:26 LR:-43.02 LO:56.47);ALT=]chr8:71016305]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr18	5227885	+	chr4	101860821	+	.	0	10	2116717_1	21.0	.	EVDNC=ASSMB;HOMSEQ=ACATCACTAATT;MAPQ=60;MATEID=2116717_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_4_101846501_101871501_283C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:10 DR:0 LR:-21.63 LO:23.53);ALT=]chr18:5227885]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	102336327	+	chr20	47019890	+	.	10	30	7039494_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;HOMSEQ=GAAGGAAGGAAGGAAG;MAPQ=53;MATEID=7039494_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_47015501_47040501_290C;SPAN=-1;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:20 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:30 DR:10 LR:-115.5 LO:115.5);ALT=G[chr20:47019890[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	5273545	+	chr4	103748338	+	.	57	0	2122682_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2122682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:103748338(-)-20:5273545(+)__4_103733001_103758001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:93 GQ:60.8 PL:[163.1, 0.0, 60.8] SR:0 DR:57 LR:-165.4 LO:165.4);ALT=]chr20:5273545]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr4	103790344	+	chr4	103806371	+	.	0	24	2122482_1	47.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2122482_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_103782001_103807001_362C;SPAN=16027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:117 GQ:47.6 PL:[47.6, 0.0, 235.7] SR:24 DR:0 LR:-47.53 LO:54.69);ALT=G[chr4:103806371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	103790566	+	chr4	103806406	+	.	25	0	2122903_1	72.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2122903_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:103790566(+)-4:103806406(-)__4_103806501_103831501D;SPAN=15840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:2 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:0 DR:25 LR:-72.62 LO:72.62);ALT=G[chr4:103806406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	104316046	-	chr4	104317168	+	.	9	0	2124344_1	4.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=2124344_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:104316046(-)-4:104317168(-)__4_104296501_104321501D;SPAN=1122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:0 DR:9 LR:-3.971 LO:17.23);ALT=[chr4:104317168[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	106290912	+	chr4	106307721	+	TCTTCATTACTTTCTTTATTTGGTGAAGATGA	3	37	2129852_1	99.0	.	DISC_MAPQ=40;EVDNC=TSI_G;HOMSEQ=TACC;INSERTION=TCTTCATTACTTTCTTTATTTGGTGAAGATGA;MAPQ=60;MATEID=2129852_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_106281001_106306001_46C;SPAN=16809;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:45 GQ:5.4 PL:[118.8, 5.4, 0.0] SR:37 DR:3 LR:-121.4 LO:121.4);ALT=T[chr4:106307721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106317493	+	chr4	106320193	+	.	3	8	2130034_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2130034_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_106305501_106330501_61C;SPAN=2700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:80 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:8 DR:3 LR:-4.734 LO:15.51);ALT=T[chr4:106320193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106345483	+	chr4	106359107	+	.	3	6	2130296_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTTT;MAPQ=60;MATEID=2130296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_106354501_106379501_149C;SPAN=13624;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:6 DR:3 LR:-15.08 LO:19.6);ALT=T[chr4:106359107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106367661	+	chr4	106370507	+	.	2	16	2130334_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2130334_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_106354501_106379501_129C;SPAN=2846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:106 GQ:30.8 PL:[30.8, 0.0, 225.5] SR:16 DR:2 LR:-30.7 LO:39.37);ALT=T[chr4:106370507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106367661	+	chr4	106374755	+	CCATTTTAGCATTTGTCCACCGAGGTATTTCTACAATCATATTAAACAGATT	3	26	2130335_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCATTTTAGCATTTGTCCACCGAGGTATTTCTACAATCATATTAAACAGATT;MAPQ=60;MATEID=2130335_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_106354501_106379501_129C;SPAN=7094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:109 GQ:62.9 PL:[62.9, 0.0, 201.5] SR:26 DR:3 LR:-62.9 LO:66.96);ALT=T[chr4:106374755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106370608	+	chr4	106395094	+	.	8	0	2130348_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2130348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:106370608(+)-4:106395094(-)__4_106354501_106379501D;SPAN=24486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=T[chr4:106395094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106377956	+	chr4	106395145	+	.	13	0	2130371_1	30.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2130371_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:106377956(+)-4:106395145(-)__4_106354501_106379501D;SPAN=17189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:46 GQ:30.5 PL:[30.5, 0.0, 80.0] SR:0 DR:13 LR:-30.45 LO:31.73);ALT=G[chr4:106395145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	106482669	-	chr8	111740547	+	.	10	0	4023193_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4023193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:106482669(-)-8:111740547(-)__8_111720001_111745001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=[chr8:111740547[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	107056578	+	chr4	107063363	+	CA	32	33	2132529_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CA;MAPQ=60;MATEID=2132529_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_107040501_107065501_326C;SPAN=6785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:51 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:33 DR:32 LR:-148.5 LO:148.5);ALT=C[chr4:107063363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107237794	+	chr4	107248607	+	.	42	0	2133059_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2133059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107237794(+)-4:107248607(-)__4_107236501_107261501D;SPAN=10813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:105 GQ:99 PL:[110.3, 0.0, 143.3] SR:0 DR:42 LR:-110.2 LO:110.5);ALT=T[chr4:107248607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107237795	+	chr4	107246141	+	.	19	0	2133060_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2133060_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107237795(+)-4:107246141(-)__4_107236501_107261501D;SPAN=8346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:89 GQ:38.6 PL:[38.6, 0.0, 177.2] SR:0 DR:19 LR:-38.61 LO:43.67);ALT=T[chr4:107246141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107246275	+	chr4	107248608	+	.	2	53	2133083_1	99.0	.	DISC_MAPQ=28;EVDNC=ASDIS;MAPQ=60;MATEID=2133083_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_107236501_107261501_66C;SPAN=2333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:102 GQ:94.7 PL:[150.8, 0.0, 94.7] SR:53 DR:2 LR:-151.2 LO:151.2);ALT=A[chr4:107248608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107249443	+	chr4	107252848	+	.	10	0	2133092_1	3.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2133092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107249443(+)-4:107252848(-)__4_107236501_107261501D;SPAN=3405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:111 GQ:3.2 PL:[3.2, 0.0, 263.9] SR:0 DR:10 LR:-2.937 LO:18.91);ALT=T[chr4:107252848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	107317322	-	chr4	107320347	+	.	15	0	2132923_1	24.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=2132923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:107317322(-)-4:107320347(-)__4_107310001_107335001D;SPAN=3025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:94 GQ:24.2 PL:[24.2, 0.0, 202.4] SR:0 DR:15 LR:-24.05 LO:32.36);ALT=[chr4:107320347[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	108127828	+	chr4	108131715	+	.	93	61	2135501_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AAAACATTAGGATTCTCTTT;MAPQ=60;MATEID=2135501_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108118501_108143501_113C;SPAN=3887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:127 DP:34 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:61 DR:93 LR:-376.3 LO:376.3);ALT=T[chr4:108131715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108276701	+	chr4	108279505	+	.	61	66	2135779_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAC;MAPQ=60;MATEID=2135779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108265501_108290501_170C;SPAN=2804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:41 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:66 DR:61 LR:-310.3 LO:310.3);ALT=C[chr4:108279505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108615164	+	chr4	108622326	+	.	0	13	2136741_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2136741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108608501_108633501_339C;SPAN=7162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:105 GQ:14.6 PL:[14.6, 0.0, 239.0] SR:13 DR:0 LR:-14.47 LO:26.49);ALT=T[chr4:108622326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108615204	+	chr4	108641277	+	.	13	0	2137019_1	30.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2137019_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:108615204(+)-4:108641277(-)__4_108633001_108658001D;SPAN=26073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:46 GQ:30.5 PL:[30.5, 0.0, 80.0] SR:0 DR:13 LR:-30.45 LO:31.73);ALT=G[chr4:108641277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108622442	+	chr4	108641275	+	.	14	6	2137020_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2137020_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_4_108633001_108658001_275C;SPAN=18833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:47 GQ:40.1 PL:[40.1, 0.0, 73.1] SR:6 DR:14 LR:-40.08 LO:40.64);ALT=C[chr4:108641275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108911222	+	chr4	108930913	+	.	24	25	2137794_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2137794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108927001_108952001_159C;SPAN=19691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:70 GQ:56.9 PL:[113.0, 0.0, 56.9] SR:25 DR:24 LR:-114.1 LO:114.1);ALT=T[chr4:108930913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	108931038	+	chr4	108935585	+	CTA	0	13	2137806_1	17.0	.	EVDNC=ASSMB;INSERTION=CTA;MAPQ=60;MATEID=2137806_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_108927001_108952001_295C;SPAN=4547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:96 GQ:17 PL:[17.0, 0.0, 215.0] SR:13 DR:0 LR:-16.9 LO:27.04);ALT=C[chr4:108935585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	109397798	+	chr12	1115362	+	.	24	0	5065390_1	69.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=5065390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:109397798(+)-12:1115362(-)__12_1102501_1127501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:36 GQ:16.7 PL:[69.5, 0.0, 16.7] SR:0 DR:24 LR:-71.17 LO:71.17);ALT=G[chr12:1115362[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	109571889	+	chr4	109578602	+	.	17	0	2140289_1	21.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2140289_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:109571889(+)-4:109578602(-)__4_109564001_109589001D;SPAN=6713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:127 GQ:21.8 PL:[21.8, 0.0, 285.8] SR:0 DR:17 LR:-21.71 LO:35.26);ALT=C[chr4:109578602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	109571951	+	chr4	109576718	+	.	0	85	2140290_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=27;MATEID=2140290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_109564001_109589001_286C;SPAN=4767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:134 GQ:79.4 PL:[244.4, 0.0, 79.4] SR:85 DR:0 LR:-248.8 LO:248.8);ALT=G[chr4:109576718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	109578804	+	chr4	109588403	+	.	9	18	2140318_1	61.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=G;MAPQ=15;MATEID=2140318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_109564001_109589001_57C;SPAN=9599;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:102 GQ:61.7 PL:[61.7, 0.0, 183.8] SR:18 DR:9 LR:-61.49 LO:64.98);ALT=G[chr4:109588403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115437012	-	chr10	72451334	+	.	11	0	4625756_1	29.0	.	DISC_MAPQ=8;EVDNC=DSCRD;IMPRECISE;MAPQ=8;MATEID=4625756_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:115437012(-)-10:72451334(-)__10_72446501_72471501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:8 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:11 LR:-29.71 LO:29.71);ALT=[chr10:72451334[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	115507821	+	chr4	115511041	+	.	12	45	2158820_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2158820_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_4_115493001_115518001_217C;SPAN=3220;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:69 GQ:27.5 PL:[139.7, 0.0, 27.5] SR:45 DR:12 LR:-144.0 LO:144.0);ALT=G[chr4:115511041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115507821	+	chr4	115513865	+	TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT	33	61	2158821_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TAACCCTTTATACCCTTTAGTCCAGAAAGGCATATTTGGCTTTAGTATTGTCAGGTTGAGT;MAPQ=60;MATEID=2158821_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_115493001_115518001_217C;SPAN=6044;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:66 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:61 DR:33 LR:-241.0 LO:241.0);ALT=G[chr4:115513865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115511096	+	chr4	115513865	+	GTTGAGT	12	33	2158823_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=AG;INSERTION=GTTGAGT;MAPQ=44;MATEID=2158823_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_4_115493001_115518001_217C;SPAN=2769;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:76 GQ:75.2 PL:[108.2, 0.0, 75.2] SR:33 DR:12 LR:-108.4 LO:108.4);ALT=G[chr4:115513865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	115928723	+	chr4	115931874	+	.	48	36	2160360_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GTGA;MAPQ=60;MATEID=2160360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_115909501_115934501_351C;SPAN=3151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:61 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:36 DR:48 LR:-201.3 LO:201.3);ALT=A[chr4:115931874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	130066137	+	chr4	130068441	+	.	10	0	2204511_1	29.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2204511_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:130066137(+)-4:130068441(-)__4_130046001_130071001D;SPAN=2304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:13 GQ:0 PL:[29.7, 0.0, 0.0] SR:0 DR:10 LR:-30.9 LO:30.9);ALT=A[chr4:130068441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	130961892	+	chr4	131004550	+	CCT	60	55	2206992_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCT;MAPQ=60;MATEID=2206992_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_131001501_131026501_192C;SPAN=42658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:48 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:55 DR:60 LR:-274.0 LO:274.0);ALT=C[chr4:131004550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	135363636	-	chr15	77180305	+	.	8	0	5993869_1	18.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=5993869_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:135363636(-)-15:77180305(-)__15_77175001_77200001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=[chr15:77180305[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	135433002	+	chr4	135435702	+	GTACA	13	62	2220961_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GTACA;MAPQ=60;MATEID=2220961_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_4_135411501_135436501_126C;SPAN=2700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:61 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:62 DR:13 LR:-217.9 LO:217.9);ALT=A[chr4:135435702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	138966211	+	chr4	138967219	+	T	49	30	2231112_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=2231112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_138964001_138989001_336C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:63 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:30 DR:49 LR:-184.8 LO:184.8);ALT=G[chr4:138967219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	139482000	-	chr16	69788760	+	.	12	0	6240889_1	30.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=6240889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:139482000(-)-16:69788760(-)__16_69776001_69801001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:0 DR:12 LR:-30.4 LO:30.71);ALT=[chr16:69788760[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	139994722	+	chr4	140005295	+	GGCCCGG	0	11	2234527_1	4.0	.	EVDNC=ASSMB;INSERTION=GGCCCGG;MAPQ=60;MATEID=2234527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_139993001_140018001_186C;SPAN=10573;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:119 GQ:4.1 PL:[4.1, 0.0, 284.6] SR:11 DR:0 LR:-4.071 LO:20.93);ALT=C[chr4:140005295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140211246	+	chr4	140213681	+	.	2	29	2235527_1	87.0	.	DISC_MAPQ=30;EVDNC=TSI_L;HOMSEQ=TAC;MAPQ=60;MATEID=2235527_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_140213501_140238501_347C;SPAN=2435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:42 GQ:11.9 PL:[87.8, 0.0, 11.9] SR:29 DR:2 LR:-90.67 LO:90.67);ALT=C[chr4:140213681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140211246	+	chr4	140216197	+	TACATTAGTGTTTCAAAAGTTTATTCCAGCCCATTTCTTCTTTTGTACTCTAAAATATCTTCATTGTGTTGTTTGATGAG	0	60	2235528_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TAC;INSERTION=TACATTAGTGTTTCAAAAGTTTATTCCAGCCCATTTCTTCTTTTGTACTCTAAAATATCTTCATTGTGTTGTTTGATGAG;MAPQ=60;MATEID=2235528_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_140213501_140238501_347C;SPAN=4951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:52 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:60 DR:0 LR:-178.2 LO:178.2);ALT=C[chr4:140216197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140213812	+	chr4	140216899	+	.	22	0	2235532_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2235532_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:140213812(+)-4:140216899(-)__4_140213501_140238501D;SPAN=3087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:130 GQ:37.4 PL:[37.4, 0.0, 278.3] SR:0 DR:22 LR:-37.4 LO:48.08);ALT=C[chr4:140216899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140468205	+	chr4	140477251	+	.	7	4	2236333_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2236333_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_4_140458501_140483501_23C;SPAN=9046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:116 GQ:1.5 PL:[0.0, 1.5, 283.8] SR:4 DR:7 LR:1.718 LO:16.41);ALT=T[chr4:140477251[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140587233	+	chr4	140599697	+	.	35	49	2236749_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=2236749_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_140581001_140606001_221C;SPAN=12464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:131 GQ:99 PL:[189.2, 0.0, 126.5] SR:49 DR:35 LR:-189.6 LO:189.6);ALT=T[chr4:140599697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140587250	+	chr4	140616350	+	.	8	0	2237056_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2237056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:140587250(+)-4:140616350(-)__4_140605501_140630501D;SPAN=29100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=T[chr4:140616350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140599796	+	chr4	140616351	+	.	2	24	2237057_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2237057_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_140605501_140630501_12C;SPAN=16555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:53 GQ:58.4 PL:[68.3, 0.0, 58.4] SR:24 DR:2 LR:-68.19 LO:68.19);ALT=A[chr4:140616351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	140616421	+	chr4	140624607	+	.	2	17	2237103_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2237103_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_140605501_140630501_280C;SPAN=8186;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:124 GQ:26 PL:[26.0, 0.0, 273.5] SR:17 DR:2 LR:-25.82 LO:38.02);ALT=G[chr4:140624607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	141294871	+	chr4	141300273	+	.	4	3	2239222_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2239222_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_4_141291501_141316501_21C;SPAN=5402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:115 GQ:17.7 PL:[0.0, 17.7, 313.5] SR:3 DR:4 LR:17.95 LO:5.87);ALT=G[chr4:141300273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	141294903	+	chr4	141300721	+	.	8	0	2239224_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2239224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:141294903(+)-4:141300721(-)__4_141291501_141316501D;SPAN=5818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=G[chr4:141300721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	142230783	+	chr4	142233063	+	.	112	70	2241959_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGCC;MAPQ=60;MATEID=2241959_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_142222501_142247501_77C;SPAN=2280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:38 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:70 DR:112 LR:-445.6 LO:445.6);ALT=C[chr4:142233063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	144894147	+	chr4	144773023	+	.	17	0	2250041_1	48.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=2250041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:144773023(-)-4:144894147(+)__4_144893001_144918001D;SPAN=121124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:27 GQ:15.8 PL:[48.8, 0.0, 15.8] SR:0 DR:17 LR:-49.67 LO:49.67);ALT=]chr4:144894147]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	144905468	+	chr4	145008810	+	.	8	0	2250095_1	16.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2250095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:144905468(+)-4:145008810(-)__4_144893001_144918001D;SPAN=103342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:0 DR:8 LR:-16.65 LO:18.55);ALT=G[chr4:145008810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	145316447	+	chr4	145319906	+	.	19	23	2251772_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=0;MATEID=2251772_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_4_145309501_145334501_424C;SECONDARY;SPAN=3459;SUBN=10;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:63 GQ:35.9 PL:[115.1, 0.0, 35.9] SR:23 DR:19 LR:-117.1 LO:117.1);ALT=C[chr4:145319906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	146019571	+	chr4	146025536	+	.	10	4	2253507_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2253507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_145995501_146020501_385C;SPAN=5965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:4 DR:10 LR:-22.81 LO:27.0);ALT=G[chr4:146025536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	146438813	+	chr4	146440451	+	.	0	42	2254758_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TTGGCCA;MAPQ=60;MATEID=2254758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_146436501_146461501_76C;SPAN=1638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:76 GQ:65.3 PL:[118.1, 0.0, 65.3] SR:42 DR:0 LR:-118.8 LO:118.8);ALT=A[chr4:146440451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	146620415	+	chr10	53798921	-	.	2	16	2256007_1	52.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=TTGCTCACACAAAGCCTGTTTGGTGGTCTCTTCACACGGA;MAPQ=60;MATEID=2256007_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_146608001_146633001_421C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:10 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:16 DR:2 LR:-52.81 LO:52.81);ALT=A]chr10:53798921];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr4	146621100	+	chr7	83089943	+	.	19	61	2256013_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GCTTTTCTGGGGGAGGGGCAAGCACCCC;MAPQ=60;MATEID=2256013_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_146608001_146633001_352C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:64 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:61 DR:19 LR:-234.4 LO:234.4);ALT=C[chr7:83089943[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr4	146919581	+	chr4	146927741	+	.	46	28	2256404_1	99.0	.	DISC_MAPQ=14;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=0;MATEID=2256404_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TT;SCTG=c_4_146926501_146951501_360C;SECONDARY;SPAN=8160;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:36 GQ:18 PL:[198.0, 18.0, 0.0] SR:28 DR:46 LR:-198.0 LO:198.0);ALT=T[chr4:146927741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147096964	+	chr4	147104062	+	.	14	5	2256918_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2256918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_147098001_147123001_83C;SPAN=7098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:50 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:5 DR:14 LR:-39.27 LO:40.1);ALT=G[chr4:147104062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147097007	+	chr4	147108422	+	.	22	0	2256920_1	56.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2256920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:147097007(+)-4:147108422(-)__4_147098001_147123001D;SPAN=11415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:60 GQ:56.3 PL:[56.3, 0.0, 89.3] SR:0 DR:22 LR:-56.37 LO:56.77);ALT=G[chr4:147108422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147104168	+	chr4	147110773	+	GGTCCTGGCTTGCCTGGATGGCTACATGAATATAGCCCTGGAGCAGACAGAAGAATATGTAAATGGACAACTGAAGAATAAGTATGGGGATGCATTTATCCGAGGAAACAAT	0	37	2256935_1	95.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GGTCCTGGCTTGCCTGGATGGCTACATGAATATAGCCCTGGAGCAGACAGAAGAATATGTAAATGGACAACTGAAGAATAAGTATGGGGATGCATTTATCCGAGGAAACAAT;MAPQ=60;MATEID=2256935_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_147098001_147123001_217C;SPAN=6605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:101 GQ:95 PL:[95.0, 0.0, 147.8] SR:37 DR:0 LR:-94.77 LO:95.46);ALT=G[chr4:147110773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147108539	+	chr4	147110773	+	.	0	18	2256957_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2256957_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_4_147098001_147123001_217C;SPAN=2234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:112 GQ:29.3 PL:[29.3, 0.0, 240.5] SR:18 DR:0 LR:-29.07 LO:38.89);ALT=G[chr4:147110773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	147208406	+	chr4	147206794	+	.	91	0	2257297_1	99.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=2257297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:147206794(-)-4:147208406(+)__4_147196001_147221001D;SPAN=1612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:101 GQ:27 PL:[297.0, 27.0, 0.0] SR:0 DR:91 LR:-297.1 LO:297.1);ALT=]chr4:147208406]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr4	154579691	-	chrX	48937461	+	.	13	0	7419059_1	36.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=7419059_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:154579691(-)-23:48937461(-)__23_48926501_48951501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:23 GQ:17 PL:[36.8, 0.0, 17.0] SR:0 DR:13 LR:-36.98 LO:36.98);ALT=[chrX:48937461[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	155078010	+	chr4	155133914	+	.	9	0	2283447_1	26.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2283447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:155078010(+)-4:155133914(-)__4_155134001_155159001D;SPAN=55904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:7 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=T[chr4:155133914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	155469036	+	chr4	155471466	+	.	11	0	2284219_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2284219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:155469036(+)-4:155471466(-)__4_155452501_155477501D;SPAN=2430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:98 GQ:9.8 PL:[9.8, 0.0, 227.6] SR:0 DR:11 LR:-9.76 LO:21.91);ALT=T[chr4:155471466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	157768893	-	chr6	155707847	+	.	16	0	2291158_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2291158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:157768893(-)-6:155707847(-)__4_157755501_157780501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:40 GQ:41.9 PL:[41.9, 0.0, 55.1] SR:0 DR:16 LR:-41.98 LO:42.08);ALT=[chr6:155707847[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr4	158169733	+	chr15	65008157	-	.	7	44	2292398_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATATATA;MAPQ=60;MATEID=2292398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_158147501_158172501_264C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:29 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:44 DR:7 LR:-145.2 LO:145.2);ALT=A]chr15:65008157];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	218547	+	chr5	224474	+	.	20	0	2398023_1	57.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2398023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:218547(+)-5:224474(-)__5_220501_245501D;SPAN=5927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:33 GQ:20.9 PL:[57.2, 0.0, 20.9] SR:0 DR:20 LR:-57.87 LO:57.87);ALT=G[chr5:224474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	271876	+	chr5	306716	+	.	8	0	2398158_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2398158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:271876(+)-5:306716(-)__5_294001_319001D;SPAN=34840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:33 GQ:17.6 PL:[17.6, 0.0, 60.5] SR:0 DR:8 LR:-17.47 LO:18.9);ALT=C[chr5:306716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	306876	+	chr5	311407	+	.	2	3	2398179_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=2398179_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_5_294001_319001_307C;SPAN=4531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:45 GQ:4.4 PL:[4.4, 0.0, 103.4] SR:3 DR:2 LR:-4.313 LO:9.938);ALT=G[chr5:311407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	795415	+	chr5	710186	+	.	12	0	2399335_1	34.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2399335_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:710186(-)-5:795415(+)__5_686001_711001D;SPAN=85229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:21 GQ:14.3 PL:[34.1, 0.0, 14.3] SR:0 DR:12 LR:-34.22 LO:34.22);ALT=]chr5:795415]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1043012	+	chr5	1041007	+	.	50	0	2400174_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2400174_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:1041007(-)-5:1043012(+)__5_1029001_1054001D;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:42 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=]chr5:1043012]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	1094364	+	chr5	1111982	+	.	0	9	2399910_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=2399910_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_1078001_1103001_131C;SPAN=17618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:20 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:9 DR:0 LR:-24.29 LO:24.29);ALT=C[chr5:1111982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	1178294	+	chr5	1180733	+	.	51	30	2400027_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=2400027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_1176001_1201001_111C;SPAN=2439;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:15 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:30 DR:51 LR:-211.3 LO:211.3);ALT=T[chr5:1180733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	1801690	+	chr5	1814450	+	.	84	0	2401318_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2401318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:1801690(+)-5:1814450(-)__5_1813001_1838001D;SPAN=12760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:67 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=C[chr5:1814450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	1814576	+	chr5	1815964	+	.	0	117	2401323_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=2401323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_1813001_1838001_207C;SPAN=1388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:117 DP:156 GQ:33.8 PL:[344.0, 0.0, 33.8] SR:117 DR:0 LR:-358.7 LO:358.7);ALT=G[chr5:1815964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	8749528	+	chr20	23697169	+	.	0	25	2411798_1	72.0	.	EVDNC=ASSMB;HOMSEQ=TAATG;MAPQ=60;MATEID=2411798_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_8746501_8771501_98C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:18 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:25 DR:0 LR:-72.62 LO:72.62);ALT=G[chr20:23697169[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	22863403	+	chr5	9024533	+	.	10	0	6959400_1	27.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=6959400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:9024533(-)-20:22863403(+)__20_22858501_22883501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:19 GQ:17.9 PL:[27.8, 0.0, 17.9] SR:0 DR:10 LR:-27.97 LO:27.97);ALT=]chr20:22863403]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	16451895	+	chr5	16453121	+	.	0	6	2422436_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2422436_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_16439501_16464501_103C;SPAN=1226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:53 GQ:5.6 PL:[5.6, 0.0, 121.1] SR:6 DR:0 LR:-5.447 LO:11.98);ALT=T[chr5:16453121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	17024220	-	chr7	101571683	+	.	14	20	2423795_1	99.0	.	DISC_MAPQ=41;EVDNC=TSI_L;HOMSEQ=CGCCACTGCACTCCAGCCTAGGTGACAGAG;MAPQ=60;MATEID=2423795_2;MATENM=3;NM=0;NUMPARTS=3;SCTG=c_5_17003001_17028001_279C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:28 GQ:9 PL:[99.0, 9.0, 0.0] SR:20 DR:14 LR:-99.02 LO:99.02);ALT=[chr7:101571683[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	32420211	+	chr5	32444335	+	.	0	9	2446606_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CTA;MAPQ=60;MATEID=2446606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32438001_32463001_86C;SPAN=24124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:9 DR:0 LR:-23.75 LO:23.78);ALT=A[chr5:32444335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32420229	+	chr5	32444730	+	.	11	0	2446607_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2446607_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:32420229(+)-5:32444730(-)__5_32438001_32463001D;SPAN=24501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:18 GQ:11.6 PL:[31.4, 0.0, 11.6] SR:0 DR:11 LR:-31.89 LO:31.89);ALT=A[chr5:32444730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32585763	+	chr5	32599063	+	.	15	0	2446916_1	30.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2446916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:32585763(+)-5:32599063(-)__5_32585001_32610001D;SPAN=13300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:69 GQ:30.8 PL:[30.8, 0.0, 136.4] SR:0 DR:15 LR:-30.82 LO:34.61);ALT=T[chr5:32599063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32585763	+	chr5	32591666	+	.	79	0	2446915_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2446915_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:32585763(+)-5:32591666(-)__5_32585001_32610001D;SPAN=5903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:70 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=T[chr5:32591666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32591794	+	chr5	32601109	+	.	2	5	2446927_1	0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=2446927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32585001_32610001_266C;SPAN=9315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:90 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:5 DR:2 LR:1.276 LO:12.77);ALT=A[chr5:32601109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32712651	+	chr5	32724802	+	.	7	5	2447100_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2447100_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32707501_32732501_276C;SPAN=12151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:5 DR:7 LR:-8.577 LO:18.05);ALT=G[chr5:32724802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	32774951	+	chr5	32780826	+	.	2	6	2447269_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2447269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_32756501_32781501_105C;SPAN=5875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:50 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:6 DR:2 LR:-9.561 LO:14.67);ALT=T[chr5:32780826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32655777	+	chr5	33234469	+	.	12	0	2778434_1	33.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=2778434_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:33234469(-)-6:32655777(+)__6_32634001_32659001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:23 GQ:20.3 PL:[33.5, 0.0, 20.3] SR:0 DR:12 LR:-33.5 LO:33.5);ALT=]chr6:32655777]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	33441223	+	chr5	33448644	+	.	11	0	2448094_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2448094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:33441223(+)-5:33448644(-)__5_33442501_33467501D;SPAN=7421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:31 GQ:28.1 PL:[28.1, 0.0, 44.6] SR:0 DR:11 LR:-27.91 LO:28.19);ALT=G[chr5:33448644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	33441249	+	chr5	33445429	+	.	9	11	2448095_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2448095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_33442501_33467501_228C;SPAN=4180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:29 GQ:28.4 PL:[41.6, 0.0, 28.4] SR:11 DR:9 LR:-41.78 LO:41.78);ALT=G[chr5:33445429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	33445510	+	chr5	33448645	+	.	0	11	2448106_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2448106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_33442501_33467501_3C;SPAN=3135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:11 DR:0 LR:-21.14 LO:24.83);ALT=G[chr5:33448645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	33453519	+	chr5	33455050	+	.	2	3	2448117_1	2.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=2448117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_33442501_33467501_242C;SPAN=1531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:51 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:3 DR:2 LR:-2.688 LO:9.65);ALT=T[chr5:33455050[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	105505772	+	chr5	34776912	+	.	2	22	5632322_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAA;MAPQ=60;MATEID=5632322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_105497001_105522001_148C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:36 GQ:23.3 PL:[62.9, 0.0, 23.3] SR:22 DR:2 LR:-63.79 LO:63.79);ALT=]chr13:105505772]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	34916003	+	chr5	34918467	+	.	0	12	2450441_1	26.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2450441_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_34912501_34937501_182C;SPAN=2464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:48 GQ:26.6 PL:[26.6, 0.0, 89.3] SR:12 DR:0 LR:-26.61 LO:28.53);ALT=G[chr5:34918467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	39134489	+	chr5	39137701	+	.	9	0	2457321_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2457321_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:39134489(+)-5:39137701(-)__5_39126501_39151501D;SPAN=3212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=A[chr5:39137701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	39135135	+	chr5	39137701	+	.	16	0	2457323_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2457323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:39135135(+)-5:39137701(-)__5_39126501_39151501D;SPAN=2566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:0 DR:16 LR:-39.54 LO:40.27);ALT=A[chr5:39137701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	39203091	+	chr5	39219544	+	.	24	4	2457365_1	74.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2457365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_39200001_39225001_159C;SPAN=16453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:44 GQ:31.1 PL:[74.0, 0.0, 31.1] SR:4 DR:24 LR:-74.76 LO:74.76);ALT=T[chr5:39219544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	39203138	+	chr5	39270669	+	.	25	0	2457494_1	72.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2457494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:39203138(+)-5:39270669(-)__5_39249001_39274001D;SPAN=67531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:23 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:0 DR:25 LR:-72.62 LO:72.62);ALT=G[chr5:39270669[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	40777746	+	chr5	40798201	+	.	12	0	2459696_1	30.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2459696_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:40777746(+)-5:40798201(-)__5_40792501_40817501D;SPAN=20455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:0 DR:12 LR:-30.67 LO:30.91);ALT=C[chr5:40798201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	41861507	+	chr5	41862742	+	.	0	8	2461050_1	12.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=2461050_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_41846001_41871001_138C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.59 LO:17.19);ALT=C[chr5:41862742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	41904569	+	chr5	41907837	+	.	11	2	2461018_1	19.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2461018_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_41895001_41920001_219C;SPAN=3268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:2 DR:11 LR:-19.51 LO:24.29);ALT=G[chr5:41907837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	41907945	+	chr5	41909846	+	.	0	7	2461024_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2461024_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_41895001_41920001_120C;SPAN=1901;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:48 GQ:10.1 PL:[10.1, 0.0, 105.8] SR:7 DR:0 LR:-10.1 LO:14.8);ALT=G[chr5:41909846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	41925600	+	chr5	41927114	+	.	8	7	2460992_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2460992_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_41919501_41944501_179C;SPAN=1514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:48 GQ:26.6 PL:[26.6, 0.0, 89.3] SR:7 DR:8 LR:-26.61 LO:28.53);ALT=G[chr5:41927114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	42801434	+	chr5	42804758	+	.	5	2	2462320_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2462320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_42801501_42826501_33C;SPAN=3324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:29 GQ:11.9 PL:[11.9, 0.0, 58.1] SR:2 DR:5 LR:-11.95 LO:13.7);ALT=C[chr5:42804758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	42807210	+	chr5	42808253	+	.	0	15	2462327_1	33.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2462327_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_42801501_42826501_228C;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:59 GQ:33.5 PL:[33.5, 0.0, 109.4] SR:15 DR:0 LR:-33.53 LO:35.79);ALT=T[chr5:42808253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	42808493	+	chr5	42811936	+	.	15	0	2462330_1	35.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2462330_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:42808493(+)-5:42811936(-)__5_42801501_42826501D;SPAN=3443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:0 DR:15 LR:-35.16 LO:36.62);ALT=C[chr5:42811936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	43086350	-	chr7	80543734	+	.	29	0	3418480_1	83.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=3418480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:43086350(-)-7:80543734(-)__7_80531501_80556501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:47 GQ:30.2 PL:[83.0, 0.0, 30.2] SR:0 DR:29 LR:-84.29 LO:84.29);ALT=[chr7:80543734[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	43299078	+	chr5	43313458	+	.	10	4	2463130_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2463130_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_43291501_43316501_207C;SPAN=14380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:64 GQ:22.4 PL:[22.4, 0.0, 131.3] SR:4 DR:10 LR:-22.27 LO:26.82);ALT=C[chr5:43313458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	43700339	+	chr5	43702721	+	.	3	4	2463754_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2463754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_43683501_43708501_84C;SPAN=2382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:67 GQ:1.5 PL:[0.0, 1.5, 165.0] SR:4 DR:3 LR:1.647 LO:9.03);ALT=G[chr5:43702721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	54603976	+	chr5	54618154	+	.	12	4	2474426_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2474426_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_54586001_54611001_243C;SPAN=14178;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:23 GQ:17 PL:[36.8, 0.0, 17.0] SR:4 DR:12 LR:-36.98 LO:36.98);ALT=G[chr5:54618154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	58988184	-	chr7	80802156	+	.	13	0	3419191_1	28.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=3419191_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:58988184(-)-7:80802156(-)__7_80801001_80826001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:0 DR:13 LR:-28.55 LO:30.78);ALT=[chr7:80802156[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	64065017	+	chr5	64070516	+	.	3	7	2487555_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2487555_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_64043001_64068001_212C;SPAN=5499;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:22 GQ:20.6 PL:[20.6, 0.0, 30.5] SR:7 DR:3 LR:-20.45 LO:20.61);ALT=T[chr5:64070516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	64070614	+	chr5	64077746	+	.	0	8	2487497_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2487497_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_64067501_64092501_70C;SPAN=7132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.86 LO:17.27);ALT=G[chr5:64077746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	64096154	+	chr5	64100056	+	TGAAAAAGGTGATGCAGCAGATTTAGTTGAT	3	3	2487563_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGAAAAAGGTGATGCAGCAGATTTAGTTGAT;MAPQ=60;MATEID=2487563_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_64092001_64117001_138C;SPAN=3902;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:45 GQ:7.7 PL:[7.7, 0.0, 100.1] SR:3 DR:3 LR:-7.614 LO:12.43);ALT=G[chr5:64100056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	64850817	+	chr5	64858922	+	.	12	0	2488780_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2488780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:64850817(+)-5:64858922(-)__5_64851501_64876501D;SPAN=8105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:28 GQ:32 PL:[32.0, 0.0, 35.3] SR:0 DR:12 LR:-32.03 LO:32.04);ALT=A[chr5:64858922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	65028099	+	chr5	65030381	+	.	0	26	2488972_1	75.0	.	EVDNC=ASSMB;HOMSEQ=AGAAAGACTCTGCCCA;MAPQ=60;MATEID=2488972_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_5_65023001_65048001_101C;SPAN=2282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:17 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:26 DR:0 LR:-75.92 LO:75.92);ALT=A[chr5:65030381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	65222634	+	chr5	65284461	+	.	2	5	2489427_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2489427_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_65268001_65293001_229C;SPAN=61827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:32 GQ:8 PL:[8.0, 0.0, 67.4] SR:5 DR:2 LR:-7.835 LO:10.74);ALT=G[chr5:65284461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	65440365	+	chr5	65449291	+	.	0	11	2489640_1	19.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2489640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_65439501_65464501_65C;SPAN=8926;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:11 DR:0 LR:-19.24 LO:24.2);ALT=A[chr5:65449291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	74063202	+	chr5	74064758	+	.	18	0	2504480_1	59.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2504480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:74063202(+)-5:74064758(-)__5_74063501_74088501D;SPAN=1556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:21 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:18 LR:-57.84 LO:57.84);ALT=C[chr5:74064758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	74066653	+	chr5	74069691	+	.	10	0	2504484_1	19.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2504484_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:74066653(+)-5:74069691(-)__5_74063501_74088501D;SPAN=3038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:0 DR:10 LR:-19.73 LO:22.76);ALT=T[chr5:74069691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	75046591	+	chr12	115330202	+	.	2	37	2505826_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATCTATCTATCTATCTATCTA;MAPQ=60;MATEID=2505826_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_75043501_75068501_245C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:25 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:37 DR:2 LR:-112.2 LO:112.2);ALT=A[chr12:115330202[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr19	33072234	+	chr5	75576783	+	.	27	24	6790035_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=11;MATEID=6790035_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_33050501_33075501_85C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:31 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:24 DR:27 LR:-102.3 LO:102.3);ALT=]chr19:33072234]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	34725363	+	chr5	75672508	+	.	11	0	2789368_1	22.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=2789368_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:75672508(-)-6:34725363(+)__6_34716501_34741501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:0 DR:11 LR:-22.49 LO:25.34);ALT=]chr6:34725363]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	75672575	+	chr6	34738067	+	.	8	0	2789369_1	8.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2789369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:75672575(+)-6:34738067(-)__6_34716501_34741501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=A[chr6:34738067[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	75672583	+	chr6	34735684	+	.	13	0	2789370_1	28.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=2789370_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:75672583(+)-6:34735684(-)__6_34716501_34741501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:54 GQ:28.4 PL:[28.4, 0.0, 101.0] SR:0 DR:13 LR:-28.28 LO:30.66);ALT=G[chr6:34735684[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	75699416	+	chr5	75757395	+	.	2	6	2506732_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2506732_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_75680501_75705501_25C;SPAN=57979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:6 DR:2 LR:-19.91 LO:20.23);ALT=T[chr5:75757395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	75858377	+	chr5	75866403	+	.	3	7	2507109_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2507109_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_75852001_75877001_277C;SPAN=8026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:7 DR:3 LR:-16.48 LO:21.7);ALT=G[chr5:75866403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	75886411	+	chr5	75888661	+	.	2	3	2507159_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2507159_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_5_75876501_75901501_170C;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:49 GQ:0 PL:[0.0, 0.0, 118.8] SR:3 DR:2 LR:0.0713 LO:7.387);ALT=G[chr5:75888661[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76145980	+	chr5	76166020	+	.	63	6	2507680_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2507680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_76146001_76171001_250C;SPAN=20040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:60 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:6 DR:63 LR:-194.7 LO:194.7);ALT=G[chr5:76166020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76146022	+	chr5	76171125	+	.	50	0	2507682_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2507682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:76146022(+)-5:76171125(-)__5_76146001_76171001D;SPAN=25103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:20 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=A[chr5:76171125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76166109	+	chr5	76171127	+	.	2	68	2507723_1	99.0	.	DISC_MAPQ=37;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2507723_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_5_76146001_76171001_91C;SPAN=5018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:43 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:68 DR:2 LR:-204.7 LO:204.7);ALT=G[chr5:76171127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76171325	+	chr5	76173498	+	.	0	19	2507581_1	45.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2507581_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_5_76170501_76195501_258C;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:63 GQ:45.8 PL:[45.8, 0.0, 105.2] SR:19 DR:0 LR:-45.65 LO:47.02);ALT=G[chr5:76173498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76173674	+	chr5	76216538	+	.	10	0	2507631_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2507631_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:76173674(+)-5:76216538(-)__5_76195001_76220001D;SPAN=42864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:30 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:0 DR:10 LR:-24.88 LO:25.28);ALT=C[chr5:76216538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76760685	+	chr5	76787994	+	.	9	0	2508741_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2508741_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:76760685(+)-5:76787994(-)__5_76758501_76783501D;SPAN=27309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:25 GQ:23 PL:[23.0, 0.0, 36.2] SR:0 DR:9 LR:-22.94 LO:23.13);ALT=T[chr5:76787994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	76785399	+	chr5	76787995	+	.	9	3	2508492_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2508492_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_5_76783001_76808001_168C;SPAN=2596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:3 DR:9 LR:-19.51 LO:24.29);ALT=T[chr5:76787995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	77004178	+	chr5	77072040	+	.	22	0	2508890_1	62.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=2508890_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:77004178(+)-5:77072040(-)__5_77052501_77077501D;SPAN=67862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:36 GQ:23.3 PL:[62.9, 0.0, 23.3] SR:0 DR:22 LR:-63.79 LO:63.79);ALT=A[chr5:77072040[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	77081450	-	chr7	5567946	+	.	19	0	3147659_1	8.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=3147659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:77081450(-)-7:5567946(-)__7_5561501_5586501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:201 GQ:8.5 PL:[8.5, 0.0, 477.2] SR:0 DR:19 LR:-8.263 LO:36.35);ALT=[chr7:5567946[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	77081571	+	chr7	5567782	-	.	9	0	3147661_1	0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=3147661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:77081571(+)-7:5567782(+)__7_5561501_5586501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:150 GQ:10.9 PL:[0.0, 10.9, 386.1] SR:0 DR:9 LR:10.93 LO:15.37);ALT=T]chr7:5567782];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	77409748	+	chr5	77411950	+	.	0	7	2509535_1	6.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2509535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_77395501_77420501_249C;SPAN=2202;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:61 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:7 DR:0 LR:-6.581 LO:14.02);ALT=C[chr5:77411950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	77656553	+	chr5	77684659	+	.	11	10	2509925_1	40.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=2509925_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_5_77640501_77665501_222C;SPAN=28106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:22 GQ:10.7 PL:[40.4, 0.0, 10.7] SR:10 DR:11 LR:-41.01 LO:41.01);ALT=G[chr5:77684659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	77656553	+	chr5	77711344	+	ATCCATCAGTTACACAAGTGACAAGAAATGTTCCACCAGGACTTGATGAATATAATCCATTCTCGGATTCTAGAACA	3	17	2509926_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATCCATCAGTTACACAAGTGACAAGAAATGTTCCACCAGGACTTGATGAATATAATCCATTCTCGGATTCTAGAACA;MAPQ=60;MATEID=2509926_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_77640501_77665501_222C;SPAN=54791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:22 GQ:2.4 PL:[56.1, 2.4, 0.0] SR:17 DR:3 LR:-56.8 LO:56.8);ALT=G[chr5:77711344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	80064822	+	chr5	80071511	+	.	2	3	2513966_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2513966_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_5_80066001_80091001_160C;SPAN=6689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:25 GQ:6.5 PL:[6.5, 0.0, 52.7] SR:3 DR:2 LR:-6.431 LO:8.634);ALT=G[chr5:80071511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	80809536	+	chr5	81046798	+	GTAATCATGGAAGGCTTTTGCTTCACTTGAGTGTTCACATGTTTCACGTCTCTCTGGAGCTGCACAGTAGAGATCCCAAAATACACACCACCAAGAATGTAAGAATCCTGGTGGTTCCCCCAATGTGATGTTTTTTTCCCATCTTATCTCTGATAAAAATGTTTGAGCTGATTTCTGAGCTCCTACATGGAGCAGATATTCATATACGTAGAGTGCTA	3	20	2515396_1	69.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=GTAATCATGGAAGGCTTTTGCTTCACTTGAGTGTTCACATGTTTCACGTCTCTCTGGAGCTGCACAGTAGAGATCCCAAAATACACACCACCAAGAATGTAAGAATCCTGGTGGTTCCCCCAATGTGATGTTTTTTTCCCATCTTATCTCTGATAAAAATGTTTGAGCTGATTTCTGAGCTCCTACATGGAGCAGATATTCATATACGTAGAGTGCTA;MAPQ=60;MATEID=2515396_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_5_81046001_81071001_232C;SPAN=237262;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:24 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:20 DR:3 LR:-69.32 LO:69.32);ALT=T[chr5:81046798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	80911425	+	chr5	81046806	+	.	25	0	2515658_1	72.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2515658_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:80911425(+)-5:81046806(-)__5_80899001_80924001D;SPAN=135381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:18 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:0 DR:25 LR:-72.62 LO:72.62);ALT=T[chr5:81046806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	80932482	+	chr5	81046807	+	.	19	0	2515448_1	59.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2515448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:80932482(+)-5:81046807(-)__5_80923501_80948501D;SPAN=114325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:23 GQ:2.7 PL:[59.4, 2.7, 0.0] SR:0 DR:19 LR:-60.16 LO:60.16);ALT=T[chr5:81046807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	80946158	+	chr5	81046798	+	.	10	4	2515465_1	30.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AC;MAPQ=60;MATEID=2515465_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TCTC;SCTG=c_5_80923501_80948501_203C;SPAN=100640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:23 GQ:23.6 PL:[30.2, 0.0, 23.6] SR:4 DR:10 LR:-30.1 LO:30.1);ALT=C[chr5:81046798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	81572337	+	chr5	81573523	+	.	10	0	2516214_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=2516214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:81572337(+)-5:81573523(-)__5_81560501_81585501D;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:470 GQ:94.2 PL:[0.0, 94.2, 1330.0] SR:0 DR:10 LR:94.33 LO:12.54);ALT=T[chr5:81573523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	81572339	+	chr5	81574137	+	.	60	0	2516215_1	0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2516215_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:81572339(+)-5:81574137(-)__5_81560501_81585501D;SPAN=1798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:60 DP:1079 GQ:94 PL:[0.0, 94.0, 2809.0] SR:0 DR:60 LR:94.27 LO:100.5);ALT=T[chr5:81574137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	82352973	+	chr5	82373139	+	.	21	0	2517269_1	56.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2517269_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:82352973(+)-5:82373139(-)__5_82369001_82394001D;SPAN=20166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:49 GQ:56 PL:[56.0, 0.0, 62.6] SR:0 DR:21 LR:-56.05 LO:56.07);ALT=C[chr5:82373139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	82352974	+	chr5	82360827	+	AATTCTGGCACACTTCCAAAATATACCCAACAAT	0	24	2517150_1	63.0	.	EVDNC=ASSMB;INSERTION=AATTCTGGCACACTTCCAAAATATACCCAACAAT;MAPQ=60;MATEID=2517150_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_82344501_82369501_154C;SPAN=7853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:57 GQ:63.8 PL:[63.8, 0.0, 73.7] SR:24 DR:0 LR:-63.78 LO:63.83);ALT=C[chr5:82360827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	82373139	-	chr19	14903115	+	.	11	0	6743518_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6743518_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:82373139(-)-19:14903115(-)__19_14896001_14921001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=[chr19:14903115[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	82789752	+	chr5	82807921	+	.	6	3	2517690_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2517690_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_82785501_82810501_177C;SPAN=18169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:3 DR:6 LR:-9.832 LO:14.73);ALT=T[chr5:82807921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64289967	+	chr5	92975971	+	.	8	0	3344752_1	18.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=3344752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:92975971(-)-7:64289967(+)__7_64288001_64313001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:29 GQ:18.5 PL:[18.5, 0.0, 51.5] SR:0 DR:8 LR:-18.55 LO:19.42);ALT=]chr7:64289967]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	93386536	+	chr5	93388831	+	.	0	7	2530972_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2530972_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_93369501_93394501_134C;SPAN=2295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:43 GQ:11.6 PL:[11.6, 0.0, 90.8] SR:7 DR:0 LR:-11.46 LO:15.17);ALT=T[chr5:93388831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	94275903	+	chr5	94278051	+	.	0	8	2532041_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CCTGT;MAPQ=60;MATEID=2532041_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_94276001_94301001_5C;SPAN=2148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:30 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:8 DR:0 LR:-18.28 LO:19.28);ALT=T[chr5:94278051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	94353190	+	chr5	94417130	+	.	27	24	2532200_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2532200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_94398501_94423501_6C;SPAN=63940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:45 GQ:5.4 PL:[118.8, 5.4, 0.0] SR:24 DR:27 LR:-121.4 LO:121.4);ALT=T[chr5:94417130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	94415670	+	chr5	94417129	+	.	0	6	2532241_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2532241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_94398501_94423501_207C;SPAN=1459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:64 GQ:2.6 PL:[2.6, 0.0, 151.1] SR:6 DR:0 LR:-2.467 LO:11.46);ALT=T[chr5:94417129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	95152331	+	chr5	95158157	+	.	0	18	2533185_1	53.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=57;MATEID=2533185_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_95158001_95183001_198C;SPAN=5826;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:23 GQ:0.5 PL:[53.3, 0.0, 0.5] SR:18 DR:0 LR:-55.93 LO:55.93);ALT=C[chr5:95158157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	95998178	+	chr5	96031537	+	.	11	0	2534312_1	27.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2534312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:95998178(+)-5:96031537(-)__5_96015501_96040501D;SPAN=33359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:33 GQ:27.5 PL:[27.5, 0.0, 50.6] SR:0 DR:11 LR:-27.37 LO:27.81);ALT=G[chr5:96031537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	95998201	+	chr5	96011241	+	.	14	26	2534358_1	92.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2534358_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_95991001_96016001_323C;SPAN=13040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:49 GQ:26.3 PL:[92.3, 0.0, 26.3] SR:26 DR:14 LR:-94.38 LO:94.38);ALT=G[chr5:96011241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	96101850	+	chr5	96103609	+	ACAAACCAGTGAAGCCACCTACAAAGAAATCAGAGGATTCAA	3	8	2534480_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACAAACCAGTGAAGCCACCTACAAAGAAATCAGAGGATTCAA;MAPQ=60;MATEID=2534480_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_96089001_96114001_131C;SPAN=1759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:8 DR:3 LR:-14.0 LO:19.3);ALT=G[chr5:96103609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	96106306	+	chr5	96108343	+	ACAACAGAGGAAACTTCCAAGCCAAAAGATGACTAAAGAAATACAAGTTAAGGTATCT	2	10	2534494_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GGTA;INSERTION=ACAACAGAGGAAACTTCCAAGCCAAAAGATGACTAAAGAAATACAAGTTAAGGTATCT;MAPQ=60;MATEID=2534494_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_96089001_96114001_5C;SPAN=2037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:10 DR:2 LR:-27.42 LO:28.93);ALT=G[chr5:96108343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	96139655	+	chr5	96143558	+	.	14	0	2534683_1	31.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2534683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:96139655(+)-5:96143558(-)__5_96138001_96163001D;SPAN=3903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:54 GQ:31.7 PL:[31.7, 0.0, 97.7] SR:0 DR:14 LR:-31.58 LO:33.55);ALT=A[chr5:96143558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	96225009	+	chr5	96228002	+	.	2	4	2534598_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2534598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_96211501_96236501_85C;SPAN=2993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:62 GQ:0 PL:[0.0, 0.0, 148.5] SR:4 DR:2 LR:0.2923 LO:9.206);ALT=G[chr5:96228002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	96271921	+	chr5	96314840	+	.	10	0	2534831_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2534831_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:96271921(+)-5:96314840(-)__5_96309501_96334501D;SPAN=42919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:29 GQ:25.1 PL:[25.1, 0.0, 44.9] SR:0 DR:10 LR:-25.15 LO:25.47);ALT=C[chr5:96314840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108120765	-	chr5	180668490	+	.	9	0	2660728_1	19.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=2660728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:108120765(-)-5:180668490(-)__5_180663001_180688001D;SPAN=72547725;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:0 DR:9 LR:-19.41 LO:21.15);ALT=[chr5:180668490[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	108120899	+	chr5	180665239	-	.	17	0	2660730_1	34.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=2660730_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:108120899(+)-5:180665239(+)__5_180663001_180688001D;SPAN=72544340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:79 GQ:34.7 PL:[34.7, 0.0, 156.8] SR:0 DR:17 LR:-34.71 LO:39.14);ALT=A]chr5:180665239];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	108230344	+	chr6	31774531	+	.	85	0	2775157_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=2775157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:108230344(+)-6:31774531(-)__6_31752001_31777001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:77 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:0 DR:85 LR:-250.9 LO:250.9);ALT=T[chr6:31774531[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	108595089	+	chr5	108601122	+	.	63	36	2550904_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAAATAAGAATGG;MAPQ=60;MATEID=2550904_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_108584001_108609001_141C;SPAN=6033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:40 GQ:21 PL:[231.0, 21.0, 0.0] SR:36 DR:63 LR:-231.1 LO:231.1);ALT=G[chr5:108601122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108679075	+	chr10	70973334	-	.	2	10	4622956_1	31.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTT;MAPQ=60;MATEID=4622956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70952001_70977001_260C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:19 GQ:14.6 PL:[31.1, 0.0, 14.6] SR:10 DR:2 LR:-31.47 LO:31.47);ALT=A]chr10:70973334];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr5	108691729	+	chr5	108698541	+	.	3	3	2550678_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2550678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_108682001_108707001_80C;SPAN=6812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:47 GQ:3.8 PL:[3.8, 0.0, 109.4] SR:3 DR:3 LR:-3.772 LO:9.838);ALT=T[chr5:108698541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108714957	+	chr5	108717202	+	.	4	6	2550767_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=2550767_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_108706501_108731501_154C;SPAN=2245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:6 DR:4 LR:-15.35 LO:19.68);ALT=T[chr5:108717202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108717407	+	chr5	108719104	+	.	0	12	2550773_1	25.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=2550773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_108706501_108731501_184C;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:12 DR:0 LR:-25.52 LO:28.05);ALT=G[chr5:108719104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	108719239	+	chr5	108745555	+	.	10	0	2550839_1	26.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2550839_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:108719239(+)-5:108745555(-)__5_108731001_108756001D;SPAN=26316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:0 DR:10 LR:-26.24 LO:26.3);ALT=A[chr5:108745555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	112197123	+	chr18	56835763	+	.	40	0	6640949_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6640949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:112197123(+)-18:56835763(-)__18_56815501_56840501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:40 LR:-130.9 LO:130.9);ALT=T[chr18:56835763[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chrX	15808690	+	chr5	112227382	+	.	10	0	7370943_1	25.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=7370943_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:112227382(-)-23:15808690(+)__23_15802501_15827501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:28 GQ:25.4 PL:[25.4, 0.0, 41.9] SR:0 DR:10 LR:-25.42 LO:25.66);ALT=]chrX:15808690]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	112238215	+	chr5	112256860	+	.	0	8	2555468_1	7.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2555468_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_112234501_112259501_154C;SPAN=18645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:8 DR:0 LR:-7.172 LO:15.95);ALT=T[chr5:112256860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	112312675	+	chr5	112321529	+	CTCTG	8	5	2555603_1	14.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=CTCTG;MAPQ=60;MATEID=2555603_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_112308001_112333001_250C;SPAN=8854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:5 DR:8 LR:-14.59 LO:21.18);ALT=T[chr5:112321529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	112321683	+	chr5	112327818	+	.	0	8	2555612_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2555612_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_112308001_112333001_156C;SPAN=6135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.59 LO:17.19);ALT=G[chr5:112327818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131746735	+	chr5	131755513	+	.	34	11	2582387_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2582387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_131736501_131761501_94C;SPAN=8778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:70 GQ:63.5 PL:[106.4, 0.0, 63.5] SR:11 DR:34 LR:-107.1 LO:107.1);ALT=T[chr5:131755513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131746757	+	chr5	131811356	+	.	10	0	2582547_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2582547_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:131746757(+)-5:131811356(-)__5_131810001_131835001D;SPAN=64599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:20 GQ:20.9 PL:[27.5, 0.0, 20.9] SR:0 DR:10 LR:-27.64 LO:27.64);ALT=G[chr5:131811356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131755635	+	chr5	131811357	+	CCAGAGTTTGTAGCCTATTGGAGGAAAACACACCA	3	23	2582549_1	69.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCAGAGTTTGTAGCCTATTGGAGGAAAACACACCA;MAPQ=60;MATEID=2582549_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_5_131810001_131835001_189C;SPAN=55722;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:20 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:23 DR:3 LR:-69.32 LO:69.32);ALT=G[chr5:131811357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131820191	+	chr5	131821359	+	.	2	4	2582573_1	7.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2582573_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_131810001_131835001_328C;SPAN=1168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:47 GQ:7.1 PL:[7.1, 0.0, 106.1] SR:4 DR:2 LR:-7.073 LO:12.31);ALT=T[chr5:131821359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131823719	+	chr5	131826236	+	.	9	9	2582585_1	31.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2582585_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_131810001_131835001_42C;SPAN=2517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:68 GQ:31.1 PL:[31.1, 0.0, 133.4] SR:9 DR:9 LR:-31.09 LO:34.72);ALT=T[chr5:131826236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	131825177	+	chr5	131826237	+	.	39	48	2582587_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2582587_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TGCTGC;SCTG=c_5_131810001_131835001_214C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:69 GQ:18.5 PL:[161.2, 18.5, 0.0] SR:48 DR:39 LR:-161.3 LO:161.3);ALT=T[chr5:131826237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	132060525	+	chr19	38248879	+	.	2	7	2582970_1	19.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=ATATATATATATATATATATATATATA;MAPQ=20;MATEID=2582970_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_132055001_132080001_226C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:15 GQ:15.8 PL:[19.1, 0.0, 15.8] SR:7 DR:2 LR:-19.05 LO:19.05);ALT=A[chr19:38248879[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	132388082	+	chr5	132403121	+	.	8	0	2583651_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2583651_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:132388082(+)-5:132403121(-)__5_132373501_132398501D;SPAN=15039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:0 DR:8 LR:-16.11 LO:18.33);ALT=G[chr5:132403121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	132400733	+	chr5	132403107	+	.	2	3	2583567_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGTAA;MAPQ=60;MATEID=2583567_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_5_132398001_132423001_68C;SPAN=2374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:51 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:3 DR:2 LR:0.6132 LO:7.314);ALT=A[chr5:132403107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133134710	+	chr5	133136486	+	.	51	0	2584716_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2584716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133134710(+)-5:133136486(-)__5_133133001_133158001D;SPAN=1776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:10 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:51 LR:-148.5 LO:148.5);ALT=A[chr5:133136486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133295744	+	chr5	133304217	+	.	25	0	2584929_1	66.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2584929_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133295744(+)-5:133304217(-)__5_133280001_133305001D;SPAN=8473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:61 GQ:66.2 PL:[66.2, 0.0, 79.4] SR:0 DR:25 LR:-66.0 LO:66.1);ALT=T[chr5:133304217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133326842	+	chr5	133340337	+	.	24	0	2585010_1	69.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=2585010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133326842(+)-5:133340337(-)__5_133329001_133354001D;SPAN=13495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:16 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=A[chr5:133340337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49397979	+	chr5	133340188	+	.	98	0	7419751_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7419751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133340188(-)-23:49397979(+)__23_49392001_49417001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:36 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:0 DR:98 LR:-290.5 LO:290.5);ALT=]chrX:49397979]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	133496836	+	chr5	133512576	+	.	39	0	2585645_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2585645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133496836(+)-5:133512576(-)__5_133500501_133525501D;SPAN=15740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:98 GQ:99 PL:[102.2, 0.0, 135.2] SR:0 DR:39 LR:-102.2 LO:102.4);ALT=G[chr5:133512576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133502964	+	chr5	133512578	+	.	9	0	2585652_1	0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2585652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133502964(+)-5:133512578(-)__5_133500501_133525501D;SPAN=9614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:134 GQ:6.3 PL:[0.0, 6.3, 336.6] SR:0 DR:9 LR:6.595 LO:15.83);ALT=C[chr5:133512578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133509713	+	chr5	133512546	+	.	61	43	2585664_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;MAPQ=20;MATEID=2585664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133500501_133525501_277C;SPAN=2833;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:63 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:43 DR:61 LR:-270.7 LO:270.7);ALT=T[chr5:133512546[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133533535	+	chr5	133534777	+	.	5	5	2585497_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2585497_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133525001_133550001_215C;SPAN=1242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:5 DR:5 LR:-20.55 LO:23.07);ALT=G[chr5:133534777[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133541824	+	chr5	133561450	+	.	2	22	2585525_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2585525_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133525001_133550001_285C;SPAN=19626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:28 GQ:0.9 PL:[69.3, 0.9, 0.0] SR:22 DR:2 LR:-72.68 LO:72.68);ALT=T[chr5:133561450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133541866	+	chr5	133561684	+	.	10	0	2585526_1	26.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2585526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133541866(+)-5:133561684(-)__5_133525001_133550001D;SPAN=19818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:0 DR:10 LR:-26.78 LO:26.78);ALT=A[chr5:133561684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133707332	+	chr5	133710073	+	.	26	20	2585731_1	97.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2585731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133696501_133721501_190C;SPAN=2741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:67 GQ:64.4 PL:[97.4, 0.0, 64.4] SR:20 DR:26 LR:-97.72 LO:97.72);ALT=T[chr5:133710073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133707348	+	chr5	133716408	+	.	8	0	2585733_1	12.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2585733_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133707348(+)-5:133716408(-)__5_133696501_133721501D;SPAN=9060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=C[chr5:133716408[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133710154	+	chr5	133724015	+	ACCAGAAGGGACACCTTTTGAAGATGGTACTTTTAAACTAGTAATAGAATTTTCTGAAGAATATCCAAATAAACCACCAACTGTTAGGTTTTTATCCAAAATGTTTCATCCAAAT	0	21	2585740_1	59.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACCAGAAGGGACACCTTTTGAAGATGGTACTTTTAAACTAGTAATAGAATTTTCTGAAGAATATCCAAATAAACCACCAACTGTTAGGTTTTTATCCAAAATGTTTCATCCAAAT;MAPQ=60;MATEID=2585740_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_133696501_133721501_64C;SPAN=13861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:37 GQ:29.6 PL:[59.3, 0.0, 29.6] SR:21 DR:0 LR:-59.79 LO:59.79);ALT=G[chr5:133724015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133716499	+	chr5	133724015	+	ACCAGAAGGGACACCTTTTGAAGAT	2	6	2585750_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;INSERTION=ACCAGAAGGGACACCTTTTGAAGAT;MAPQ=60;MATEID=2585750_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_133696501_133721501_64C;SPAN=7516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:17 GQ:15.2 PL:[15.2, 0.0, 25.1] SR:6 DR:2 LR:-15.2 LO:15.36);ALT=G[chr5:133724015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133948446	+	chr5	133956623	+	.	0	7	2586439_1	8.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2586439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_133941501_133966501_251C;SPAN=8177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:56 GQ:8 PL:[8.0, 0.0, 126.8] SR:7 DR:0 LR:-7.935 LO:14.3);ALT=G[chr5:133956623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	133956790	+	chr5	133968419	+	.	8	0	2586545_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2586545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:133956790(+)-5:133968419(-)__5_133966001_133991001D;SPAN=11629;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=T[chr5:133968419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134074482	+	chr5	134086448	+	.	12	12	2586641_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2586641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134064001_134089001_260C;SPAN=11966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:81 GQ:41 PL:[41.0, 0.0, 153.2] SR:12 DR:12 LR:-40.77 LO:44.56);ALT=G[chr5:134086448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134074482	+	chr5	134076752	+	.	13	15	2586638_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2586638_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134064001_134089001_117C;SPAN=2270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:82 GQ:47.3 PL:[47.3, 0.0, 149.6] SR:15 DR:13 LR:-47.11 LO:50.19);ALT=G[chr5:134076752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134094645	+	chr5	134102605	+	CCACTATCGAAAACGATCGGCATCCCGGGGTCGCTCTGGAAGTCGGTCTAGAAGTCGCTCACCCTCAGACAAAAGAAGTAAACGTGGAGATGACAGACGGTCTAGAAGTAGAGATAGAGATAGGAGGAGAGAGAGGTCTCGTAGCAGGGATAAAAGAAGATCTCGGTCAAGGGACAGGAAGCGTCTG	0	122	2586728_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCACTATCGAAAACGATCGGCATCCCGGGGTCGCTCTGGAAGTCGGTCTAGAAGTCGCTCACCCTCAGACAAAAGAAGTAAACGTGGAGATGACAGACGGTCTAGAAGTAGAGATAGAGATAGGAGGAGAGAGAGGTCTCGTAGCAGGGATAAAAGAAGATCTCGGTCAAGGGACAGGAAGCGTCTG;MAPQ=60;MATEID=2586728_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_134088501_134113501_116C;SPAN=7960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:92 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:122 DR:0 LR:-359.8 LO:359.8);ALT=G[chr5:134102605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134094645	+	chr5	134099593	+	.	79	53	2586727_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2586727_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_134088501_134113501_116C;SPAN=4948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:86 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:53 DR:79 LR:-307.0 LO:307.0);ALT=G[chr5:134099593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134099782	+	chr5	134102605	+	.	5	68	2586734_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2586734_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_134088501_134113501_116C;SPAN=2823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:91 GQ:5.3 PL:[213.2, 0.0, 5.3] SR:68 DR:5 LR:-224.5 LO:224.5);ALT=G[chr5:134102605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134102750	+	chr5	134109386	+	ATCTAGGTCCAAAGAGAAAACTGATGGTGGGGAAAGTTCTAAAGAGAAGAAAAAAGACAAAGATGACAAGGAGGATGAAAAAGAAAAAGATGCTGGC	4	58	2586741_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TAG;INSERTION=ATCTAGGTCCAAAGAGAAAACTGATGGTGGGGAAAGTTCTAAAGAGAAGAAAAAAGACAAAGATGACAAGGAGGATGAAAAAGAAAAAGATGCTGGC;MAPQ=60;MATEID=2586741_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_134088501_134113501_267C;SPAN=6636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:72 GQ:6 PL:[184.8, 6.0, 0.0] SR:58 DR:4 LR:-190.6 LO:190.6);ALT=G[chr5:134109386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134119203	+	chr9	133575626	+	.	17	0	2586770_1	52.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2586770_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:134119203(+)-9:133575626(-)__5_134113001_134138001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:18 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:17 LR:-52.81 LO:52.81);ALT=A[chr9:133575626[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	134181902	+	chr5	134190586	+	.	11	13	2587010_1	49.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2587010_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134162001_134187001_127C;SPAN=8684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:25 GQ:9.8 PL:[49.4, 0.0, 9.8] SR:13 DR:11 LR:-50.68 LO:50.68);ALT=G[chr5:134190586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134210220	+	chr5	134223384	+	.	7	5	2586915_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2586915_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134211001_134236001_58C;SPAN=13164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:32 GQ:27.8 PL:[27.8, 0.0, 47.6] SR:5 DR:7 LR:-27.64 LO:28.0);ALT=G[chr5:134223384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134670834	+	chr5	134678949	+	.	15	27	2587689_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=2587689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134652001_134677001_11C;SPAN=8115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:46 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:27 DR:15 LR:-134.4 LO:134.4);ALT=G[chr5:134678949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134679126	+	chr5	134681658	+	.	10	9	2587703_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2587703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134676501_134701501_222C;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:61 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:9 DR:10 LR:-42.89 LO:44.34);ALT=T[chr5:134681658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134681749	+	chr5	134696186	+	.	7	3	2587709_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2587709_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134676501_134701501_59C;SPAN=14437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:3 DR:7 LR:-11.24 LO:16.84);ALT=T[chr5:134696186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134681751	+	chr5	134688635	+	.	0	11	2587710_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CCTAG;MAPQ=60;MATEID=2587710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134676501_134701501_152C;SPAN=6884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:64 GQ:19.1 PL:[19.1, 0.0, 134.6] SR:11 DR:0 LR:-18.97 LO:24.12);ALT=G[chr5:134688635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134681788	+	chr5	134705095	+	.	8	0	2587711_1	19.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2587711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:134681788(+)-5:134705095(-)__5_134676501_134701501D;SPAN=23307;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:0 DR:8 LR:-19.36 LO:19.88);ALT=C[chr5:134705095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134688737	+	chr5	134696187	+	.	6	12	2587722_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2587722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134676501_134701501_287C;SPAN=7450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:49 GQ:29.6 PL:[29.6, 0.0, 89.0] SR:12 DR:6 LR:-29.64 LO:31.3);ALT=T[chr5:134696187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134696301	+	chr5	134705096	+	.	5	5	2587734_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTTG;MAPQ=60;MATEID=2587734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134676501_134701501_100C;SPAN=8795;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:5 DR:5 LR:-19.41 LO:21.15);ALT=G[chr5:134705096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134705836	+	chr5	134724612	+	.	3	35	2587640_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGT;MAPQ=60;MATEID=2587640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134701001_134726001_8C;SPAN=18776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:76 GQ:81.8 PL:[101.6, 0.0, 81.8] SR:35 DR:3 LR:-101.6 LO:101.6);ALT=T[chr5:134724612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134705878	+	chr5	134734798	+	.	13	0	2587826_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2587826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:134705878(+)-5:134734798(-)__5_134725501_134750501D;SPAN=28920;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:0 DR:13 LR:-22.32 LO:28.48);ALT=T[chr5:134734798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	134724816	+	chr5	134734752	+	.	135	30	2587827_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=2587827_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_134725501_134750501_2C;SPAN=9936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:165 DP:47 GQ:44.5 PL:[488.5, 44.5, 0.0] SR:30 DR:135 LR:-488.5 LO:488.5);ALT=A[chr5:134734752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	136854719	+	chr5	136856379	+	.	58	0	2590927_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2590927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:136854719(+)-5:136856379(-)__5_136857001_136882001D;SPAN=1660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:0 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=T[chr5:136856379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	137674038	+	chr5	137676887	+	.	8	0	2592154_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2592154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:137674038(+)-5:137676887(-)__5_137665501_137690501D;SPAN=2849;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=G[chr5:137676887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	137854557	+	chr5	137878522	+	.	0	9	2592912_1	23.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2592912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_137837001_137862001_273C;SPAN=23965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:25 GQ:23 PL:[23.0, 0.0, 36.2] SR:9 DR:0 LR:-22.94 LO:23.13);ALT=C[chr5:137878522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	137854603	+	chr5	137878782	+	.	11	0	2592913_1	30.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=2592913_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:137854603(+)-5:137878782(-)__5_137837001_137862001D;SPAN=24179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:22 GQ:20.6 PL:[30.5, 0.0, 20.6] SR:0 DR:11 LR:-30.4 LO:30.4);ALT=T[chr5:137878782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	137909542	+	chr5	137910927	+	.	14	3	2592874_1	33.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2592874_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_137886001_137911001_223C;SPAN=1385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:61 GQ:33.2 PL:[33.2, 0.0, 112.4] SR:3 DR:14 LR:-32.99 LO:35.54);ALT=G[chr5:137910927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	137909817	+	chr5	137910926	+	.	5	9	2592875_1	27.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2592875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_137886001_137911001_318C;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:9 DR:5 LR:-27.52 LO:31.83);ALT=T[chr5:137910926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138089206	+	chr5	138117609	+	.	8	0	2593267_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2593267_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138089206(+)-5:138117609(-)__5_138106501_138131501D;SPAN=28403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=T[chr5:138117609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138356984	+	chr5	138362490	+	.	3	2	2593642_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2593642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138351501_138376501_93C;SPAN=5506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:54 GQ:2 PL:[2.0, 0.0, 127.4] SR:2 DR:3 LR:-1.875 LO:9.519);ALT=G[chr5:138362490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138386737	+	chr5	138456723	+	.	2	7	2593760_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2593760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138376001_138401001_50C;SPAN=69986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:7 DR:2 LR:-17.2 LO:18.78);ALT=T[chr5:138456723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138456863	+	chr5	138463428	+	.	2	8	2593869_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2593869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138449501_138474501_71C;SPAN=6565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:8 DR:2 LR:-11.83 LO:18.75);ALT=C[chr5:138463428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138456906	+	chr5	138533955	+	.	20	0	2594039_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2594039_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138456906(+)-5:138533955(-)__5_138523001_138548001D;SPAN=77049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:30 GQ:14.9 PL:[57.8, 0.0, 14.9] SR:0 DR:20 LR:-59.31 LO:59.31);ALT=C[chr5:138533955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138463544	+	chr5	138533955	+	.	9	0	2594040_1	21.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2594040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138463544(+)-5:138533955(-)__5_138523001_138548001D;SPAN=70411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:30 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.58 LO:22.25);ALT=T[chr5:138533955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138609886	+	chr5	138614737	+	.	15	0	2594116_1	35.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2594116_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138609886(+)-5:138614737(-)__5_138596501_138621501D;SPAN=4851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:52 GQ:35.6 PL:[35.6, 0.0, 88.4] SR:0 DR:15 LR:-35.43 LO:36.77);ALT=T[chr5:138614737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138629758	+	chr5	138642921	+	.	30	0	2594162_1	83.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2594162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138629758(+)-5:138642921(-)__5_138621001_138646001D;SPAN=13163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:56 GQ:50.9 PL:[83.9, 0.0, 50.9] SR:0 DR:30 LR:-84.26 LO:84.26);ALT=C[chr5:138642921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138658697	+	chr5	138661124	+	.	9	0	2594299_1	17.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=2594299_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138658697(+)-5:138661124(-)__5_138645501_138670501D;SPAN=2427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=A[chr5:138661124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138677671	+	chr5	138699447	+	.	99	31	2594459_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2594459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138694501_138719501_118C;SPAN=21776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:42 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:31 DR:99 LR:-343.3 LO:343.3);ALT=T[chr5:138699447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138677675	+	chr5	138700252	+	.	15	0	2594460_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2594460_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138677675(+)-5:138700252(-)__5_138694501_138719501D;SPAN=22577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:32 GQ:34.4 PL:[41.0, 0.0, 34.4] SR:0 DR:15 LR:-40.86 LO:40.86);ALT=G[chr5:138700252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138699611	+	chr5	138704421	+	ATAGAAGAGGAGTTATGGGAAGAAGAATTTATTGAACGCTGTTTCCAAGAAATGCTGGAAGAGGAAGAAGAGCATGAATGGTTTATTCCAGCTCGAGATCTCCCACAAACTATGGACCAAATCCAAGACCAGTTTAATGACCTTGTTATCAGTGATGGCTCTTCTCTGGAAGATCTTGT	0	52	2594474_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=ATAGAAGAGGAGTTATGGGAAGAAGAATTTATTGAACGCTGTTTCCAAGAAATGCTGGAAGAGGAAGAAGAGCATGAATGGTTTATTCCAGCTCGAGATCTCCCACAAACTATGGACCAAATCCAAGACCAGTTTAATGACCTTGTTATCAGTGATGGCTCTTCTCTGGAAGATCTTGT;MAPQ=60;MATEID=2594474_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_138694501_138719501_225C;SPAN=4810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:75 GQ:29.3 PL:[151.4, 0.0, 29.3] SR:52 DR:0 LR:-155.8 LO:155.8);ALT=A[chr5:138704421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138700434	+	chr5	138704421	+	.	11	15	2594476_1	64.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=2594476_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_5_138694501_138719501_225C;SPAN=3987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:67 GQ:64.4 PL:[64.4, 0.0, 97.4] SR:15 DR:11 LR:-64.37 LO:64.76);ALT=T[chr5:138704421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138724385	+	chr5	138725493	+	.	17	0	2594418_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2594418_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138724385(+)-5:138725493(-)__5_138719001_138744001D;SPAN=1108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:66 GQ:38.3 PL:[38.3, 0.0, 120.8] SR:0 DR:17 LR:-38.24 LO:40.68);ALT=G[chr5:138725493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138856040	+	chr5	138857855	+	.	6	4	2594640_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2594640_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_5_138841501_138866501_88C;SPAN=1815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:63 GQ:16.1 PL:[16.1, 0.0, 134.9] SR:4 DR:6 LR:-15.94 LO:21.55);ALT=C[chr5:138857855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138858096	+	chr5	138860375	+	.	6	4	2594646_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2594646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138841501_138866501_81C;SPAN=2279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:4 DR:6 LR:-5.818 LO:15.7);ALT=G[chr5:138860375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138941401	+	chr5	138979955	+	.	18	24	2594976_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=2594976_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_5_138964001_138989001_53C;SPAN=38554;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:24 DR:18 LR:-99.02 LO:99.02);ALT=G[chr5:138979955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138941452	+	chr5	138994281	+	.	25	0	2594911_1	74.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2594911_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:138941452(+)-5:138994281(-)__5_138988501_139013501D;SPAN=52829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:32 GQ:1.4 PL:[74.0, 0.0, 1.4] SR:0 DR:25 LR:-77.64 LO:77.64);ALT=C[chr5:138994281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138980020	+	chr5	138994282	+	TGTTCCATTGGCAAGCTACAATAATGGGGCCA	3	34	2595008_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;INSERTION=TGTTCCATTGGCAAGCTACAATAATGGGGCCA;MAPQ=60;MATEID=2595008_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_138964001_138989001_53C;SPAN=14262;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:30 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:34 DR:3 LR:-102.3 LO:102.3);ALT=A[chr5:138994282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	138994551	+	chr5	139002951	+	.	0	38	2594925_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2594925_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138988501_139013501_98C;SPAN=8400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:62 GQ:39.5 PL:[108.8, 0.0, 39.5] SR:38 DR:0 LR:-110.3 LO:110.3);ALT=G[chr5:139002951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139003049	+	chr5	139006341	+	.	3	30	2594942_1	85.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GTA;MAPQ=60;MATEID=2594942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_138988501_139013501_172C;SPAN=3292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:74 GQ:85.7 PL:[85.7, 0.0, 92.3] SR:30 DR:3 LR:-85.58 LO:85.61);ALT=A[chr5:139006341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139028622	+	chr5	139059944	+	.	10	0	2595104_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2595104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:139028622(+)-5:139059944(-)__5_139037501_139062501D;SPAN=31322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:30 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:0 DR:10 LR:-24.88 LO:25.28);ALT=G[chr5:139059944[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139061032	+	chr5	139062446	+	.	3	12	2595137_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2595137_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_139062001_139087001_250C;SPAN=1414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:26 GQ:26 PL:[35.9, 0.0, 26.0] SR:12 DR:3 LR:-35.93 LO:35.93);ALT=G[chr5:139062446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139554873	+	chr5	139574029	+	.	28	6	2596020_1	81.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=2596020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_139552001_139577001_94C;SPAN=19156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:65 GQ:74.9 PL:[81.5, 0.0, 74.9] SR:6 DR:28 LR:-81.43 LO:81.43);ALT=G[chr5:139574029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139680169	+	chr5	139682625	+	.	7	10	2596090_1	26.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2596090_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_139674501_139699501_132C;SPAN=2456;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:10 DR:7 LR:-26.71 LO:31.54);ALT=T[chr5:139682625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139825561	+	chr5	139828793	+	.	2	4	2596518_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=2596518_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_139821501_139846501_146C;SPAN=3232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:52 GQ:2.6 PL:[2.6, 0.0, 121.4] SR:4 DR:2 LR:-2.417 LO:9.606);ALT=G[chr5:139828793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139927426	+	chr5	139928489	+	.	25	11	2596560_1	76.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2596560_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_139919501_139944501_78C;SPAN=1063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:58 GQ:63.5 PL:[76.7, 0.0, 63.5] SR:11 DR:25 LR:-76.77 LO:76.77);ALT=G[chr5:139928489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	139931771	+	chr5	139936732	+	.	0	21	2596567_1	54.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2596567_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_139919501_139944501_204C;SPAN=4961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:54 GQ:54.8 PL:[54.8, 0.0, 74.6] SR:21 DR:0 LR:-54.69 LO:54.89);ALT=T[chr5:139936732[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140025311	+	chr5	140026841	+	.	40	3	2596901_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2596901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_140017501_140042501_157C;SPAN=1530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:85 GQ:89.3 PL:[115.7, 0.0, 89.3] SR:3 DR:40 LR:-115.8 LO:115.8);ALT=C[chr5:140026841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140062809	+	chr5	140070439	+	.	0	15	2596803_1	41.0	.	EVDNC=ASSMB;HOMSEQ=CCTTGG;MAPQ=60;MATEID=2596803_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_140066501_140091501_106C;SPAN=7630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:30 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:15 DR:0 LR:-41.46 LO:41.46);ALT=G[chr5:140070439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140062855	+	chr5	140070844	+	.	10	0	2596804_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2596804_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140062855(+)-5:140070844(-)__5_140066501_140091501D;SPAN=7989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:29 GQ:25.1 PL:[25.1, 0.0, 44.9] SR:0 DR:10 LR:-25.15 LO:25.47);ALT=A[chr5:140070844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140080115	+	chr5	140081588	+	.	53	0	2596835_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2596835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140080115(+)-5:140081588(-)__5_140066501_140091501D;SPAN=1473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:65 GQ:0.9 PL:[158.4, 0.9, 0.0] SR:0 DR:53 LR:-167.0 LO:167.0);ALT=A[chr5:140081588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140080116	+	chr5	140083501	+	.	12	0	2596837_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2596837_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140080116(+)-5:140083501(-)__5_140066501_140091501D;SPAN=3385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:69 GQ:20.9 PL:[20.9, 0.0, 146.3] SR:0 DR:12 LR:-20.92 LO:26.38);ALT=G[chr5:140083501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140080498	+	chr5	140081590	+	.	0	25	2596839_1	65.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=2596839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_140066501_140091501_162C;SPAN=1092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:64 GQ:65.3 PL:[65.3, 0.0, 88.4] SR:25 DR:0 LR:-65.19 LO:65.41);ALT=G[chr5:140081590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140081714	+	chr5	140083502	+	.	4	42	2596842_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2596842_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_5_140066501_140091501_55C;SPAN=1788;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:76 GQ:58.7 PL:[124.7, 0.0, 58.7] SR:42 DR:4 LR:-125.9 LO:125.9);ALT=G[chr5:140083502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140081714	+	chr5	140084011	+	ATATTACTGCAATGTCTGTGACTGTGTGGTGAAGGACTCCATCAACTTTCTGGATCACATTAATGGAAAGAAAC	8	69	2596843_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATATTACTGCAATGTCTGTGACTGTGTGGTGAAGGACTCCATCAACTTTCTGGATCACATTAATGGAAAGAAAC;MAPQ=60;MATEID=2596843_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_140066501_140091501_55C;SPAN=2297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:84 GQ:9.3 PL:[221.1, 9.3, 0.0] SR:69 DR:8 LR:-226.8 LO:226.8);ALT=G[chr5:140084011[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140084191	+	chr5	140085214	+	.	10	0	2596847_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2596847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140084191(+)-5:140085214(-)__5_140066501_140091501D;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:0 DR:10 LR:-15.67 LO:21.47);ALT=T[chr5:140085214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	140594447	+	chr5	140558343	+	.	8	0	2597779_1	23.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2597779_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:140558343(-)-5:140594447(+)__5_140556501_140581501D;SPAN=36104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:7 GQ:2.1 PL:[23.1, 2.1, 0.0] SR:0 DR:8 LR:-23.11 LO:23.11);ALT=]chr5:140594447]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr5	140951609	+	chr5	140953059	+	.	0	10	2598427_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2598427_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_140948501_140973501_286C;SPAN=1450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:10 DR:0 LR:-19.19 LO:22.57);ALT=T[chr5:140953059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141011830	+	chr5	141579496	+	.	13	0	2599588_1	36.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=2599588_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:141011830(+)-5:141579496(-)__5_141561001_141586001D;SPAN=567666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:13 DP:12 GQ:3.3 PL:[36.3, 3.3, 0.0] SR:0 DR:13 LR:-36.31 LO:36.31);ALT=G[chr5:141579496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141014520	+	chr5	141016302	+	GATCATCTTCTTATAGAGACCGTAATGCAGGACCAGGCTATGGGTCAATGCCAGGCGATGGGGCTTCATAGGGTGTCCAGCT	12	14	2598576_1	52.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GATCATCTTCTTATAGAGACCGTAATGCAGGACCAGGCTATGGGTCAATGCCAGGCGATGGGGCTTCATAGGGTGTCCAGCT;MAPQ=60;MATEID=2598576_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_5_140997501_141022501_209C;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:63 GQ:52.4 PL:[52.4, 0.0, 98.6] SR:14 DR:12 LR:-52.25 LO:53.09);ALT=C[chr5:141016302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141303520	+	chr5	141304972	+	.	12	0	2599092_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2599092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:141303520(+)-5:141304972(-)__5_141291501_141316501D;SPAN=1452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:0 DR:12 LR:-22.81 LO:27.0);ALT=C[chr5:141304972[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141305093	+	chr5	141307715	+	.	0	8	2599097_1	9.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=2599097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141291501_141316501_143C;SPAN=2622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:8 DR:0 LR:-9.34 LO:16.4);ALT=G[chr5:141307715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141456960	+	chr13	82367698	+	C	12	62	5574246_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;INSERTION=C;MAPQ=41;MATEID=5574246_2;MATENM=1;NM=18;NUMPARTS=2;SCTG=c_13_82344501_82369501_305C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:38 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:62 DR:12 LR:-191.4 LO:191.4);ALT=C[chr13:82367698[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	141488602	+	chr5	141511371	+	.	0	81	2599505_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2599505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141487501_141512501_12C;SPAN=22769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:120 GQ:56.6 PL:[234.8, 0.0, 56.6] SR:81 DR:0 LR:-241.0 LO:241.0);ALT=G[chr5:141511371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141488604	+	chr5	141511772	+	.	11	0	2599506_1	9.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2599506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:141488604(+)-5:141511772(-)__5_141487501_141512501D;SPAN=23168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:0 DR:11 LR:-9.219 LO:21.81);ALT=T[chr5:141511772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141511460	+	chr5	141515295	+	CATATTTTGACTACAAGGATGAGTCTGGGTTTCCAAAGCCCCCATCTTACAATGTAGCTACAACACTGCCCAGTTATGATGAAGCGGAGAGGACCAAGGCTGAAGCTACTATCCCTTTGGTTCCTGGGAGA	0	30	2599537_1	92.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CATATTTTGACTACAAGGATGAGTCTGGGTTTCCAAAGCCCCCATCTTACAATGTAGCTACAACACTGCCCAGTTATGATGAAGCGGAGAGGACCAAGGCTGAAGCTACTATCCCTTTGGTTCCTGGGAGA;MAPQ=60;MATEID=2599537_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_141487501_141512501_25C;SPAN=3835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:32 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:30 DR:0 LR:-92.42 LO:92.42);ALT=G[chr5:141515295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141511908	+	chr5	141515295	+	.	5	6	2599450_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2599450_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_5_141512001_141537001_163C;SPAN=3387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:6 DR:5 LR:-26.24 LO:26.3);ALT=G[chr5:141515295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141515382	+	chr5	141517299	+	.	0	7	2599454_1	7.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2599454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141512001_141537001_243C;SPAN=1917;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:57 GQ:7.7 PL:[7.7, 0.0, 129.8] SR:7 DR:0 LR:-7.664 LO:14.24);ALT=A[chr5:141517299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141515382	+	chr5	141520128	+	.	2	3	2599455_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2599455_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141512001_141537001_77C;SPAN=4746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:56 GQ:1.4 PL:[1.4, 0.0, 133.4] SR:3 DR:2 LR:-1.333 LO:9.437);ALT=A[chr5:141520128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141520195	+	chr5	141524132	+	.	0	21	2599469_1	54.0	.	EVDNC=ASSMB;HOMSEQ=TTAGG;MAPQ=60;MATEID=2599469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141512001_141537001_181C;SPAN=3937;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:55 GQ:54.5 PL:[54.5, 0.0, 77.6] SR:21 DR:0 LR:-54.42 LO:54.67);ALT=G[chr5:141524132[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	141524241	+	chr5	141531294	+	.	3	15	2599474_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2599474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_141512001_141537001_141C;SPAN=7053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:63 GQ:39.2 PL:[39.2, 0.0, 111.8] SR:15 DR:3 LR:-39.05 LO:41.08);ALT=G[chr5:141531294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	175085185	+	chr5	175109708	+	.	16	0	2649616_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2649616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:175085185(+)-5:175109708(-)__5_175077001_175102001D;SPAN=24523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:19 GQ:1.8 PL:[49.5, 1.8, 0.0] SR:0 DR:16 LR:-51.04 LO:51.04);ALT=G[chr5:175109708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	175786923	+	chr5	175788605	+	.	0	16	2650953_1	44.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2650953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_175787501_175812501_11C;SPAN=1682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:31 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:16 DR:0 LR:-44.55 LO:44.55);ALT=T[chr5:175788605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	175825050	+	chr5	175843178	+	GAAACACATCTCCATTGACTGTGGTCCCCATGTCCTCAGAACCAG	3	16	2651116_1	59.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GAAACACATCTCCATTGACTGTGGTCCCCATGTCCTCAGAACCAG;MAPQ=60;MATEID=2651116_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_175836501_175861501_144C;SPAN=18128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:21 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:16 DR:3 LR:-57.84 LO:57.84);ALT=T[chr5:175843178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176258026	+	chr5	176259412	+	AAGTTC	59	57	2652125_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=AAGTTC;MAPQ=60;MATEID=2652125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176253001_176278001_254C;SPAN=1386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:31 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:57 DR:59 LR:-280.6 LO:280.6);ALT=A[chr5:176259412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176387587	+	chr5	176390181	+	.	44	27	2652209_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAAAAA;MAPQ=60;MATEID=2652209_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176375501_176400501_273C;SPAN=2594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:51 DP:725 GQ:27.7 PL:[0.0, 27.7, 1815.0] SR:27 DR:44 LR:28.07 LO:90.75);ALT=A[chr5:176390181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176402483	+	chr5	176409469	+	GTGCA	2	11	2652416_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;INSERTION=GTGCA;MAPQ=60;MATEID=2652416_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_176400001_176425001_221C;SPAN=6986;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:49 GQ:26.3 PL:[26.3, 0.0, 92.3] SR:11 DR:2 LR:-26.34 LO:28.41);ALT=T[chr5:176409469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176409624	+	chr5	176433651	+	.	20	5	2652429_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2652429_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176400001_176425001_311C;SPAN=24027;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:23 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:5 DR:20 LR:-69.32 LO:69.32);ALT=T[chr5:176433651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176560955	+	chr5	176562087	+	.	5	8	2652558_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=2652558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176547001_176572001_204C;SPAN=1132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:44 GQ:24.5 PL:[24.5, 0.0, 80.6] SR:8 DR:5 LR:-24.39 LO:26.15);ALT=T[chr5:176562087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176730323	+	chr5	176734781	+	.	0	8	2652962_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2652962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176718501_176743501_288C;SPAN=4458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:8 DR:0 LR:-10.42 LO:16.64);ALT=T[chr5:176734781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176759249	+	chr5	176764137	+	TTGGGCGACTTGAGGAAGTTGACGCTGGGCTCGATCTTGGTCCAGTCGATGCTCTCCTCGTCGGGCGTGTGCTCCACCATCAGCTGGAACAGCTTCATGGAGATGATGTCATGATTGT	3	20	2653040_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTGGGCGACTTGAGGAAGTTGACGCTGGGCTCGATCTTGGTCCAGTCGATGCTCTCCTCGTCGGGCGTGTGCTCCACCATCAGCTGGAACAGCTTCATGGAGATGATGTCATGATTGT;MAPQ=60;MATEID=2653040_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_176743001_176768001_123C;SPAN=4888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:76 GQ:48.8 PL:[48.8, 0.0, 134.6] SR:20 DR:3 LR:-48.73 LO:51.01);ALT=T[chr5:176764137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176759249	+	chr5	176761285	+	.	8	11	2653039_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2653039_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_176743001_176768001_123C;SPAN=2036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:58 GQ:47 PL:[47.0, 0.0, 93.2] SR:11 DR:8 LR:-47.01 LO:47.86);ALT=T[chr5:176761285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176761405	+	chr5	176764137	+	.	0	9	2653044_1	6.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2653044_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_176743001_176768001_123C;SPAN=2732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:85 GQ:6.8 PL:[6.8, 0.0, 198.2] SR:9 DR:0 LR:-6.68 LO:17.69);ALT=C[chr5:176764137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176765610	+	chr5	176778174	+	.	3	23	2653292_1	74.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=2653292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176767501_176792501_122C;SPAN=12564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:41 GQ:22.1 PL:[74.9, 0.0, 22.1] SR:23 DR:3 LR:-76.1 LO:76.1);ALT=G[chr5:176778174[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176765650	+	chr5	176778451	+	.	13	0	2653293_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2653293_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:176765650(+)-5:176778451(-)__5_176767501_176792501D;SPAN=12801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:56 GQ:27.8 PL:[27.8, 0.0, 107.0] SR:0 DR:13 LR:-27.74 LO:30.42);ALT=T[chr5:176778451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176785072	+	chr5	176793176	+	TCTGGCTGTGTCAGATGG	37	20	2653323_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCTGGCTGTGTCAGATGG;MAPQ=60;MATEID=2653323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176767501_176792501_208C;SPAN=8104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:38 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:20 DR:37 LR:-118.8 LO:118.8);ALT=T[chr5:176793176[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176919679	+	chr5	176923418	+	.	0	13	2653342_1	28.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2653342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_176914501_176939501_224C;SPAN=3739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:54 GQ:28.4 PL:[28.4, 0.0, 101.0] SR:13 DR:0 LR:-28.28 LO:30.66);ALT=C[chr5:176923418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	176919728	+	chr5	176924539	+	.	28	0	2653343_1	75.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2653343_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:176919728(+)-5:176924539(-)__5_176914501_176939501D;SPAN=4811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:64 GQ:75.2 PL:[75.2, 0.0, 78.5] SR:0 DR:28 LR:-75.09 LO:75.1);ALT=A[chr5:176924539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177019400	+	chr5	177020649	+	AAACTACCGGACGCAGCTGTATGACAAGCAGCGGGAGGAGTACCAGCCGGCCACCCCGGGGCTTGGCATGTTTGTGGAGGTGAAGGACCCAGAGGACA	15	98	2653474_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=AAACTACCGGACGCAGCTGTATGACAAGCAGCGGGAGGAGTACCAGCCGGCCACCCCGGGGCTTGGCATGTTTGTGGAGGTGAAGGACCCAGAGGACA;MAPQ=60;MATEID=2653474_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_177012501_177037501_269C;SPAN=1249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:89 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:98 DR:15 LR:-307.0 LO:307.0);ALT=G[chr5:177020649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177027263	+	chr5	177031177	+	.	24	3	2653499_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=2653499_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_177012501_177037501_195C;SPAN=3914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:55 GQ:61.1 PL:[71.0, 0.0, 61.1] SR:3 DR:24 LR:-70.95 LO:70.95);ALT=T[chr5:177031177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177580808	-	chr10	93976191	+	.	41	0	2654873_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2654873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:177580808(-)-10:93976191(-)__5_177576001_177601001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:74 GQ:62.6 PL:[115.4, 0.0, 62.6] SR:0 DR:41 LR:-116.1 LO:116.1);ALT=[chr10:93976191[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr5	177595870	+	chr18	46198355	+	.	14	40	6616153_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=AGCCACTGTG;MAPQ=60;MATEID=6616153_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_46182501_46207501_312C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:17 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:40 DR:14 LR:-125.4 LO:125.4);ALT=G[chr18:46198355[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr5	177635919	+	chr5	177638891	+	.	0	8	2654943_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=2654943_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_177625001_177650001_212C;SPAN=2972;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:69 GQ:7.7 PL:[7.7, 0.0, 159.5] SR:8 DR:0 LR:-7.714 LO:16.06);ALT=G[chr5:177638891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177636450	+	chr5	177637552	+	.	0	6	2654945_1	2.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=2654945_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_177625001_177650001_44C;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:64 GQ:2.6 PL:[2.6, 0.0, 151.1] SR:6 DR:0 LR:-2.467 LO:11.46);ALT=T[chr5:177637552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	177821913	+	chr5	177823871	+	.	15	0	2655325_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2655325_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:177821913(+)-5:177823871(-)__5_177821001_177846001D;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:44 GQ:37.7 PL:[37.7, 0.0, 67.4] SR:0 DR:15 LR:-37.59 LO:38.11);ALT=T[chr5:177823871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	178050451	+	chr5	178053969	+	.	11	0	2655632_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2655632_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:178050451(+)-5:178053969(-)__5_178041501_178066501D;SPAN=3518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:59 GQ:20.3 PL:[20.3, 0.0, 122.6] SR:0 DR:11 LR:-20.33 LO:24.55);ALT=T[chr5:178053969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	178109066	+	chr5	178113412	+	.	24	30	2655782_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GAGAT;MAPQ=60;MATEID=2655782_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_178090501_178115501_232C;SPAN=4346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:12 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:30 DR:24 LR:-138.6 LO:138.6);ALT=T[chr5:178113412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	178860409	-	chr5	179217043	+	.	10	0	2658113_1	29.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=2658113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:178860409(-)-5:179217043(-)__5_179193001_179218001D;SPAN=356634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:14 GQ:2.9 PL:[29.3, 0.0, 2.9] SR:0 DR:10 LR:-30.22 LO:30.22);ALT=[chr5:179217043[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr5	178860539	+	chr5	179216893	-	.	10	0	2658114_1	28.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2658114_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:178860539(+)-5:179216893(+)__5_179193001_179218001D;SPAN=356354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:18 GQ:14.9 PL:[28.1, 0.0, 14.9] SR:0 DR:10 LR:-28.33 LO:28.33);ALT=G]chr5:179216893];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr5	179046410	+	chr5	179047892	+	.	4	7	2657769_1	18.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2657769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179046001_179071001_326C;SPAN=1482;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:66 GQ:18.5 PL:[18.5, 0.0, 140.6] SR:7 DR:4 LR:-18.43 LO:23.96);ALT=T[chr5:179047892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179048399	+	chr5	179050038	+	.	0	23	2657775_1	62.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2657775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179046001_179071001_12C;SPAN=1639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:49 GQ:56 PL:[62.6, 0.0, 56.0] SR:23 DR:0 LR:-62.67 LO:62.67);ALT=C[chr5:179050038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179048440	+	chr5	179050611	+	.	20	0	2657776_1	50.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=2657776_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179048440(+)-5:179050611(-)__5_179046001_179071001D;SPAN=2171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:59 GQ:50 PL:[50.0, 0.0, 92.9] SR:0 DR:20 LR:-50.04 LO:50.75);ALT=A[chr5:179050611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179126103	+	chr5	179132678	+	.	68	14	2657864_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2657864_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_5_179119501_179144501_79C;SPAN=6575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:56 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:14 DR:68 LR:-208.0 LO:208.0);ALT=G[chr5:179132678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179126124	+	chr5	179133256	+	.	8	0	2657865_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2657865_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179126124(+)-5:179133256(-)__5_179119501_179144501D;SPAN=7132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.59 LO:17.19);ALT=G[chr5:179133256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179137098	+	chr5	179143105	+	.	12	0	2657893_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2657893_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179137098(+)-5:179143105(-)__5_179119501_179144501D;SPAN=6007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=G[chr5:179143105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179147562	+	chr5	179149803	+	.	5	6	2657923_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2657923_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_5_179144001_179169001_179C;SPAN=2241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:6 DR:5 LR:-14.27 LO:19.37);ALT=G[chr5:179149803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179150055	+	chr5	179151655	+	.	11	0	2657931_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2657931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179150055(+)-5:179151655(-)__5_179144001_179169001D;SPAN=1600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:52 GQ:22.4 PL:[22.4, 0.0, 101.6] SR:0 DR:11 LR:-22.22 LO:25.23);ALT=A[chr5:179151655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179151833	+	chr5	179155589	+	.	8	0	2657938_1	11.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2657938_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179151833(+)-5:179155589(-)__5_179144001_179169001D;SPAN=3756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=G[chr5:179155589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179153766	+	chr5	179155601	+	.	8	0	2657948_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2657948_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179153766(+)-5:179155601(-)__5_179144001_179169001D;SPAN=1835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=G[chr5:179155601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179221139	+	chr5	179222583	+	.	56	16	2658165_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2658165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179217501_179242501_156C;SPAN=1444;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:50 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:16 DR:56 LR:-168.3 LO:168.3);ALT=G[chr5:179222583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179248141	+	chr5	179249957	+	.	0	28	2658346_1	63.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=2658346_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179242001_179267001_78C;SPAN=1816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:108 GQ:63.2 PL:[63.2, 0.0, 198.5] SR:28 DR:0 LR:-63.17 LO:67.09);ALT=G[chr5:179249957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179326308	+	chr5	179334702	+	ACACGCCACTGTCCAGTAGACCTGGGAGTCCTGGGTCTGGTGCAGGATGCGGTAAGGGGCCACGCGGGCACTGGAGTCCAGCACCACGTCCAGGGTGCCCACGAGAAG	0	19	2658309_1	54.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=ACACGCCACTGTCCAGTAGACCTGGGAGTCCTGGGTCTGGTGCAGGATGCGGTAAGGGGCCACGCGGGCACTGGAGTCCAGCACCACGTCCAGGGTGCCCACGAGAAG;MAPQ=60;MATEID=2658309_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_179315501_179340501_250C;SPAN=8394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:29 GQ:15.2 PL:[54.8, 0.0, 15.2] SR:19 DR:0 LR:-56.08 LO:56.08);ALT=C[chr5:179334702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179331858	+	chr5	179334794	+	.	13	0	2658323_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2658323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:179331858(+)-5:179334794(-)__5_179315501_179340501D;SPAN=2936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:28 GQ:32 PL:[35.3, 0.0, 32.0] SR:0 DR:13 LR:-35.33 LO:35.33);ALT=C[chr5:179334794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179382669	+	chr5	179390470	+	.	4	53	2658692_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2658692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179364501_179389501_258C;SPAN=7801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:37 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:53 DR:4 LR:-168.3 LO:168.3);ALT=C[chr5:179390470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179390564	+	chr5	179393806	+	.	0	44	2658454_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2658454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179389001_179414001_166C;SPAN=3242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:83 GQ:76.7 PL:[122.9, 0.0, 76.7] SR:44 DR:0 LR:-123.3 LO:123.3);ALT=T[chr5:179393806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179397506	+	chr5	179405202	+	.	3	8	2658467_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2658467_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_179389001_179414001_295C;SPAN=7696;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:8 DR:3 LR:-19.51 LO:24.29);ALT=C[chr5:179405202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179405287	+	chr5	179407128	+	.	2	9	2658481_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2658481_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_179389001_179414001_295C;SPAN=1841;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:9 DR:2 LR:-17.3 LO:21.94);ALT=T[chr5:179407128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179407202	+	chr5	179440061	+	.	3	6	2658748_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2658748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179438001_179463001_290C;SPAN=32859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:6 DR:3 LR:-16.93 LO:18.66);ALT=T[chr5:179440061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179440314	+	chr5	179467452	+	.	6	8	2658752_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=2658752_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179438001_179463001_117C;SPAN=27138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:29 GQ:31.7 PL:[31.7, 0.0, 38.3] SR:8 DR:6 LR:-31.76 LO:31.79);ALT=G[chr5:179467452[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	179467649	+	chr5	179498456	+	.	38	52	2658587_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2658587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_179487001_179512001_255C;SPAN=30807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:25 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:52 DR:38 LR:-217.9 LO:217.9);ALT=T[chr5:179498456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180220099	+	chr5	180230600	+	.	0	7	2660053_1	16.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=2660053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_180222001_180247001_93C;SPAN=10501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:26 GQ:16.1 PL:[16.1, 0.0, 45.8] SR:7 DR:0 LR:-16.06 LO:16.91);ALT=T[chr5:180230600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180665241	+	chr5	180666485	+	TGCCTCCAGAAGCACAGAGGGATCCATCTGGAGAGACAGTCACCGTGTTCAGATAGCCTGTGTGGCCAATGTGGTTGGTCTTCAGCTTGCAGTTAGCCAGGTTCCAT	2	125	2660753_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TAAAGGTGTTTGCCTTCGTTGAGATCCCATAACATGGCCTGGCCATCCTTGCCTCCAGAAGCACAGAGGGATCCATCTGGAGAGACAGTCACCGTGTTCAGATAGCCTGTGTGGCCAATGTGGTTGGTCTTCAGCTTGCAGTTAGCCAGGTTCCATACCT;INSERTION=TGCCTCCAGAAGCACAGAGGGATCCATCTGGAGAGACAGTCACCGTGTTCAGATAGCCTGTGTGGCCAATGTGGTTGGTCTTCAGCTTGCAGTTAGCCAGGTTCCAT;MAPQ=60;MATEID=2660753_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_5_180663001_180688001_19C;SECONDARY;SPAN=1244;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:106 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:125 DR:2 LR:-373.0 LO:373.0);ALT=T[chr5:180666485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180666202	+	chr5	180668490	+	.	11	0	2660757_1	17.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2660757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:180666202(+)-5:180668490(-)__5_180663001_180688001D;SPAN=2288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:71 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:0 DR:11 LR:-17.08 LO:23.58);ALT=T[chr5:180668490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180666584	+	chr5	180668491	+	.	18	47	2660758_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2660758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_180663001_180688001_52C;SPAN=1907;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:91 GQ:51.5 PL:[167.0, 0.0, 51.5] SR:47 DR:18 LR:-170.0 LO:170.0);ALT=T[chr5:180668491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180666629	+	chr5	180669282	+	.	13	0	2660759_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2660759_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:180666629(+)-5:180669282(-)__5_180663001_180688001D;SPAN=2653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:13 DP:505 GQ:93.6 PL:[0.0, 93.6, 1413.0] SR:0 DR:13 LR:93.9 LO:17.37);ALT=A[chr5:180669282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180668687	+	chr5	180670762	+	.	56	0	2660767_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2660767_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:180668687(+)-5:180670762(-)__5_180663001_180688001D;SPAN=2075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:492 GQ:51.8 PL:[51.8, 0.0, 1141.0] SR:0 DR:56 LR:-51.56 LO:111.9);ALT=T[chr5:180670762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180669347	+	chr5	180670692	+	.	127	131	2660770_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2660770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_180663001_180688001_277C;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:195 DP:604 GQ:99 PL:[480.3, 0.0, 985.3] SR:131 DR:127 LR:-480.1 LO:489.6);ALT=T[chr5:180670692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	180688385	+	chr5	180690625	+	.	21	7	2660804_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=2660804_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_180687501_180712501_184C;SPAN=2240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:61 GQ:62.9 PL:[62.9, 0.0, 82.7] SR:7 DR:21 LR:-62.7 LO:62.89);ALT=G[chr5:180690625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	292610	+	chr6	311877	+	.	8	0	2662042_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2662042_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:292610(+)-6:311877(-)__6_269501_294501D;SPAN=19267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:0 DR:8 LR:-10.97 LO:16.77);ALT=G[chr6:311877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	292610	+	chr6	345851	+	.	12	0	2662222_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2662222_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:292610(+)-6:345851(-)__6_343001_368001D;SPAN=53241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:57 GQ:24.2 PL:[24.2, 0.0, 113.3] SR:0 DR:12 LR:-24.17 LO:27.5);ALT=G[chr6:345851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	345928	+	chr6	348102	+	.	0	17	2662244_1	14.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=2662244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_343001_368001_173C;SPAN=2174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:154 GQ:14.6 PL:[14.6, 0.0, 357.8] SR:17 DR:0 LR:-14.39 LO:33.74);ALT=G[chr6:348102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	666376	+	chr6	667822	+	.	0	50	2663149_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2663149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_661501_686501_35C;SPAN=1446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:80 GQ:50.9 PL:[143.3, 0.0, 50.9] SR:50 DR:0 LR:-145.8 LO:145.8);ALT=A[chr6:667822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	1274201	-	chr6	1275263	+	.	11	0	2665744_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2665744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:1274201(-)-6:1275263(-)__6_1249501_1274501D;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=[chr6:1275263[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	1624809	+	chr6	1626361	+	.	21	0	2666626_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2666626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:1624809(+)-6:1626361(-)__6_1617001_1642001D;SPAN=1552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:115 GQ:38.3 PL:[38.3, 0.0, 239.6] SR:0 DR:21 LR:-38.17 LO:46.66);ALT=G[chr6:1626361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2125022	+	chr6	2245714	+	.	12	0	2668549_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2668549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2125022(+)-6:2245714(-)__6_2229501_2254501D;SPAN=120692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=T[chr6:2245714[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2246164	+	chr6	2249069	+	.	12	10	2668619_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2668619_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2229501_2254501_282C;SPAN=2905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:102 GQ:28.7 PL:[28.7, 0.0, 216.8] SR:10 DR:12 LR:-28.48 LO:37.03);ALT=G[chr6:2249069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2249160	+	chr6	2263833	+	.	0	11	2668640_1	19.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2668640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2229501_2254501_436C;SPAN=14673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:11 DR:0 LR:-19.51 LO:24.29);ALT=G[chr6:2263833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2834248	+	chr6	2836090	+	.	67	39	2670598_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2670598_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2817501_2842501_366C;SPAN=1842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:86 DP:130 GQ:67.1 PL:[248.6, 0.0, 67.1] SR:39 DR:67 LR:-254.5 LO:254.5);ALT=T[chr6:2836090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2836486	+	chr6	2838782	+	TCTGTCTGTCCTTTGACCCACTGGTTTATGGTCTTCCTTGCATCTTCAGAGGCATGCTGAAAATCCACACTGGCCAGGTCAGCACCATATGTTTTCTGAGTCGAAACCAAGAACT	16	83	2670612_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCTGTCTGTCCTTTGACCCACTGGTTTATGGTCTTCCTTGCATCTTCAGAGGCATGCTGAAAATCCACACTGGCCAGGTCAGCACCATATGTTTTCTGAGTCGAAACCAAGAACT;MAPQ=60;MATEID=2670612_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_2817501_2842501_174C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:130 GQ:63.8 PL:[251.9, 0.0, 63.8] SR:83 DR:16 LR:-258.3 LO:258.3);ALT=T[chr6:2838782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2836486	+	chr6	2838115	+	.	18	30	2670611_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2670611_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTGTCTGT;SCTG=c_6_2817501_2842501_174C;SPAN=1629;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:119 GQ:60 PL:[60.0, 0.0, 89.9] SR:30 DR:18 LR:-59.76 LO:60.29);ALT=T[chr6:2838115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2838275	+	chr6	2842045	+	.	15	0	2670625_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2670625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2838275(+)-6:2842045(-)__6_2817501_2842501D;SPAN=3770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:15 DP:365 GQ:49.1 PL:[0.0, 49.1, 983.6] SR:0 DR:15 LR:49.37 LO:23.11);ALT=C[chr6:2842045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2838922	+	chr6	2840653	+	.	2	95	2670627_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2670627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2817501_2842501_5C;SPAN=1731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:315 GQ:99 PL:[235.0, 0.0, 528.8] SR:95 DR:2 LR:-234.9 LO:241.1);ALT=T[chr6:2840653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2838979	+	chr6	2842045	+	.	120	0	2670628_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2670628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2838979(+)-6:2842045(-)__6_2817501_2842501D;SPAN=3066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:120 DP:362 GQ:99 PL:[298.3, 0.0, 578.9] SR:0 DR:120 LR:-298.0 LO:303.0);ALT=C[chr6:2842045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2840854	+	chr6	2842043	+	.	136	0	2670639_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2670639_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2840854(+)-6:2842043(-)__6_2817501_2842501D;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:136 DP:333 GQ:99 PL:[358.9, 0.0, 448.0] SR:0 DR:136 LR:-358.7 LO:359.3);ALT=G[chr6:2842043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2949305	+	chr6	2955758	+	TGCTGACTTTAAACAGTCTCTCCTCGGTGTTCTCCTTGTCAAACTGTTCATCCCAGTTTCCTCTGAAATAGACAGCATTCACCAGAACCAGCCTTGTCAATGGATCCACTGAGCCCGGAGAGAGCAACTCCGCAATTTTACCTTCTGTCTTTTCAGCTACCCAGGTGTTTATGTGTTTTCTGGACTTCTCTACGGCGCTGATAAAGTCAAGCTCCTCCATCTCTGCTTGGTAGAATTTTTGGCAGGAATCTCTAAAAGA	0	27	2670885_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=TGCTGACTTTAAACAGTCTCTCCTCGGTGTTCTCCTTGTCAAACTGTTCATCCCAGTTTCCTCTGAAATAGACAGCATTCACCAGAACCAGCCTTGTCAATGGATCCACTGAGCCCGGAGAGAGCAACTCCGCAATTTTACCTTCTGTCTTTTCAGCTACCCAGGTGTTTATGTGTTTTCTGGACTTCTCTACGGCGCTGATAAAGTCAAGCTCCTCCATCTCTGCTTGGTAGAATTTTTGGCAGGAATCTCTAAAAGA;MAPQ=60;MATEID=2670885_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_2940001_2965001_317C;SPAN=6453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:121 GQ:56.6 PL:[56.6, 0.0, 234.8] SR:27 DR:0 LR:-56.35 LO:62.65);ALT=T[chr6:2955758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2949305	+	chr6	2953278	+	.	12	16	2670884_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2670884_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_2940001_2965001_317C;SPAN=3973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:107 GQ:37.1 PL:[37.1, 0.0, 221.9] SR:16 DR:12 LR:-37.03 LO:44.67);ALT=T[chr6:2953278[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2953422	+	chr6	2954824	+	.	0	5	2670905_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=2670905_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_2940001_2965001_317C;SPAN=1402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:85 GQ:6.3 PL:[0.0, 6.3, 217.8] SR:5 DR:0 LR:6.524 LO:8.497);ALT=T[chr6:2954824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2955907	+	chr6	2959402	+	.	9	31	2670914_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2670914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2940001_2965001_75C;SPAN=3495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:124 GQ:98.6 PL:[98.6, 0.0, 200.9] SR:31 DR:9 LR:-98.45 LO:100.4);ALT=G[chr6:2959402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2955953	+	chr6	2971764	+	.	10	0	2671031_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2671031_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2955953(+)-6:2971764(-)__6_2964501_2989501D;SPAN=15811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=T[chr6:2971764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2955956	+	chr6	2971348	+	.	16	0	2671032_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2671032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:2955956(+)-6:2971348(-)__6_2964501_2989501D;SPAN=15392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:40 GQ:41.9 PL:[41.9, 0.0, 55.1] SR:0 DR:16 LR:-41.98 LO:42.08);ALT=A[chr6:2971348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2959576	+	chr6	2971765	+	.	37	13	2671034_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=2671034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2964501_2989501_302C;SPAN=12189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:52 GQ:0.6 PL:[125.4, 0.6, 0.0] SR:13 DR:37 LR:-131.9 LO:131.9);ALT=C[chr6:2971765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	2959579	+	chr6	2971349	+	.	22	8	2671035_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=2671035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_2964501_2989501_167C;SPAN=11770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:40 GQ:28.7 PL:[68.3, 0.0, 28.7] SR:8 DR:22 LR:-69.27 LO:69.27);ALT=G[chr6:2971349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	3000319	+	chr6	3006700	+	.	0	16	2671170_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2671170_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_2989001_3014001_428C;SPAN=6381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:130 GQ:17.6 PL:[17.6, 0.0, 298.1] SR:16 DR:0 LR:-17.6 LO:32.56);ALT=G[chr6:3006700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	3017219	+	chr6	3019711	+	.	3	9	2671239_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2671239_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_3013501_3038501_378C;SPAN=2492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:133 GQ:3.8 PL:[3.8, 0.0, 317.3] SR:9 DR:3 LR:-3.579 LO:22.71);ALT=G[chr6:3019711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	3259430	+	chr6	3267825	+	.	2	4	2672321_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2672321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_3258501_3283501_321C;SPAN=8395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:116 GQ:14.7 PL:[0.0, 14.7, 310.2] SR:4 DR:2 LR:14.92 LO:7.808);ALT=C[chr6:3267825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	3259431	+	chr6	3263918	+	.	0	18	2672322_1	28.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=2672322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_3258501_3283501_82C;SPAN=4487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:116 GQ:28.1 PL:[28.1, 0.0, 252.5] SR:18 DR:0 LR:-27.99 LO:38.59);ALT=G[chr6:3263918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	3263993	+	chr6	3267822	+	.	0	13	2672335_1	9.0	.	EVDNC=ASSMB;HOMSEQ=TAG;MAPQ=60;MATEID=2672335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_3258501_3283501_183C;SPAN=3829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:123 GQ:9.8 PL:[9.8, 0.0, 287.0] SR:13 DR:0 LR:-9.589 LO:25.54);ALT=G[chr6:3267822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131934791	+	chr6	3978390	+	.	19	0	4721038_1	56.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=4721038_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:3978390(-)-10:131934791(+)__10_131932501_131957501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:16 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:0 DR:19 LR:-56.11 LO:56.11);ALT=]chr10:131934791]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	4021701	+	chr6	4031793	+	.	23	6	2674905_1	57.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2674905_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_4018001_4043001_15C;SPAN=10092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:94 GQ:57.2 PL:[57.2, 0.0, 169.4] SR:6 DR:23 LR:-57.06 LO:60.23);ALT=G[chr6:4031793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	4130796	+	chr6	4133782	+	TGGGCAGGCTGCCAAGGGCATTCCATGCGTCCCATTTGGCCTTGTTGATCAAGTCAAATACACCTGGTTTGGGCATGTTACAAGGTCCTTCAGTGG	0	23	2675300_1	47.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=TGGGCAGGCTGCCAAGGGCATTCCATGCGTCCCATTTGGCCTTGTTGATCAAGTCAAATACACCTGGTTTGGGCATGTTACAAGGTCCTTCAGTGG;MAPQ=60;MATEID=2675300_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_6_4116001_4141001_218C;SPAN=2986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:106 GQ:47.3 PL:[47.3, 0.0, 209.0] SR:23 DR:0 LR:-47.21 LO:53.05);ALT=T[chr6:4133782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	4131141	+	chr6	4135743	+	.	12	0	2675303_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2675303_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:4131141(+)-6:4135743(-)__6_4116001_4141001D;SPAN=4602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:96 GQ:13.7 PL:[13.7, 0.0, 218.3] SR:0 DR:12 LR:-13.6 LO:24.51);ALT=A[chr6:4135743[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	4133940	+	chr6	4135743	+	.	17	0	2675316_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2675316_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:4133940(+)-6:4135743(-)__6_4116001_4141001D;SPAN=1803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:94 GQ:30.8 PL:[30.8, 0.0, 195.8] SR:0 DR:17 LR:-30.65 LO:37.69);ALT=A[chr6:4135743[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	4475582	-	chr8	125476342	+	.	2	2	2676341_1	0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGAG;MAPQ=60;MATEID=2676341_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_4459001_4484001_296C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:49 GQ:0 PL:[0.0, 0.0, 118.8] SR:2 DR:2 LR:0.0713 LO:7.387);ALT=[chr8:125476342[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	5002527	+	chr6	5004184	+	.	9	0	2678236_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2678236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:5002527(+)-6:5004184(-)__6_4998001_5023001D;SPAN=1657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:0 DR:9 LR:-1.262 LO:16.82);ALT=A[chr6:5004184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	5037249	+	chr6	5039187	+	AAAATCTGCTTC	0	50	2678688_1	99.0	.	EVDNC=ASSMB;INSERTION=AAAATCTGCTTC;MAPQ=60;MATEID=2678688_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_5022501_5047501_409C;SPAN=1938;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:35 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:50 DR:0 LR:-148.5 LO:148.5);ALT=T[chr6:5039187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	5109775	+	chr6	5260914	+	.	14	0	2679257_1	32.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2679257_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:5109775(+)-6:5260914(-)__6_5243001_5268001D;SPAN=151139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:52 GQ:32.3 PL:[32.3, 0.0, 91.7] SR:0 DR:14 LR:-32.13 LO:33.82);ALT=T[chr6:5260914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	5216973	+	chr6	5260881	+	.	9	6	2679259_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2679259_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_5243001_5268001_420C;SPAN=43908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:42 GQ:31.7 PL:[31.7, 0.0, 68.0] SR:6 DR:9 LR:-31.53 LO:32.35);ALT=T[chr6:5260881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	5261893	+	chr6	5368782	+	.	19	6	2679575_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2679575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_5365501_5390501_68C;SPAN=106889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:68 GQ:44.3 PL:[44.3, 0.0, 120.2] SR:6 DR:19 LR:-44.3 LO:46.26);ALT=G[chr6:5368782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	5852781	-	chr13	21899458	+	.	13	0	5414304_1	34.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5414304_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:5852781(-)-13:21899458(-)__13_21878501_21903501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:31 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:0 DR:13 LR:-34.51 LO:34.54);ALT=[chr13:21899458[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	5853738	+	chr13	21899458	-	.	11	0	5414306_1	28.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5414306_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:5853738(+)-13:21899458(+)__13_21878501_21903501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:31 GQ:28.1 PL:[28.1, 0.0, 44.6] SR:0 DR:11 LR:-27.91 LO:28.19);ALT=T]chr13:21899458];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	6243461	-	chr22	49000956	+	.	8	0	7336747_1	7.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7336747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6243461(-)-22:49000956(-)__22_49000001_49025001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=[chr22:49000956[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	6267043	+	chr6	6305582	+	.	3	4	2683110_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=2683110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_6296501_6321501_27C;SPAN=38539;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:53 GQ:5.6 PL:[5.6, 0.0, 121.1] SR:4 DR:3 LR:-5.447 LO:11.98);ALT=C[chr6:6305582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6312664	+	chr6	9434113	-	.	20	75	2683165_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACTTTGG;MAPQ=60;MATEID=2683165_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_6_6296501_6321501_279C;SPAN=3121449;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:27 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:75 DR:20 LR:-247.6 LO:247.6);ALT=G]chr6:9434113];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	6318948	+	chr6	6320831	+	.	12	0	2683194_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2683194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6318948(+)-6:6320831(-)__6_6296501_6321501D;SPAN=1883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:121 GQ:7.1 PL:[7.1, 0.0, 284.3] SR:0 DR:12 LR:-6.83 LO:23.22);ALT=A[chr6:6320831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6589103	+	chr6	6625158	+	.	72	60	2683742_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2683742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_6566001_6591001_182C;SPAN=36055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:74 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:60 DR:72 LR:-307.0 LO:307.0);ALT=G[chr6:6625158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6589120	+	chr6	6626525	+	.	46	0	2683744_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2683744_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6589120(+)-6:6626525(-)__6_6566001_6591001D;SPAN=37405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:54 GQ:7.8 PL:[145.2, 7.8, 0.0] SR:0 DR:46 LR:-147.4 LO:147.4);ALT=C[chr6:6626525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6625246	+	chr6	6626526	+	.	9	110	2683786_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2683786_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_6615001_6640001_91C;SPAN=1280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:118 DP:162 GQ:45.5 PL:[345.8, 0.0, 45.5] SR:110 DR:9 LR:-358.7 LO:358.7);ALT=G[chr6:6626526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	6626654	+	chr6	6654774	+	AGCAGATTTACTATGCTGGGCCTGTCAATAATCCTGAATTTACTATTCCT	11	41	2683903_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=AGCAGATTTACTATGCTGGGCCTGTCAATAATCCTGAATTTACTATTCCT;MAPQ=60;MATEID=2683903_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_6639501_6664501_88C;SPAN=28120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:61 GQ:3 PL:[151.8, 3.0, 0.0] SR:41 DR:11 LR:-157.9 LO:157.9);ALT=G[chr6:6654774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7299056	+	chr6	7301542	+	.	0	10	2686565_1	17.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2686565_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_7301001_7326001_29C;SPAN=2486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:10 DR:0 LR:-17.03 LO:21.86);ALT=C[chr6:7301542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7301807	+	chr6	7303783	+	.	5	4	2686570_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2686570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_7301001_7326001_181C;SPAN=1976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:4 DR:5 LR:0.9554 LO:14.66);ALT=T[chr6:7303783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7303915	+	chr6	7313328	+	.	8	0	2686578_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2686578_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:7303915(+)-6:7313328(-)__6_7301001_7326001D;SPAN=9413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:0 DR:8 LR:3.123 LO:14.39);ALT=A[chr6:7313328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7310308	+	chr6	7313328	+	.	43	0	2686608_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2686608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:7310308(+)-6:7313328(-)__6_7301001_7326001D;SPAN=3020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:99 GQ:99 PL:[115.1, 0.0, 125.0] SR:0 DR:43 LR:-115.1 LO:115.1);ALT=A[chr6:7313328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	7590647	+	chr6	7593965	+	.	0	7	2687803_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2687803_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_7570501_7595501_4C;SPAN=3318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:120 GQ:9.3 PL:[0.0, 9.3, 310.2] SR:7 DR:0 LR:9.404 LO:11.87);ALT=G[chr6:7593965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	8097702	+	chr6	8102668	+	.	38	8	2689588_1	58.0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2689588_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCGCTCGC;SCTG=c_6_8085001_8110001_71C;SPAN=4966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:96 GQ:58.3 PL:[58.3, 0.0, 62.2] SR:8 DR:38 LR:-57.99 LO:58.02);ALT=T[chr6:8102668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10695302	+	chr6	10697555	+	.	7	4	2698044_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2698044_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10682001_10707001_118C;SPAN=2253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:4 DR:7 LR:-3.971 LO:17.23);ALT=G[chr6:10697555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10697419	-	chr6	10702601	+	ACTGTGATGCACTAGAGCCCCATGCTCAATCTTCTTTTTCATGTCATAAATGTGAATTGTTTCATCTTTGCTCCCAGTGACCACAAAACGACTATTTACAGCTACTGCTGACAAGGAGGCAGTGTGAGCATGGTGAGTGAAGTCAGCCACAAGAGTCCATTGCTGCTGAAGATGAAAACATACAATTAATGCCAGTCACACCACAGTTCTACCAACTCTATCCACTGG	0	20	2698050_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TAGTTTTCATGAATC;INSERTION=ACTGTGATGCACTAGAGCCCCATGCTCAATCTTCTTTTTCATGTCATAAATGTGAATTGTTTCATCTTTGCTCCCAGTGACCACAAAACGACTATTTACAGCTACTGCTGACAAGGAGGCAGTGTGAGCATGGTGAGTGAAGTCAGCCACAAGAGTCCATTGCTGCTGAAGATGAAAACATACAATTAATGCCAGTCACACCACAGTTCTACCAACTCTATCCACTGG;MAPQ=60;MATEID=2698050_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_10682001_10707001_6C;SPAN=5182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:102 GQ:38.6 PL:[38.6, 0.0, 206.9] SR:20 DR:0 LR:-38.39 LO:45.13);ALT=[chr6:10702601[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	10723474	+	chr6	10724788	+	.	36	17	2698243_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2698243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_394C;SPAN=1314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:155 GQ:99 PL:[113.3, 0.0, 261.8] SR:17 DR:36 LR:-113.2 LO:116.4);ALT=G[chr6:10724788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723474	+	chr6	10725193	+	.	46	3	2698244_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2698244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_153C;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:180 GQ:99 PL:[113.0, 0.0, 324.2] SR:3 DR:46 LR:-113.0 LO:118.6);ALT=G[chr6:10725193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723511	+	chr6	10726136	+	.	32	0	2698248_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2698248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10723511(+)-6:10726136(-)__6_10706501_10731501D;SPAN=2625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:106 GQ:77 PL:[77.0, 0.0, 179.3] SR:0 DR:32 LR:-76.91 LO:79.21);ALT=C[chr6:10726136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10723513	+	chr10	70304558	-	.	25	0	2698249_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2698249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10723513(+)-10:70304558(+)__6_10706501_10731501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:50 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:0 DR:25 LR:-69.1 LO:69.1);ALT=T]chr10:70304558];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	10723515	+	chr6	10728870	+	.	13	0	2698250_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2698250_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10723515(+)-6:10728870(-)__6_10706501_10731501D;SPAN=5355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:104 GQ:14.9 PL:[14.9, 0.0, 236.0] SR:0 DR:13 LR:-14.74 LO:26.55);ALT=T[chr6:10728870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10726241	+	chr6	10728871	+	.	0	33	2698267_1	79.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2698267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_60C;SPAN=2630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:110 GQ:79.1 PL:[79.1, 0.0, 188.0] SR:33 DR:0 LR:-79.13 LO:81.57);ALT=G[chr6:10728871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10728960	+	chr6	10730845	+	.	7	11	2698282_1	27.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=2698282_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_10706501_10731501_406C;SPAN=1885;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:107 GQ:27.2 PL:[27.2, 0.0, 231.8] SR:11 DR:7 LR:-27.13 LO:36.64);ALT=G[chr6:10730845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10748147	+	chr6	10751363	+	.	25	0	2698155_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2698155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10748147(+)-6:10751363(-)__6_10731001_10756001D;SPAN=3216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:109 GQ:53 PL:[53.0, 0.0, 211.4] SR:0 DR:25 LR:-52.99 LO:58.35);ALT=A[chr6:10751363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	10748157	+	chr10	70304647	-	.	111	0	4621447_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4621447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:10748157(+)-10:70304647(+)__10_70290501_70315501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:37 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:111 LR:-326.8 LO:326.8);ALT=A]chr10:70304647];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	13191492	+	chr17	64637274	+	.	37	0	6472096_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6472096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:13191492(+)-17:64637274(-)__17_64631001_64656001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:47 GQ:3.8 PL:[109.4, 0.0, 3.8] SR:0 DR:37 LR:-115.2 LO:115.2);ALT=T[chr17:64637274[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	13305419	+	chr6	13306630	+	.	0	8	2707004_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2707004_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_13303501_13328501_167C;SPAN=1211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:8 DR:0 LR:-1.483 LO:15.0);ALT=T[chr6:13306630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	13321332	+	chr6	13327019	+	AGCACCTTCCATACCAATGCACGGTACATGGACGGGAGAGGGAACCTCTGACTAAAAGTACAAAGTTTCTCAGTAT	0	14	2707061_1	18.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGCACCTTCCATACCAATGCACGGTACATGGACGGGAGAGGGAACCTCTGACTAAAAGTACAAAGTTTCTCAGTAT;MAPQ=60;MATEID=2707061_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_13303501_13328501_213C;SPAN=5687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:14 DR:0 LR:-18.58 LO:29.2);ALT=A[chr6:13327019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	13327168	+	chr6	13328664	+	.	10	0	2707357_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2707357_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:13327168(+)-6:13328664(-)__6_13328001_13353001D;SPAN=1496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:0 DR:10 LR:-18.11 LO:22.2);ALT=G[chr6:13328664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	13579841	+	chr6	13584302	+	.	0	8	2708187_1	0	.	EVDNC=ASSMB;HOMSEQ=CTAAAG;MAPQ=60;MATEID=2708187_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_13573001_13598001_403C;SPAN=4461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:104 GQ:1.5 PL:[0.0, 1.5, 254.1] SR:8 DR:0 LR:1.768 LO:14.56);ALT=G[chr6:13584302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	13618371	+	chr6	13620437	+	.	0	11	2708398_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=2708398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_13597501_13622501_432C;SPAN=2066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:107 GQ:7.4 PL:[7.4, 0.0, 251.6] SR:11 DR:0 LR:-7.322 LO:21.47);ALT=G[chr6:13620437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	13807278	+	chr6	13814247	+	.	0	10	2709171_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2709171_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_13793501_13818501_72C;SPAN=6969;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:10 DR:0 LR:-5.918 LO:19.39);ALT=T[chr6:13814247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	14118296	+	chr6	14131749	+	.	0	7	2710512_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2710512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_14112001_14137001_400C;SPAN=13453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:122 GQ:9.6 PL:[0.0, 9.6, 313.5] SR:7 DR:0 LR:9.946 LO:11.82);ALT=G[chr6:14131749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	19765125	+	chr6	19771185	+	.	115	29	2731437_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGAAAAAAAAACTAACTGG;MAPQ=60;MATEID=2731437_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_19747001_19772001_100C;SECONDARY;SPAN=6060;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:131 DP:4255 GQ:99 PL:[0.0, 719.4, 11770.0] SR:29 DR:115 LR:720.4 LO:185.3);ALT=G[chr6:19771185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	20168872	-	chr6	149031800	+	.	2	4	2732566_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTCTCCTCTCCTCTC;MAPQ=60;MATEID=2732566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_20163501_20188501_104C;SPAN=128862928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:19 GQ:11.3 PL:[11.3, 0.0, 34.4] SR:4 DR:2 LR:-11.36 LO:12.02);ALT=[chr6:149031800[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	20404059	+	chr6	20431339	+	.	8	0	2733324_1	18.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2733324_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:20404059(+)-6:20431339(-)__6_20384001_20409001D;SPAN=27280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=A[chr6:20431339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	27748738	+	chr15	55489062	+	.	61	0	5956060_1	99.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=5956060_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:27748738(+)-15:55489062(-)__15_55468001_55493001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:49 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:61 LR:-178.2 LO:178.2);ALT=C[chr15:55489062[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	28090990	+	chr6	28104522	+	.	22	13	2761215_1	92.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2761215_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_28077001_28102001_280C;SPAN=13532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:62 GQ:56 PL:[92.3, 0.0, 56.0] SR:13 DR:22 LR:-92.54 LO:92.54);ALT=C[chr6:28104522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29034334	+	chr9	109235259	+	.	5	21	2764495_1	56.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=TGTTTCCTGACTTTTTAATGATCGTCATTC;MAPQ=21;MATEID=2764495_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_29032501_29057501_218C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:58 GQ:56.9 PL:[56.9, 0.0, 83.3] SR:21 DR:5 LR:-56.91 LO:57.19);ALT=C[chr9:109235259[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	29643902	+	chr6	29645574	-	.	3	26	2766229_1	79.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGTGTGTGTGTGT;MAPQ=60;MATEID=2766229_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_6_29620501_29645501_186C;SPAN=1672;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:48 GQ:36.5 PL:[79.4, 0.0, 36.5] SR:26 DR:3 LR:-80.26 LO:80.26);ALT=T]chr6:29645574];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	29685488	+	chr6	29688081	+	.	105	24	2766515_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAGAAAGACCCAAGCCT;MAPQ=60;MATEID=2766515_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_29669501_29694501_51C;SPAN=2593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:112 DP:2059 GQ:99 PL:[0.0, 187.7, 5377.0] SR:24 DR:105 LR:188.1 LO:186.4);ALT=T[chr6:29688081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29923065	+	chr6	29766577	+	.	21	0	2766996_1	61.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=2766996_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29766577(-)-6:29923065(+)__6_29914501_29939501D;SPAN=156488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:30 GQ:11.6 PL:[61.1, 0.0, 11.6] SR:0 DR:21 LR:-63.11 LO:63.11);ALT=]chr6:29923065]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	29766711	+	chr6	29923300	+	.	12	0	2766997_1	29.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2766997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29766711(+)-6:29923300(-)__6_29914501_29939501D;SPAN=156589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:0 DR:12 LR:-29.05 LO:29.82);ALT=A[chr6:29923300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29814678	-	chr12	133066751	+	C	4	12	5401471_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=5401471_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_133059501_133084501_306C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:13 DP:10 GQ:3.3 PL:[36.3, 3.3, 0.0] SR:12 DR:4 LR:-36.31 LO:36.31);ALT=[chr12:133066751[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	29814750	+	chr12	133088578	-	.	36	0	5401718_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5401718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29814750(+)-12:133088578(+)__12_133084001_133109001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:22 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=G]chr12:133088578];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	29843498	+	chr6	29849137	+	.	18	0	2767236_1	53.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=2767236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29843498(+)-6:29849137(-)__6_29841001_29866001D;SPAN=5639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:24 GQ:3.5 PL:[53.0, 0.0, 3.5] SR:0 DR:18 LR:-55.19 LO:55.19);ALT=A[chr6:29849137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29843530	+	chr6	29849543	+	.	8	0	2767237_1	14.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2767237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29843530(+)-6:29849543(-)__6_29841001_29866001D;SPAN=6013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:0 DR:8 LR:-14.49 LO:17.76);ALT=T[chr6:29849543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29884497	+	chr6	29970026	+	GGTTTT	2	12	2767193_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GGTTTT;MAPQ=60;MATEID=2767193_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_6_29865501_29890501_263C;SPAN=85529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:45 GQ:34.1 PL:[34.1, 0.0, 73.7] SR:12 DR:2 LR:-34.02 LO:34.88);ALT=G[chr6:29970026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29970132	+	chr6	29884590	+	.	16	0	2767195_1	41.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2767195_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29884590(-)-6:29970132(+)__6_29865501_29890501D;SPAN=85542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:44 GQ:41 PL:[41.0, 0.0, 64.1] SR:0 DR:16 LR:-40.9 LO:41.22);ALT=]chr6:29970132]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	29899782	+	chr6	29901527	+	.	109	86	2767610_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=AAGAATTGAGGAGC;MAPQ=60;MATEID=2767610_2;MATENM=7;NM=1;NUMPARTS=2;SCTG=c_6_29890001_29915001_228C;SPAN=1745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:172 DP:37 GQ:46.3 PL:[508.3, 46.3, 0.0] SR:86 DR:109 LR:-508.3 LO:508.3);ALT=C[chr6:29901527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	29911403	+	chr6	29902295	+	.	15	0	2767618_1	29.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2767618_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:29902295(-)-6:29911403(+)__6_29890001_29915001D;SPAN=9108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:75 GQ:29.3 PL:[29.3, 0.0, 151.4] SR:0 DR:15 LR:-29.2 LO:34.0);ALT=]chr6:29911403]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	30029796	+	chr6	30032450	+	TGACAGGCGCTGCCCTCGATGTGGTCATGAAGGAATGGCATACCACACCAGACAGATGCGTTCAGCCGATGAAGGGCAAACTGTCTTCTACACCTGTACCAACTGCAA	0	36	2767527_1	89.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=TGACAGGCGCTGCCCTCGATGTGGTCATGAAGGAATGGCATACCACACCAGACAGATGCGTTCAGCCGATGAAGGGCAAACTGTCTTCTACACCTGTACCAACTGCAA;MAPQ=60;MATEID=2767527_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_30012501_30037501_253C;SPAN=2654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:110 GQ:89 PL:[89.0, 0.0, 178.1] SR:36 DR:0 LR:-89.04 LO:90.66);ALT=T[chr6:30032450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30035210	+	chr6	30036364	+	.	9	0	2767544_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2767544_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30035210(+)-6:30036364(-)__6_30012501_30037501D;SPAN=1154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:111 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.3636 LO:16.59);ALT=T[chr6:30036364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30262743	+	chr6	30263908	+	.	0	4	2768681_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2768681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30257501_30282501_246C;SPAN=1165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:115 GQ:17.7 PL:[0.0, 17.7, 313.5] SR:4 DR:0 LR:17.95 LO:5.87);ALT=T[chr6:30263908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30436718	-	chr13	48575314	+	.	6	4	5488733_1	9.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=ACCTGAGCAGCAGCCCGC;MAPQ=34;MATEID=5488733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48559001_48584001_159C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:50 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:4 DR:6 LR:-9.561 LO:14.67);ALT=[chr13:48575314[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	30459434	+	chr6	30460524	+	AAAAGGAGGGAGCTACTCTAAGGCTGAGTGGAGCGACAGTGCCCAGGGGTCTGAGTCTCACAGCTTGTAA	6	27	2769602_1	68.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAAAGGAGGGAGCTACTCTAAGGCTGAGTGGAGCGACAGTGCCCAGGGGTCTGAGTCTCACAGCTTGTAA;MAPQ=60;MATEID=2769602_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_30453501_30478501_404C;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:112 GQ:68.9 PL:[68.9, 0.0, 200.9] SR:27 DR:6 LR:-68.69 LO:72.39);ALT=G[chr6:30460524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30539337	+	chr6	30545594	+	ACAAAGTGGTGAAGAAAGGGAAGAAGGACAAGAAGATCAAAAAAAC	6	14	2769509_1	27.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACAAAGTGGTGAAGAAAGGGAAGAAGGACAAGAAGATCAAAAAAAC;MAPQ=57;MATEID=2769509_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_30527001_30552001_62C;SPAN=6257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:106 GQ:27.5 PL:[27.5, 0.0, 228.8] SR:14 DR:6 LR:-27.4 LO:36.71);ALT=G[chr6:30545594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30539337	+	chr6	30545184	+	.	4	8	2769508_1	0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=57;MATEID=2769508_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_30527001_30552001_62C;SPAN=5847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:8 DR:4 LR:5.29 LO:14.13);ALT=G[chr6:30545184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30546355	+	chr6	30547706	+	.	2	10	2769543_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2769543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30527001_30552001_281C;SPAN=1351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:111 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:10 DR:2 LR:-9.539 LO:23.7);ALT=G[chr6:30547706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30585720	+	chr6	30587483	+	.	31	0	2769820_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2769820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30585720(+)-6:30587483(-)__6_30576001_30601001D;SPAN=1763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:108 GQ:73.1 PL:[73.1, 0.0, 188.6] SR:0 DR:31 LR:-73.07 LO:75.91);ALT=G[chr6:30587483[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30585722	+	chr6	30587268	+	.	16	4	2769821_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2769821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30576001_30601001_381C;SPAN=1546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:99 GQ:32.6 PL:[32.6, 0.0, 207.5] SR:4 DR:16 LR:-32.6 LO:39.96);ALT=T[chr6:30587268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30639053	+	chr6	30640410	+	.	0	5	2770065_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=2770065_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30625001_30650001_75C;SPAN=1357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:105 GQ:11.7 PL:[0.0, 11.7, 277.2] SR:5 DR:0 LR:11.94 LO:8.028);ALT=T[chr6:30640410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30645066	+	chr6	30646956	+	.	8	5	2770090_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2770090_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30625001_30650001_378C;SPAN=1890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:102 GQ:12.2 PL:[12.2, 0.0, 233.3] SR:5 DR:8 LR:-11.98 LO:24.17);ALT=C[chr6:30646956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30647169	+	chr6	30652185	+	.	24	29	2770113_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2770113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_30649501_30674501_379C;SPAN=5016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:64 GQ:29 PL:[124.7, 0.0, 29.0] SR:29 DR:24 LR:-127.8 LO:127.8);ALT=G[chr6:30652185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30656753	+	chr6	30658640	+	.	9	0	2770129_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2770129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30656753(+)-6:30658640(-)__6_30649501_30674501D;SPAN=1887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:120 GQ:2.7 PL:[0.0, 2.7, 297.0] SR:0 DR:9 LR:2.802 LO:16.28);ALT=A[chr6:30658640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30688282	+	chr6	30690311	+	.	21	0	2770616_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2770616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30688282(+)-6:30690311(-)__6_30674001_30699001D;SPAN=2029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:175 GQ:22 PL:[22.0, 0.0, 401.6] SR:0 DR:21 LR:-21.91 LO:42.49);ALT=C[chr6:30690311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	30775307	+	chr6	34237082	-	.	8	0	2787433_1	12.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=2787433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:30775307(+)-6:34237082(+)__6_34226501_34251501D;SPAN=3461775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=C]chr6:34237082];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	31211630	+	chr6	31213117	+	.	118	39	2772820_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AATACCCACCACCC;MAPQ=60;MATEID=2772820_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_31188501_31213501_461C;SPAN=1487;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:219 GQ:99 PL:[402.8, 0.0, 128.8] SR:39 DR:118 LR:-410.6 LO:410.6);ALT=C[chr6:31213117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31292074	+	chr6	31294055	+	.	8	0	2774013_1	10.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2774013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31292074(+)-6:31294055(-)__6_31286501_31311501D;SPAN=1981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=G[chr6:31294055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31337861	+	chr6	31341967	+	.	34	34	2773094_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCCA;MAPQ=60;MATEID=2773094_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_31335501_31360501_28C;SPAN=4106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:56 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:34 DR:34 LR:-178.2 LO:178.2);ALT=A[chr6:31341967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31421503	+	chr6	31424387	+	.	24	23	2773396_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TTATAT;MAPQ=60;MATEID=2773396_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_31409001_31434001_331C;SPAN=2884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:23 DR:24 LR:-128.7 LO:128.7);ALT=T[chr6:31424387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31503263	+	chr6	31504277	+	.	6	3	2773720_1	0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2773720_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31482501_31507501_160C;SPAN=1014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:138 GQ:14.1 PL:[0.0, 14.1, 363.0] SR:3 DR:6 LR:14.28 LO:11.44);ALT=C[chr6:31504277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31507053	+	chr6	31508099	+	.	0	23	2773748_1	44.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2773748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31507001_31532001_84C;SPAN=1046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:118 GQ:44 PL:[44.0, 0.0, 242.0] SR:23 DR:0 LR:-43.95 LO:51.84);ALT=T[chr6:31508099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31507096	+	chr6	31509726	+	.	15	0	2773742_1	32.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2773742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31507096(+)-6:31509726(-)__6_31482501_31507501D;SPAN=2630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:0 DR:15 LR:-31.91 LO:35.06);ALT=A[chr6:31509726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31555096	+	chr6	31556294	+	.	127	31	2773950_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2773950_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31531501_31556501_153C;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:148 DP:232 GQ:99 PL:[425.9, 0.0, 135.4] SR:31 DR:127 LR:-433.8 LO:433.8);ALT=G[chr6:31556294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31588636	+	chr6	31590501	+	.	10	6	2774178_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=2774178_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31580501_31605501_80C;SPAN=1865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:102 GQ:18.8 PL:[18.8, 0.0, 226.7] SR:6 DR:10 LR:-18.58 LO:29.2);ALT=G[chr6:31590501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31633966	+	chr6	31636314	+	.	16	0	2774551_1	24.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2774551_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31633966(+)-6:31636314(-)__6_31629501_31654501D;SPAN=2348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:105 GQ:24.5 PL:[24.5, 0.0, 229.1] SR:0 DR:16 LR:-24.37 LO:34.16);ALT=T[chr6:31636314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31633994	+	chr6	31635642	+	.	86	0	2774553_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2774553_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31633994(+)-6:31635642(-)__6_31629501_31654501D;SPAN=1648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:103 GQ:7.8 PL:[264.0, 7.8, 0.0] SR:0 DR:86 LR:-273.4 LO:273.4);ALT=G[chr6:31635642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31635747	+	chr6	31636873	+	ATGAAGAACTGGAAGACAACCCCAACCAGAGTGACCTGATTGAGCAGGCAGCCGAGATGCTTTATGGATTGATCCACGCCCGCTACATCCTTACCAACCGTGGCATCGCCCAGAT	0	71	2774557_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGAAGAACTGGAAGACAACCCCAACCAGAGTGACCTGATTGAGCAGGCAGCCGAGATGCTTTATGGATTGATCCACGCCCGCTACATCCTTACCAACCGTGGCATCGCCCAGAT;MAPQ=60;MATEID=2774557_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_31629501_31654501_37C;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:111 GQ:62.6 PL:[204.5, 0.0, 62.6] SR:71 DR:0 LR:-208.3 LO:208.3);ALT=G[chr6:31636873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31647047	+	chr6	31649005	+	.	0	7	2774605_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=2774605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31629501_31654501_95C;SPAN=1958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:147 GQ:16.6 PL:[0.0, 16.6, 389.4] SR:7 DR:0 LR:16.72 LO:11.24);ALT=T[chr6:31649005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31669118	+	chr6	31670926	+	AGTGCCAGGATGCTGTCAGCATGTTTCTCCAGGGCACGGGGCTGATAGTACGTAT	0	10	2774688_1	1.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AGTGCCAGGATGCTGTCAGCATGTTTCTCCAGGGCACGGGGCTGATAGTACGTAT;MAPQ=60;MATEID=2774688_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_31654001_31679001_82C;SPAN=1808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:116 GQ:1.7 PL:[1.7, 0.0, 278.9] SR:10 DR:0 LR:-1.583 LO:18.71);ALT=C[chr6:31670926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31696763	+	chr6	31697828	+	.	0	4	2774789_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2774789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31678501_31703501_227C;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:115 GQ:17.7 PL:[0.0, 17.7, 313.5] SR:4 DR:0 LR:17.95 LO:5.87);ALT=T[chr6:31697828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31702042	+	chr6	31704038	+	.	166	17	2774836_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2774836_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31678501_31703501_77C;SPAN=1996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:74 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:17 DR:166 LR:-514.9 LO:514.9);ALT=T[chr6:31704038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31745441	+	chr6	31746744	+	.	0	13	2774893_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2774893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31727501_31752501_391C;SPAN=1303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:100 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:13 DR:0 LR:-15.82 LO:26.79);ALT=T[chr6:31746744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31765660	+	chr6	31774532	+	ATGTGAGGGTATTTCTCAGGGTCTGTGACACTGATGTCAGTTAGTTTGATGTTGAGATACTGATCCACAGAATGGAGGGTTCCACAGATGCTCAGGTCATTCTTTAGTTCCACGACCACATCCTTGCCCACAAGGGACTTGAAAAAAGAATAGAAGAG	0	140	2775236_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATGTGAGGGTATTTCTCAGGGTCTGTGACACTGATGTCAGTTAGTTTGATGTTGAGATACTGATCCACAGAATGGAGGGTTCCACAGATGCTCAGGTCATTCTTTAGTTCCACGACCACATCCTTGCCCACAAGGGACTTGAAAAAAGAATAGAAGAG;MAPQ=60;MATEID=2775236_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_31752001_31777001_275C;SPAN=8872;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:131 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:140 DR:0 LR:-415.9 LO:415.9);ALT=C[chr6:31774532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31765887	+	chr6	31774529	+	.	32	0	2775239_1	74.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2775239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31765887(+)-6:31774529(-)__6_31752001_31777001D;SPAN=8642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:115 GQ:74.6 PL:[74.6, 0.0, 203.3] SR:0 DR:32 LR:-74.48 LO:77.84);ALT=T[chr6:31774529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31802978	+	chr6	31804199	+	AGTTGTAAGACGTTCATCGCCGTGTTATCCTTGAGTAA	4	27	2776010_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGTTGTAAGACGTTCATCGCCGTGTTATCCTTGAGTAA;MAPQ=60;MATEID=2776010_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_31801001_31826001_141C;SPAN=1221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:147 GQ:56 PL:[56.0, 0.0, 300.2] SR:27 DR:4 LR:-55.9 LO:65.53);ALT=G[chr6:31804199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31802978	+	chr6	31805011	+	AGTTGTAAGACGTTCATCGCCGTGTTATCCTTGAGTAA	15	42	2776011_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGTTGTAAGACGTTCATCGCCGTGTTATCCTTGAGTAA;MAPQ=60;MATEID=2776011_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_31801001_31826001_108C;SPAN=2033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:144 GQ:99 PL:[129.5, 0.0, 218.6] SR:42 DR:15 LR:-129.3 LO:130.6);ALT=G[chr6:31805011[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31803228	+	chr6	31805011	+	.	3	26	2776014_1	59.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2776014_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_31801001_31826001_108C;SPAN=1783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:136 GQ:59 PL:[59.0, 0.0, 270.2] SR:26 DR:3 LR:-58.88 LO:66.64);ALT=G[chr6:31805011[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31805213	+	chr6	31807319	+	.	9	127	2776030_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2776030_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31801001_31826001_85C;SPAN=2106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:133 DP:203 GQ:99 PL:[384.2, 0.0, 106.9] SR:127 DR:9 LR:-392.6 LO:392.6);ALT=G[chr6:31807319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31920176	+	chr6	31921506	+	.	3	43	2775849_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2775849_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31899001_31924001_394C;SPAN=1330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:124 GQ:99 PL:[111.8, 0.0, 187.7] SR:43 DR:3 LR:-111.7 LO:112.7);ALT=C[chr6:31921506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31923072	+	chr6	31924469	+	.	5	5	2776158_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2776158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31923501_31948501_288C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:5 DR:5 LR:-14.0 LO:19.3);ALT=T[chr6:31924469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31924789	+	chr6	31926149	+	.	2	14	2776165_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2776165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_31923501_31948501_3C;SPAN=1360;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:124 GQ:19.4 PL:[19.4, 0.0, 280.1] SR:14 DR:2 LR:-19.22 LO:32.91);ALT=T[chr6:31926149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	31924828	+	chr6	31926667	+	.	59	0	2776166_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2776166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:31924828(+)-6:31926667(-)__6_31923501_31948501D;SPAN=1839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:102 GQ:78.2 PL:[167.3, 0.0, 78.2] SR:0 DR:59 LR:-168.8 LO:168.8);ALT=G[chr6:31926667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32139284	+	chr6	32143588	+	.	0	11	2776651_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CACCT;MAPQ=60;MATEID=2776651_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32119501_32144501_343C;SPAN=4304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:107 GQ:7.4 PL:[7.4, 0.0, 251.6] SR:11 DR:0 LR:-7.322 LO:21.47);ALT=T[chr6:32143588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32407809	+	chr6	32410223	+	.	162	94	2778079_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2778079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32389001_32414001_126C;SPAN=2414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:223 DP:621 GQ:99 PL:[568.2, 0.0, 937.9] SR:94 DR:162 LR:-567.9 LO:572.9);ALT=G[chr6:32410223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32411243	+	chr6	32412427	+	AGTTTGATGCTCCAAGCCCTCTCCCAGAGACTACAGAGAACGTGGTGTGTGCCCTGGGCCTGACTGTGGGTCTGGTGGGCATCATTATTGGGACCATCTTCATCATCAAGGGATTGCGCAAAAGCAATGCAGCAGAACGCAGGGGGCCTCTGTAAGGCACATGG	0	134	2778103_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGTGA;INSERTION=AGTTTGATGCTCCAAGCCCTCTCCCAGAGACTACAGAGAACGTGGTGTGTGCCCTGGGCCTGACTGTGGGTCTGGTGGGCATCATTATTGGGACCATCTTCATCATCAAGGGATTGCGCAAAAGCAATGCAGCAGAACGCAGGGGGCCTCTGTAAGGCACATGG;MAPQ=60;MATEID=2778103_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32389001_32414001_316C;SPAN=1184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:134 DP:185 GQ:55.6 PL:[392.3, 0.0, 55.6] SR:134 DR:0 LR:-406.6 LO:406.6);ALT=G[chr6:32412427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32459955	+	chr6	32468801	+	.	16	0	2777935_1	46.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=2777935_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32459955(+)-6:32468801(-)__6_32462501_32487501D;SPAN=8846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:9 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:0 DR:16 LR:-46.21 LO:46.21);ALT=A[chr6:32468801[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32541269	+	chr6	32478605	+	.	22	0	2781664_1	61.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2781664_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32478605(-)-6:32541269(+)__6_32536001_32561001D;SPAN=62664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:41 GQ:35.3 PL:[61.7, 0.0, 35.3] SR:0 DR:22 LR:-61.81 LO:61.81);ALT=]chr6:32541269]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32543211	+	chr6	32481164	+	GATTTTAAAACAAACTATTGTACTTGTCAATTGTGGAGT	6	73	2781676_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=GATTTTAAAACAAACTATTGTACTTGTCAATTGTGGAGT;MAPQ=60;MATEID=2781676_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_6_32536001_32561001_358C;SPAN=62047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:68 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:73 DR:6 LR:-224.5 LO:224.5);ALT=]chr6:32543211]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32481243	+	chr6	32543355	+	TCGGCTATTAGA	2	39	2781678_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=TCGGCTATTAGA;MAPQ=60;MATEID=2781678_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_6_32536001_32561001_275C;SPAN=62112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:39 DR:2 LR:-109.9 LO:109.9);ALT=A[chr6:32543355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32481578	+	chr6	32543652	+	GTCACAGCTACGGTTTGGA	8	81	2781683_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=GTCACAGCTACGGTTTGGA;MAPQ=60;MATEID=2781683_2;MATENM=3;NM=2;NUMPARTS=2;SCTG=c_6_32536001_32561001_867C;SPAN=62074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:63 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:81 DR:8 LR:-257.5 LO:257.5);ALT=T[chr6:32543652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32482054	+	chr6	32544150	+	.	16	0	2781687_1	34.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=2781687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32482054(+)-6:32544150(-)__6_32536001_32561001D;SPAN=62096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:67 GQ:34.7 PL:[34.7, 0.0, 127.1] SR:0 DR:16 LR:-34.66 LO:37.67);ALT=C[chr6:32544150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32486443	+	chr6	32489682	+	TCCATTCCACTGTGAGAGGGCTCGTCACGCTTGGGTGCTCCACTTGGCAGGTGTAAACCTCTCCACTTCGAGGAACTGTTTCCAGCATCACCAGGGTCTGGAAGGTCCAGTCTCCATTCTGAATCAGGCCTGTGGACACCACCCCAGCCTTCTCTTCCTGGCTGTTCCGGAACCACCTGACTTCAATGCTGCCTGGATAGAAACCATTCACAGAGCAGACCAGGAGGTTGTGGTGCTGCAGGGTCTGGGTCCTTGCAGGATACACAGTCACCTTAGGCTCAA	0	73	2779864_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TCCATTCCACTGTGAGAGGGCTCGTCACGCTTGGGTGCTCCACTTGGCAGGTGTAAACCTCTCCACTTCGAGGAACTGTTTCCAGCATCACCAGGGTCTGGAAGGTCCAGTCTCCATTCTGAATCAGGCCTGTGGACACCACCCCAGCCTTCTCTTCCTGGCTGTTCCGGAACCACCTGACTTCAATGCTGCCTGGATAGAAACCATTCACAGAGCAGACCAGGAGGTTGTGGTGCTGCAGGGTCTGGGTCCTTGCAGGATACACAGTCACCTTAGGCTCAA;MAPQ=60;MATEID=2779864_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32487001_32512001_788C;SPAN=3239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:86 GQ:9.9 PL:[227.7, 9.9, 0.0] SR:73 DR:0 LR:-233.6 LO:233.6);ALT=C[chr6:32489682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32487430	+	chr6	32489682	+	.	51	30	2779870_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2779870_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32487001_32512001_788C;SPAN=2252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:101 GQ:29 PL:[213.8, 0.0, 29.0] SR:30 DR:51 LR:-221.4 LO:221.4);ALT=T[chr6:32489682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32549610	+	chr6	32489682	+	CTCAA	10	7	2781702_1	21.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=CTCAA;MAPQ=60;MATEID=2781702_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_32536001_32561001_456C;SPAN=59928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:116 GQ:21.5 PL:[21.5, 0.0, 259.1] SR:7 DR:10 LR:-21.39 LO:33.41);ALT=]chr6:32549610]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32489951	+	chr6	32497902	+	.	147	77	2779892_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=2779892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32487001_32512001_80C;SPAN=7951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:175 DP:376 GQ:99 PL:[475.9, 0.0, 436.3] SR:77 DR:147 LR:-475.9 LO:475.9);ALT=G[chr6:32497902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32490844	+	chr6	32526954	+	GCCTCGTGGGTGGCGTTAGGATTTTGGATTTATAGTAAGACAATGGTAAAGTATCGAAGAGTTTAAAGGACAATAAAACCATGATCCCTGTA	11	44	2779904_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;INSERTION=GCCTCGTGGGTGGCGTTAGGATTTTGGATTTATAGTAAGACAATGGTAAAGTATCGAAGAGTTTAAAGGACAATAAAACCATGATCCCTGTA;MAPQ=60;MATEID=2779904_2;MATENM=4;NM=6;NUMPARTS=2;SCTG=c_6_32487001_32512001_803C;SPAN=36110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:29 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:44 DR:11 LR:-158.4 LO:158.4);ALT=A[chr6:32526954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32538527	+	chr6	32494884	+	TGAGCCTG	4	37	2781721_1	99.0	.	DISC_MAPQ=22;EVDNC=TSI_L;INSERTION=TGAGCCTG;MAPQ=60;MATEID=2781721_2;MATENM=5;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_6_32536001_32561001_902C;SPAN=43643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:67 GQ:34.7 PL:[127.1, 0.0, 34.7] SR:37 DR:4 LR:-130.0 LO:130.0);ALT=]chr6:32538527]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32516929	+	chr14	32252018	-	CAGGGCTG	12	62	2778309_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;INSERTION=CAGGGCTG;MAPQ=10;MATEID=2778309_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_32511501_32536501_18C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:34 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:62 DR:12 LR:-201.3 LO:201.3);ALT=A]chr14:32252018];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	32523664	+	chr6	32529893	+	.	11	0	2778369_1	32.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=2778369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32523664(+)-6:32529893(-)__6_32511501_32536501D;SPAN=6229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:16 GQ:5.6 PL:[32.0, 0.0, 5.6] SR:0 DR:11 LR:-32.89 LO:32.89);ALT=A[chr6:32529893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32550879	+	chr6	32524781	+	.	17	0	2781773_1	41.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=2781773_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32524781(-)-6:32550879(+)__6_32536001_32561001D;SPAN=26098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:54 GQ:41.6 PL:[41.6, 0.0, 87.8] SR:0 DR:17 LR:-41.49 LO:42.46);ALT=]chr6:32550879]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32549617	+	chr6	32551886	+	.	30	17	2781935_1	99.0	.	DISC_MAPQ=33;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2781935_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32536001_32561001_813C;SPAN=2269;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:151 GQ:99 PL:[101.3, 0.0, 263.0] SR:17 DR:30 LR:-101.0 LO:105.1);ALT=T[chr6:32551886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32552155	+	chr6	32557420	+	.	162	48	2781961_1	99.0	.	DISC_MAPQ=36;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2781961_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32536001_32561001_813C;SPAN=5265;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:194 DP:324 GQ:99 PL:[552.8, 0.0, 232.6] SR:48 DR:162 LR:-559.7 LO:559.7);ALT=G[chr6:32557420[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32561965	+	chr6	32564609	+	.	88	68	2778886_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ATTATTTTTC;MAPQ=60;MATEID=2778886_2;MATENM=0;NM=12;NUMPARTS=2;SCTG=c_6_32560501_32585501_315C;SPAN=2644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:39 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:68 DR:88 LR:-359.8 LO:359.8);ALT=C[chr6:32564609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32567295	+	chr10	83427201	+	CCACCTGTAATTCCAGCTACGCAGGTGGA	14	90	2778908_1	99.0	.	DISC_MAPQ=47;EVDNC=TSI_L;INSERTION=CCACCTGTAATTCCAGCTACGCAGGTGGA;MAPQ=60;MATEID=2778908_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32560501_32585501_26C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:25 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:90 DR:14 LR:-274.0 LO:274.0);ALT=G[chr10:83427201[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	83427277	+	chr6	32567382	+	CCACCTGTAATTCCAGCTACGCAGGTGGA	10	86	2778915_1	99.0	.	DISC_MAPQ=52;EVDNC=TSI_L;HOMSEQ=CCACTGCACTCCAGCCTGGG;INSERTION=CCACCTGTAATTCCAGCTACGCAGGTGGA;MAPQ=60;MATEID=2778915_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ACAC;SCTG=c_6_32560501_32585501_26C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:26 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:86 DR:10 LR:-254.2 LO:254.2);ALT=]chr10:83427277]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	32605317	+	chr6	32609086	+	.	119	57	2781019_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2781019_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32585001_32610001_973C;SPAN=3769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:183 GQ:13 PL:[468.7, 13.0, 0.0] SR:57 DR:119 LR:-486.7 LO:486.7);ALT=G[chr6:32609086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32608278	+	chr6	32712105	+	AACGGTAAAAGGCTTACACGTCTTGACAGGAATGTCCAGTTCGGCTCATTTGGCTGGAGCCACATTGCAC	7	87	2781056_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CTGCCCATTAGAGGAAAAAG;INSERTION=AACGGTAAAAGGCTTACACGTCTTGACAGGAATGTCCAGTTCGGCTCATTTGGCTGGAGCCACATTGCAC;MAPQ=60;MATEID=2781056_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_32585001_32610001_474C;SPAN=103827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:25 GQ:24 PL:[264.0, 24.0, 0.0] SR:87 DR:7 LR:-264.1 LO:264.1);ALT=G[chr6:32712105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32615820	+	chr6	32718989	+	.	18	0	2780115_1	43.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=2780115_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32615820(+)-6:32718989(-)__6_32707501_32732501D;SPAN=103169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:0 DR:18 LR:-43.7 LO:44.82);ALT=G[chr6:32718989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32719382	+	chr6	32620142	+	.	36	0	2779320_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=2779320_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32620142(-)-6:32719382(+)__6_32609501_32634501D;SPAN=99240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:7 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=]chr6:32719382]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32623469	+	chr6	32722262	+	.	12	0	2779360_1	28.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=2779360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32623469(+)-6:32722262(-)__6_32609501_32634501D;SPAN=98793;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:41 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:0 DR:12 LR:-28.5 LO:29.51);ALT=C[chr6:32722262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32623587	+	chr6	32624623	+	.	31	0	2779362_1	89.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=2779362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32623587(+)-6:32624623(-)__6_32609501_32634501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:5 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=C[chr6:32624623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32626583	+	chr6	32722802	+	.	2	53	2779369_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ACTGTGAGGA;MAPQ=60;MATEID=2779369_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_32609501_32634501_83C;SPAN=96219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:53 DR:2 LR:-158.4 LO:158.4);ALT=A[chr6:32722802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32628028	+	chr6	32629130	+	TTCC	6	14	2779395_1	29.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TTCC;MAPQ=60;MATEID=2779395_2;MATENM=1;NM=5;NUMPARTS=2;SCTG=c_6_32609501_32634501_681C;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:122 GQ:29.9 PL:[29.9, 0.0, 264.2] SR:14 DR:6 LR:-29.67 LO:40.77);ALT=T[chr6:32629130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32628028	+	chr6	32629743	+	TTCTGACTCCTTTGACGGATGATAAGGCCCAGCCCAAGGAAGATCAGCCCCAGCACGAAGCCTCCAACGCCACTCAGCATCTTGCTCTGGGCAGATTCAGACTGAGCC	10	24	2779396_1	74.0	.	DISC_MAPQ=49;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTCTGACTCCTTTGACGGATGATAAGGCCCAGCCCAAGGAAGATCAGCCCCAGCACGAAGCCTCCAACGCCACTCAGCATCTTGCTCTGGGCAGATTCAGACTGAGCC;MAPQ=60;MATEID=2779396_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32609501_32634501_471C;SPAN=1715;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:115 GQ:74.6 PL:[74.6, 0.0, 203.3] SR:24 DR:10 LR:-74.48 LO:77.84);ALT=T[chr6:32629743[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32630027	+	chr6	32632575	+	.	29	12	2779412_1	98.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2779412_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32609501_32634501_416C;SPAN=2548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:62 GQ:49.4 PL:[98.9, 0.0, 49.4] SR:12 DR:29 LR:-99.53 LO:99.53);ALT=T[chr6:32632575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32630915	+	chr6	32727766	+	TCCACCTGAAATC	2	16	2779433_1	37.0	.	DISC_MAPQ=42;EVDNC=ASDIS;INSERTION=TCCACCTGAAATC;MAPQ=60;MATEID=2779433_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_6_32609501_32634501_439C;SPAN=96851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:83 GQ:37.1 PL:[37.1, 0.0, 162.5] SR:16 DR:2 LR:-36.93 LO:41.51);ALT=G[chr6:32727766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32728042	+	chr6	32631211	+	TGGAAAACAC	30	15	2779438_1	99.0	.	DISC_MAPQ=44;EVDNC=TSI_L;INSERTION=TGGAAAACAC;MAPQ=60;MATEID=2779438_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACA;SCTG=c_6_32609501_32634501_307C;SPAN=96831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:24 GQ:12 PL:[132.0, 12.0, 0.0] SR:15 DR:30 LR:-132.0 LO:132.0);ALT=]chr6:32728042]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32631611	+	chr6	32728417	+	.	2	33	2779446_1	99.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CCAAAAGCAACCTGAAACTATTTTTATCCAATAATTTAAT;MAPQ=60;MATEID=2779446_2;MATENM=5;NM=7;NUMPARTS=2;SCTG=c_6_32609501_32634501_510C;SPAN=96806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:42 GQ:4.5 PL:[108.9, 4.5, 0.0] SR:33 DR:2 LR:-111.2 LO:111.2);ALT=T[chr6:32728417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32632845	+	chr6	32634276	+	.	122	15	2778436_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=43;MATEID=2778436_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32634001_32659001_128C;SPAN=1431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:107 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:15 DR:122 LR:-402.7 LO:402.7);ALT=C[chr6:32634276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32778699	+	chr6	32779819	+	.	87	0	2780350_1	99.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=2780350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32778699(+)-6:32779819(-)__6_32756501_32781501D;SPAN=1120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:28 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:0 DR:87 LR:-257.5 LO:257.5);ALT=C[chr6:32779819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32778708	+	chr6	32853320	+	.	30	29	2780713_1	99.0	.	DISC_MAPQ=51;EVDNC=TSI_L;HOMSEQ=TTCTCCTGCCTCAGCCTCCGGAGTAGCTGGGACTACAGGCGC;MAPQ=24;MATEID=2780713_2;MATENM=2;NM=5;NUMPARTS=3;REPSEQ=CGCG;SCTG=c_6_32830001_32855001_450C;SPAN=74612;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:74 GQ:32.9 PL:[145.1, 0.0, 32.9] SR:29 DR:30 LR:-148.8 LO:148.8);ALT=C[chr6:32853320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32853410	+	chr6	32779821	+	.	0	80	2780355_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=2780355_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_32756501_32781501_22C;SPAN=73589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:21 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:80 DR:0 LR:-237.7 LO:237.7);ALT=]chr6:32853410]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	32810560	+	chr6	32811627	+	TAATGTAGGACCCAGCTGAGGCCCGAGAATCCACTGCTGCAATCACTCCATGCTGGAACTTGAAGGCGAGCGTGGTGGTGCCATGGGCCATCTCAATCTGAACGTTCCTTTCTCCGTCCCCACCCAGGGACTGGAAGAATTCTGTGGG	0	134	2780544_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TAATGTAGGACCCAGCTGAGGCCCGAGAATCCACTGCTGCAATCACTCCATGCTGGAACTTGAAGGCGAGCGTGGTGGTGCCATGGGCCATCTCAATCTGAACGTTCCTTTCTCCGTCCCCACCCAGGGACTGGAAGAATTCTGTGGG;MAPQ=60;MATEID=2780544_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32805501_32830501_177C;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:141 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:134 DR:0 LR:-415.9 LO:415.9);ALT=C[chr6:32811627[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32810905	+	chr6	32812066	+	.	9	0	2780549_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2780549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32810905(+)-6:32812066(-)__6_32805501_32830501D;SPAN=1161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:110 GQ:0 PL:[0.0, 0.0, 267.3] SR:0 DR:9 LR:0.0927 LO:16.63);ALT=T[chr6:32812066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32822052	+	chr6	32825780	+	.	8	0	2780591_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2780591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:32822052(+)-6:32825780(-)__6_32805501_32830501D;SPAN=3728;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:108 GQ:2.7 PL:[0.0, 2.7, 267.3] SR:0 DR:8 LR:2.852 LO:14.42);ALT=G[chr6:32825780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32822066	+	chr6	32823914	+	.	27	18	2780592_1	63.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2780592_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCACCA;SCTG=c_6_32805501_32830501_416C;SPAN=1848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:103 GQ:63.4 PL:[63.4, 0.0, 120.6] SR:18 DR:27 LR:-63.17 LO:64.41);ALT=G[chr6:32823914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32822066	+	chr6	32825039	+	ACCACCATCATGGCAGTGGAGTTTGACGGGGGCGTTGTGATGGGTTCTGATTCCCGAGTGTCTGCAG	90	93	2780593_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACCACCATCATGGCAGTGGAGTTTGACGGGGGCGTTGTGATGGGTTCTGATTCCCGAGTGTCTGCAG;MAPQ=60;MATEID=2780593_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_32805501_32830501_416C;SPAN=2973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:124 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:93 DR:90 LR:-435.7 LO:435.7);ALT=G[chr6:32825039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32862704	+	chr6	32868696	+	.	6	4	2780470_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2780470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32854501_32879501_115C;SPAN=5992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:4 DR:6 LR:-1.483 LO:15.0);ALT=G[chr6:32868696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32906744	+	chr6	32908528	+	.	22	40	2781104_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=2781104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32903501_32928501_359C;SPAN=1784;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:117 GQ:99 PL:[123.5, 0.0, 159.8] SR:40 DR:22 LR:-123.4 LO:123.7);ALT=T[chr6:32908528[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32918582	+	chr6	32920726	+	.	151	38	2781158_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2781158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_32903501_32928501_173C;SPAN=2144;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:164 DP:166 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:38 DR:151 LR:-491.8 LO:491.8);ALT=T[chr6:32920726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	32946166	+	chr6	32947605	+	.	6	3	2781281_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2781281_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_32928001_32953001_94C;SPAN=1439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:124 GQ:6.9 PL:[0.0, 6.9, 313.5] SR:3 DR:6 LR:7.187 LO:13.93);ALT=G[chr6:32947605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33026728	+	chr6	33028601	+	.	15	22	2782381_1	88.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2782381_2;MATENM=10;NM=4;NUMPARTS=2;REPSEQ=TTTTTT;SCTG=c_6_33026001_33051001_186C;SECONDARY;SPAN=1873;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:45 GQ:4.1 PL:[88.4, 4.1, 0.0] SR:22 DR:15 LR:-91.07 LO:91.07);ALT=T[chr6:33028601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33033126	+	chr6	33036412	+	.	18	59	2782422_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=2782422_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_344C;SPAN=3286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:192 GQ:99 PL:[169.4, 0.0, 294.8] SR:59 DR:18 LR:-169.2 LO:171.1);ALT=T[chr6:33036412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33037664	+	chr6	33041248	+	.	183	104	2782450_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2782450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_199C;SPAN=3584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:238 DP:410 GQ:99 PL:[674.5, 0.0, 321.4] SR:104 DR:183 LR:-681.4 LO:681.4);ALT=C[chr6:33041248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33043918	+	chr6	33048455	+	AGAATG	175	163	2782470_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=AGAATG;MAPQ=60;MATEID=2782470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_206C;SPAN=4537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:302 DP:539 GQ:99 PL:[850.9, 0.0, 458.1] SR:163 DR:175 LR:-857.2 LO:857.2);ALT=G[chr6:33048455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33048712	+	chr6	33052725	+	.	7	7	2782492_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2782492_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33026001_33051001_407C;SPAN=4013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:7 DR:7 LR:-28.06 LO:32.03);ALT=G[chr6:33052725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33269550	+	chr6	33271905	+	TCTTTGAATCCTTGCAGGTGGACAGGTAGACAG	0	11	2783190_1	20.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCTTTGAATCCTTGCAGGTGGACAGGTAGACAG;MAPQ=60;MATEID=2783190_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_33271001_33296001_205C;SPAN=2355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:60 GQ:20 PL:[20.0, 0.0, 125.6] SR:11 DR:0 LR:-20.06 LO:24.46);ALT=T[chr6:33271905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33273167	+	chr6	33280994	+	.	5	3	2783202_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=2783202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33271001_33296001_174C;SPAN=7827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:113 GQ:7.2 PL:[0.0, 7.2, 287.1] SR:3 DR:5 LR:7.508 LO:12.06);ALT=G[chr6:33280994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33583198	+	chr6	33585845	+	.	24	36	2784716_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2784716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33565001_33590001_160C;SPAN=2647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:60 GQ:0.2 PL:[145.4, 0.0, 0.2] SR:36 DR:24 LR:-154.5 LO:154.5);ALT=C[chr6:33585845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33665530	+	chr6	33669123	+	TGGACAGGATCAGCTTGTACTCTTCCAACGACAGGCCACTGAAGCTGGTGTCTCTGGGGCGAGGGTA	0	95	2785188_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGGACAGGATCAGCTTGTACTCTTCCAACGACAGGCCACTGAAGCTGGTGTCTCTGGGGCGAGGGTA;MAPQ=60;MATEID=2785188_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_33663001_33688001_53C;SPAN=3593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:95 DP:126 GQ:25.4 PL:[279.5, 0.0, 25.4] SR:95 DR:0 LR:-291.7 LO:291.7);ALT=G[chr6:33669123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33665576	+	chr6	33679323	+	.	10	0	2785189_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2785189_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:33665576(+)-6:33679323(-)__6_33663001_33688001D;SPAN=13747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:105 GQ:4.7 PL:[4.7, 0.0, 248.9] SR:0 DR:10 LR:-4.563 LO:19.17);ALT=G[chr6:33679323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33668339	+	chr6	33679412	+	.	19	0	2785201_1	30.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2785201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:33668339(+)-6:33679412(-)__6_33663001_33688001D;SPAN=11073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:119 GQ:30.5 PL:[30.5, 0.0, 258.2] SR:0 DR:19 LR:-30.48 LO:40.99);ALT=A[chr6:33679412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33669200	+	chr6	33679324	+	.	0	47	2785205_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=2785205_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33663001_33688001_449C;SPAN=10124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:132 GQ:99 PL:[119.6, 0.0, 198.8] SR:47 DR:0 LR:-119.4 LO:120.5);ALT=G[chr6:33679324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	33937829	+	chr6	33942698	+	GCTTTTAT	0	25	2785889_1	64.0	.	EVDNC=ASSMB;INSERTION=GCTTTTAT;MAPQ=60;MATEID=2785889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_33932501_33957501_29C;SPAN=4869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:68 GQ:64.1 PL:[64.1, 0.0, 100.4] SR:25 DR:0 LR:-64.1 LO:64.55);ALT=A[chr6:33942698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34205094	+	chr6	34208513	+	.	119	104	2787700_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=2787700_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GCGC;SCTG=c_6_34202001_34227001_392C;SPAN=3419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:188 DP:119 GQ:50.8 PL:[557.8, 50.8, 0.0] SR:104 DR:119 LR:-557.8 LO:557.8);ALT=G[chr6:34208513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34214987	+	chr6	34216754	+	.	8	0	2787753_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2787753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:34214987(+)-6:34216754(-)__6_34202001_34227001D;SPAN=1767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=C[chr6:34216754[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34215649	+	chr6	34216754	+	.	19	0	2787759_1	33.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2787759_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:34215649(+)-6:34216754(-)__6_34202001_34227001D;SPAN=1105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:108 GQ:33.5 PL:[33.5, 0.0, 228.2] SR:0 DR:19 LR:-33.46 LO:41.88);ALT=G[chr6:34216754[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34309751	+	chr6	34360038	+	.	10	18	2787814_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=2787814_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_34349001_34374001_369C;SPAN=50287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:51 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:18 DR:10 LR:-68.79 LO:68.79);ALT=T[chr6:34360038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34725363	+	chr6	34735684	+	.	8	0	2789428_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=2789428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:34725363(+)-6:34735684(-)__6_34716501_34741501D;SPAN=10321;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=G[chr6:34735684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34725374	+	chr6	34730371	+	.	10	0	2789430_1	1.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=2789430_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:34725374(+)-6:34730371(-)__6_34716501_34741501D;SPAN=4997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:116 GQ:1.7 PL:[1.7, 0.0, 278.9] SR:0 DR:10 LR:-1.583 LO:18.71);ALT=T[chr6:34730371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	34850859	+	chr6	34855564	+	.	0	14	2790166_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2790166_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_34839001_34864001_193C;SPAN=4705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:101 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:14 DR:0 LR:-18.85 LO:29.27);ALT=T[chr6:34855564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35265732	+	chr6	35277445	+	.	50	10	2791568_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=2791568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35255501_35280501_285C;SPAN=11713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:101 GQ:91.7 PL:[151.1, 0.0, 91.7] SR:10 DR:50 LR:-151.6 LO:151.6);ALT=G[chr6:35277445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35604937	+	chr6	35610497	+	.	0	7	2793298_1	19.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=2793298_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_35647501_35672501_260C;SPAN=5560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:7 DP:0 GQ:1.8 PL:[19.8, 1.8, 0.0] SR:7 DR:0 LR:-19.8 LO:19.8);ALT=T[chr6:35610497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35610623	+	chr6	35656579	+	.	8	4	2793301_1	12.0	.	DISC_MAPQ=51;EVDNC=TSI_L;HOMSEQ=ACCTG;MAPQ=60;MATEID=2793301_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CGCCGC;SCTG=c_6_35647501_35672501_260C;SPAN=45956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:12.8 PL:[12.8, 0.0, 75.2] SR:4 DR:8 LR:-12.75 LO:15.79);ALT=G[chr6:35656579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35626434	+	chr6	35629745	+	.	83	77	2793238_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=2793238_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35623001_35648001_95C;SPAN=3311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:38 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:77 DR:83 LR:-406.0 LO:406.0);ALT=G[chr6:35629745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35766788	+	chr6	35754561	+	.	96	58	2794250_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAC;MAPQ=60;MATEID=2794250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35745501_35770501_86C;SPAN=12227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:130 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:58 DR:96 LR:-386.2 LO:386.2);ALT=]chr6:35766788]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	35840505	+	chr6	35842008	+	.	0	19	2793689_1	35.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=2793689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35819001_35844001_295C;SPAN=1503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:102 GQ:35.3 PL:[35.3, 0.0, 210.2] SR:19 DR:0 LR:-35.09 LO:42.4);ALT=C[chr6:35842008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35856702	+	chr6	35858671	+	.	0	16	2794010_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=2794010_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35843501_35868501_218C;SPAN=1969;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:98 GQ:26.3 PL:[26.3, 0.0, 211.1] SR:16 DR:0 LR:-26.27 LO:34.69);ALT=T[chr6:35858671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35856723	+	chr6	35888259	+	.	8	0	2794355_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2794355_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:35856723(+)-6:35888259(-)__6_35868001_35893001D;SPAN=31536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=A[chr6:35888259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35858790	+	chr6	35888245	+	.	4	5	2794357_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2794357_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_35868001_35893001_319C;SPAN=29455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:5 DR:4 LR:-19.14 LO:21.04);ALT=T[chr6:35888245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	35858834	+	chr6	35888820	+	.	13	0	2794358_1	29.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2794358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:35858834(+)-6:35888820(-)__6_35868001_35893001D;SPAN=29986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:50 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:0 DR:13 LR:-29.37 LO:31.17);ALT=A[chr6:35888820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36410900	+	chr6	36437828	+	.	8	0	2796261_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2796261_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:36410900(+)-6:36437828(-)__6_36431501_36456501D;SPAN=26928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:0 DR:8 LR:-10.69 LO:16.71);ALT=C[chr6:36437828[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36507982	+	chr6	36514967	+	.	0	13	2796605_1	13.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2796605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36505001_36530001_355C;SPAN=6985;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:111 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:13 DR:0 LR:-12.84 LO:26.15);ALT=C[chr6:36514967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36562258	+	chr6	36564537	+	.	131	25	2797146_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2797146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36554001_36579001_207C;SPAN=2279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:135 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:25 DR:131 LR:-448.9 LO:448.9);ALT=G[chr6:36564537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36564745	+	chr6	36566624	+	.	4	22	2797160_1	47.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=14;MATEID=2797160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36554001_36579001_465C;SPAN=1879;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:116 GQ:47.9 PL:[47.9, 0.0, 232.7] SR:22 DR:4 LR:-47.8 LO:54.79);ALT=G[chr6:36566624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36646576	+	chr6	36651872	+	.	29	2	2797320_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2797320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36652001_36677001_6C;SPAN=5296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:0 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:2 DR:29 LR:-89.12 LO:89.12);ALT=G[chr6:36651872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36839634	+	chr6	36842508	+	.	8	0	2798044_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2798044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:36839634(+)-6:36842508(-)__6_36823501_36848501D;SPAN=2874;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:111 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.665 LO:14.32);ALT=A[chr6:36842508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36853846	+	chr6	36867207	+	.	12	0	2798290_1	6.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2798290_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:36853846(+)-6:36867207(-)__6_36848001_36873001D;SPAN=13361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:124 GQ:6.2 PL:[6.2, 0.0, 293.3] SR:0 DR:12 LR:-6.017 LO:23.09);ALT=C[chr6:36867207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36946388	+	chr6	36949364	+	.	0	10	2798644_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=2798644_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36946001_36971001_173C;SPAN=2976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:123 GQ:0 PL:[0.0, 0.0, 297.0] SR:10 DR:0 LR:0.3137 LO:18.45);ALT=C[chr6:36949364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	36949450	+	chr6	36953624	+	.	0	25	2798658_1	51.0	.	EVDNC=ASSMB;HOMSEQ=CCCACCT;MAPQ=60;MATEID=2798658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_36946001_36971001_53C;SPAN=4174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:115 GQ:51.5 PL:[51.5, 0.0, 226.4] SR:25 DR:0 LR:-51.37 LO:57.69);ALT=T[chr6:36953624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37225750	+	chr6	37231403	+	.	18	16	2799650_1	49.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2799650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_37215501_37240501_225C;SPAN=5653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:136 GQ:49.1 PL:[49.1, 0.0, 280.1] SR:16 DR:18 LR:-48.98 LO:58.35);ALT=G[chr6:37231403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37451066	+	chr6	37452875	+	GTAGTTGGAGGCTTTGTTCATTAGGCTGTTTTTCTCCTTCTCCAGGGACCT	0	52	2800674_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=GTAGTTGGAGGCTTTGTTCATTAGGCTGTTTTTCTCCTTCTCCAGGGACCT;MAPQ=60;MATEID=2800674_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_6_37436001_37461001_262C;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:113 GQ:99 PL:[141.2, 0.0, 131.3] SR:52 DR:0 LR:-141.0 LO:141.0);ALT=C[chr6:37452875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37451113	+	chr6	37467595	+	.	31	0	2800705_1	83.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2800705_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:37451113(+)-6:37467595(-)__6_37460501_37485501D;SPAN=16482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:68 GQ:80.6 PL:[83.9, 0.0, 80.6] SR:0 DR:31 LR:-83.91 LO:83.91);ALT=T[chr6:37467595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	37452972	+	chr6	37467598	+	.	48	8	2800707_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2800707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_37460501_37485501_440C;SPAN=14626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:72 GQ:33.5 PL:[139.1, 0.0, 33.5] SR:8 DR:48 LR:-142.3 LO:142.3);ALT=T[chr6:37467598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	38254865	-	chr8	15474649	+	.	3	14	3757909_1	44.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTT;MAPQ=60;MATEID=3757909_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_15459501_15484501_146C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:32 GQ:31.1 PL:[44.3, 0.0, 31.1] SR:14 DR:3 LR:-44.22 LO:44.22);ALT=[chr8:15474649[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	38652336	+	chr6	38670799	+	.	16	0	2805126_1	35.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2805126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:38652336(+)-6:38670799(-)__6_38661001_38686001D;SPAN=18463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:63 GQ:35.9 PL:[35.9, 0.0, 115.1] SR:0 DR:16 LR:-35.75 LO:38.17);ALT=G[chr6:38670799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	38654800	+	chr6	38670799	+	.	23	0	2805128_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2805128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:38654800(+)-6:38670799(-)__6_38661001_38686001D;SPAN=15999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:63 GQ:59 PL:[59.0, 0.0, 92.0] SR:0 DR:23 LR:-58.86 LO:59.3);ALT=C[chr6:38670799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41250482	+	chr6	41254356	+	.	21	0	2813153_1	40.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=2813153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:41250482(+)-6:41254356(-)__6_41233501_41258501D;SPAN=3874;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:108 GQ:40.1 PL:[40.1, 0.0, 221.6] SR:0 DR:21 LR:-40.06 LO:47.3);ALT=T[chr6:41254356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41658979	+	chr6	41691212	+	.	8	0	2814875_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2814875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:41658979(+)-6:41691212(-)__6_41674501_41699501D;SPAN=32233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=G[chr6:41691212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41755564	+	chr6	41756968	+	.	52	112	2814998_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2814998_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_41748001_41773001_83C;SPAN=1404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:119 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:112 DR:52 LR:-422.5 LO:422.5);ALT=G[chr6:41756968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	41755578	+	chr12	125541044	-	.	37	0	2814999_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2814999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:41755578(+)-12:125541044(+)__6_41748001_41773001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:28 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:0 DR:37 LR:-108.9 LO:108.9);ALT=G]chr12:125541044];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	41782965	-	chr6	41784616	+	.	9	0	2815111_1	3.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2815111_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:41782965(-)-6:41784616(-)__6_41772501_41797501D;SPAN=1651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:0 DR:9 LR:-3.429 LO:17.14);ALT=[chr6:41784616[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	42019251	+	chr6	42023269	+	.	0	7	2816142_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2816142_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_42017501_42042501_136C;SPAN=4018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:7 DR:0 LR:2.902 LO:12.57);ALT=T[chr6:42023269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42179696	+	chr6	42185536	+	.	13	0	2817184_1	15.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=2817184_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:42179696(+)-6:42185536(-)__6_42164501_42189501D;SPAN=5840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:101 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:0 DR:13 LR:-15.55 LO:26.73);ALT=T[chr6:42185536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42532135	+	chr6	42541471	+	.	11	11	2818357_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2818357_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42532001_42557001_87C;SPAN=9336;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:136 GQ:12.8 PL:[12.8, 0.0, 316.4] SR:11 DR:11 LR:-12.67 LO:29.76);ALT=G[chr6:42541471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42897459	+	chr6	42902211	+	.	0	72	2820435_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2820435_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42875001_42900001_395C;SPAN=4752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:76 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:72 DR:0 LR:-224.5 LO:224.5);ALT=G[chr6:42902211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42897460	+	chr6	42903310	+	.	11	8	2820437_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2820437_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42875001_42900001_325C;SPAN=5850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:74 GQ:29.6 PL:[29.6, 0.0, 148.4] SR:8 DR:11 LR:-29.47 LO:34.09);ALT=G[chr6:42903310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42903409	+	chr6	42905453	+	.	3	9	2820002_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2820002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42899501_42924501_341C;SPAN=2044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:110 GQ:3.2 PL:[3.2, 0.0, 263.9] SR:9 DR:3 LR:-3.208 LO:18.96);ALT=G[chr6:42905453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42952443	+	chr6	42957347	+	.	2	2	2820152_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2820152_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42948501_42973501_242C;SPAN=4904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:123 GQ:19.8 PL:[0.0, 19.8, 336.6] SR:2 DR:2 LR:20.12 LO:5.753);ALT=G[chr6:42957347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42982079	+	chr6	42985253	+	.	8	0	2820259_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2820259_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:42982079(+)-6:42985253(-)__6_42973001_42998001D;SPAN=3174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=C[chr6:42985253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	42982086	+	chr6	42984868	+	.	19	3	2820260_1	42.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GCAG;MAPQ=60;MATEID=2820260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_42973001_42998001_295C;SPAN=2782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:99 GQ:42.5 PL:[42.5, 0.0, 197.6] SR:3 DR:19 LR:-42.5 LO:48.2);ALT=G[chr6:42984868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	43025973	+	chr6	43027024	+	.	39	12	2820592_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2820592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_43022001_43047001_309C;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:108 GQ:99 PL:[119.3, 0.0, 142.4] SR:12 DR:39 LR:-119.3 LO:119.4);ALT=T[chr6:43027024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	43193931	+	chr6	43197049	+	.	17	0	2821444_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2821444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:43193931(+)-6:43197049(-)__6_43193501_43218501D;SPAN=3118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:126 GQ:22.1 PL:[22.1, 0.0, 282.8] SR:0 DR:17 LR:-21.98 LO:35.32);ALT=C[chr6:43197049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	43194183	+	chr6	43197134	+	.	30	0	2821448_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2821448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:43194183(+)-6:43197134(-)__6_43193501_43218501D;SPAN=2951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:114 GQ:68.3 PL:[68.3, 0.0, 206.9] SR:0 DR:30 LR:-68.15 LO:72.11);ALT=T[chr6:43197134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	43646389	+	chr6	43655460	+	.	9	0	2822753_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=2822753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:43646389(+)-6:43655460(-)__6_43634501_43659501D;SPAN=9071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:0 DR:9 LR:-0.7201 LO:16.74);ALT=G[chr6:43655460[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44081949	+	chr6	44084278	+	.	0	23	2824766_1	46.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=2824766_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44075501_44100501_221C;SPAN=2329;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:108 GQ:46.7 PL:[46.7, 0.0, 215.0] SR:23 DR:0 LR:-46.66 LO:52.84);ALT=G[chr6:44084278[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44081993	+	chr6	44095079	+	.	37	0	2824769_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2824769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44081993(+)-6:44095079(-)__6_44075501_44100501D;SPAN=13086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:136 GQ:85.4 PL:[85.4, 0.0, 243.8] SR:0 DR:37 LR:-85.29 LO:89.57);ALT=C[chr6:44095079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44084367	+	chr6	44095080	+	.	12	5	2824776_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2824776_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44075501_44100501_231C;SPAN=10713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:121 GQ:10.4 PL:[10.4, 0.0, 281.0] SR:5 DR:12 LR:-10.13 LO:25.64);ALT=C[chr6:44095080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44214926	+	chr6	44217111	+	.	34	0	2825377_1	76.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2825377_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44214926(+)-6:44217111(-)__6_44198001_44223001D;SPAN=2185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:134 GQ:76.1 PL:[76.1, 0.0, 247.7] SR:0 DR:34 LR:-75.93 LO:81.1);ALT=T[chr6:44217111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44214931	+	chr6	44216351	+	.	72	0	2825378_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2825378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:44214931(+)-6:44216351(-)__6_44198001_44223001D;SPAN=1420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:115 GQ:71.3 PL:[206.6, 0.0, 71.3] SR:0 DR:72 LR:-210.0 LO:210.0);ALT=A[chr6:44216351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44355606	+	chr6	44358003	+	.	10	11	2825748_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2825748_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44345001_44370001_19C;SPAN=2397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:108 GQ:20.3 PL:[20.3, 0.0, 241.4] SR:11 DR:10 LR:-20.26 LO:31.37);ALT=G[chr6:44358003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44364177	+	chr6	44371544	+	.	2	4	2825779_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2825779_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44345001_44370001_204C;SPAN=7367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:52 GQ:2.6 PL:[2.6, 0.0, 121.4] SR:4 DR:2 LR:-2.417 LO:9.606);ALT=G[chr6:44371544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	44394462	+	chr6	44397448	+	.	2	3	2825984_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2825984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_44394001_44419001_341C;SPAN=2986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:92 GQ:11.4 PL:[0.0, 11.4, 244.2] SR:3 DR:2 LR:11.72 LO:6.262);ALT=G[chr6:44397448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	45390696	+	chr6	45405682	+	GGTAGCCCTCGGAGAGGTACCAGATGGGACTGTGGTTACTGTCATGGCGGGTAACGATGAAAATTATTCTGCTGAGCTCCGGAATGCCTCTGCTGTTATGAAAAACCAAGTAGCAAGGTTCAACGATCTGAGATTTGTGGGCCGGAGTGGACG	4	11	2829402_1	33.0	.	DISC_MAPQ=52;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=GGTAGCCCTCGGAGAGGTACCAGATGGGACTGTGGTTACTGTCATGGCGGGTAACGATGAAAATTATTCTGCTGAGCTCCGGAATGCCTCTGCTGTTATGAAAAACCAAGTAGCAAGGTTCAACGATCTGAGATTTGTGGGCCGGAGTGGACG;MAPQ=60;MATEID=2829402_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_45374001_45399001_275C;SPAN=14986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:47 GQ:33.5 PL:[33.5, 0.0, 79.7] SR:11 DR:4 LR:-33.48 LO:34.55);ALT=T[chr6:45405682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	45390696	+	chr6	45399598	+	.	7	9	2829401_1	33.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=2829401_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_45374001_45399001_275C;SPAN=8902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:47 GQ:33.5 PL:[33.5, 0.0, 79.7] SR:9 DR:7 LR:-33.48 LO:34.55);ALT=T[chr6:45399598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	51847696	+	chr6	101194037	+	AAAAAAAA	7	13	2960137_1	56.0	.	DISC_MAPQ=26;EVDNC=ASDIS;INSERTION=AAAAAAAA;MAPQ=0;MATEID=2960137_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_101185001_101210001_53C;SPAN=49346341;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:13 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:13 DR:7 LR:-56.11 LO:56.11);ALT=A[chr6:101194037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52129587	+	chr6	52131409	+	GATTCACTCAACTCCACTTTCTGGGATTCCTTGGTCTCCTGTGAGTCTGCCGTCTTTGGAGTGTGTA	0	9	2849796_1	0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTT;INSERTION=GATTCACTCAACTCCACTTTCTGGGATTCCTTGGTCTCCTGTGAGTCTGCCGTCTTTGGAGTGTGTA;MAPQ=60;MATEID=2849796_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_52111501_52136501_30C;SPAN=1822;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:9 DR:0 LR:-0.7201 LO:16.74);ALT=G[chr6:52131409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52148206	+	chr6	52149394	+	.	12	4	2849564_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2849564_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_52136001_52161001_316C;SPAN=1188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:147 GQ:0 PL:[0.0, 0.0, 356.4] SR:4 DR:12 LR:0.2139 LO:22.16);ALT=T[chr6:52149394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52285271	+	chr6	52288743	+	.	22	17	2850121_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=2850121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_52283001_52308001_327C;SPAN=3472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:120 GQ:63.2 PL:[63.2, 0.0, 228.2] SR:17 DR:22 LR:-63.22 LO:68.45);ALT=G[chr6:52288743[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52536043	+	chr6	52541883	+	.	16	10	2851022_1	40.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=2851022_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_52528001_52553001_264C;SPAN=5840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:119 GQ:40.4 PL:[40.4, 0.0, 248.3] SR:10 DR:16 LR:-40.38 LO:49.02);ALT=G[chr6:52541883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52536094	+	chr6	52546607	+	.	23	0	2851026_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2851026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:52536094(+)-6:52546607(-)__6_52528001_52553001D;SPAN=10513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:106 GQ:47.3 PL:[47.3, 0.0, 209.0] SR:0 DR:23 LR:-47.21 LO:53.05);ALT=A[chr6:52546607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52546712	+	chr6	52548876	+	.	0	10	2851071_1	3.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2851071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_52528001_52553001_354C;SPAN=2164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:111 GQ:3.2 PL:[3.2, 0.0, 263.9] SR:10 DR:0 LR:-2.937 LO:18.91);ALT=T[chr6:52548876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52651164	+	chr6	52652644	+	.	25	0	2851467_1	49.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=2851467_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:52651164(+)-6:52652644(-)__6_52650501_52675501D;SPAN=1480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:124 GQ:49.1 PL:[49.1, 0.0, 250.4] SR:0 DR:25 LR:-48.93 LO:56.76);ALT=C[chr6:52652644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	52935944	+	chr6	52938277	+	.	2	6	2852539_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGCA;MAPQ=60;MATEID=2852539_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_6_52920001_52945001_171C;SPAN=2333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:6 DR:2 LR:3.394 LO:14.36);ALT=A[chr6:52938277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	53156763	+	chr6	53160440	+	.	0	11	2852945_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2852945_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_53140501_53165501_199C;SPAN=3677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:11 DR:0 LR:-9.219 LO:21.81);ALT=T[chr6:53160440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	53156805	+	chr6	53213612	+	.	19	0	2853442_1	51.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2853442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:53156805(+)-6:53213612(-)__6_53189501_53214501D;SPAN=56807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:43 GQ:51.2 PL:[51.2, 0.0, 51.2] SR:0 DR:19 LR:-51.07 LO:51.07);ALT=A[chr6:53213612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	53159291	+	chr6	53160437	+	.	0	11	2852964_1	4.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=2852964_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_53140501_53165501_218C;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:118 GQ:4.4 PL:[4.4, 0.0, 281.6] SR:11 DR:0 LR:-4.342 LO:20.98);ALT=T[chr6:53160437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	53159326	+	chr6	53213622	+	.	12	0	2853443_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2853443_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:53159326(+)-6:53213622(-)__6_53189501_53214501D;SPAN=54296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=A[chr6:53213622[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	53160507	+	chr6	53213613	+	.	15	13	2853444_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=2853444_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_53189501_53214501_113C;SPAN=53106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:43 GQ:47.9 PL:[47.9, 0.0, 54.5] SR:13 DR:15 LR:-47.77 LO:47.81);ALT=T[chr6:53213613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	74229149	+	chr9	118862122	-	.	18	35	2902286_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=T;MAPQ=22;MATEID=2902286_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_74210501_74235501_240C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:91 GQ:91.1 PL:[127.4, 0.0, 91.1] SR:35 DR:18 LR:-127.5 LO:127.5);ALT=T]chr9:118862122];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	74865448	+	chr6	74866585	+	.	25	19	2903459_1	96.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GAAAACCAAGTTATT;MAPQ=60;MATEID=2903459_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_74847501_74872501_157C;SPAN=1137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:57 GQ:40.7 PL:[96.8, 0.0, 40.7] SR:19 DR:25 LR:-97.99 LO:97.99);ALT=T[chr6:74866585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	44886653	+	chr6	78846111	+	.	8	0	5724419_1	20.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5724419_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:78846111(-)-14:44886653(+)__14_44884001_44909001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:21 GQ:20.9 PL:[20.9, 0.0, 27.5] SR:0 DR:8 LR:-20.72 LO:20.82);ALT=]chr14:44886653]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	79688430	+	chr6	79692603	+	.	7	1	2913918_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2913918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_79674001_79699001_92C;SPAN=4173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:66 GQ:5.3 PL:[5.3, 0.0, 153.8] SR:1 DR:7 LR:-5.226 LO:13.76);ALT=T[chr6:79692603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	79692840	+	chr6	79697925	+	CTGCCATCACTGTGCCATGCTCTCTCTTCTTCTTCGGATGTTCCACCACTGACAGCAACTACTTCGCCTT	0	18	2913934_1	37.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTGCCATCACTGTGCCATGCTCTCTCTTCTTCTTCGGATGTTCCACCACTGACAGCAACTACTTCGCCTT;MAPQ=60;MATEID=2913934_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_79674001_79699001_276C;SPAN=5085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:83 GQ:37.1 PL:[37.1, 0.0, 162.5] SR:18 DR:0 LR:-36.93 LO:41.51);ALT=A[chr6:79697925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	79727301	+	chr6	79735236	+	AGCACTAAAAGAAGAACAGATCATTTGAACTCCAGGCCGAGGGCGCTCTGTAAATTTTGCAGGTCTTGGG	6	12	2913465_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGCACTAAAAGAAGAACAGATCATTTGAACTCCAGGCCGAGGGCGCTCTGTAAATTTTGCAGGTCTTGGG;MAPQ=60;MATEID=2913465_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_79723001_79748001_252C;SPAN=7935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:12 DR:6 LR:-26.17 LO:31.35);ALT=C[chr6:79735236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	79770536	+	chr6	79787746	+	AGATTCTGGTAGGTCCTGGGATGCTCCTTCCCGGTCCAGTCGGTGCGCCGGGGCAGCAGCTCCTTCTCGGCCACCTCGCGGATCAGCACCTGAGCCGCCTGCTGACAGGGTCCATCTTCCAGGAACCGGGCGATGAGGAAGTAGAGCT	0	18	2913679_1	49.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGATTCTGGTAGGTCCTGGGATGCTCCTTCCCGGTCCAGTCGGTGCGCCGGGGCAGCAGCTCCTTCTCGGCCACCTCGCGGATCAGCACCTGAGCCGCCTGCTGACAGGGTCCATCTTCCAGGAACCGGGCGATGAGGAAGTAGAGCT;MAPQ=60;MATEID=2913679_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_6_79747501_79772501_321C;SPAN=17210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:37 GQ:39.5 PL:[49.4, 0.0, 39.5] SR:18 DR:0 LR:-49.44 LO:49.44);ALT=C[chr6:79787746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	79912141	+	chr6	79944262	+	.	29	0	2914162_1	84.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=2914162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:79912141(+)-6:79944262(-)__6_79943501_79968501D;SPAN=32121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:41 GQ:12.2 PL:[84.8, 0.0, 12.2] SR:0 DR:29 LR:-87.4 LO:87.4);ALT=T[chr6:79944262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	80071347	+	chr6	80073342	+	.	13	0	2914412_1	22.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=2914412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:80071347(+)-6:80073342(-)__6_80066001_80091001D;SPAN=1995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:77 GQ:22.1 PL:[22.1, 0.0, 164.0] SR:0 DR:13 LR:-22.05 LO:28.39);ALT=A[chr6:80073342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	80073657	+	chr6	80071662	+	.	22	0	2914416_1	57.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2914416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:80071662(-)-6:80073657(+)__6_80066001_80091001D;SPAN=1995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:55 GQ:57.8 PL:[57.8, 0.0, 74.3] SR:0 DR:22 LR:-57.72 LO:57.86);ALT=]chr6:80073657]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	87865477	+	chr6	87925618	+	.	0	7	2931270_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=2931270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_87906001_87931001_25C;SPAN=60141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:35 GQ:13.7 PL:[13.7, 0.0, 69.8] SR:7 DR:0 LR:-13.62 LO:15.86);ALT=G[chr6:87925618[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	88272505	+	chr6	88273848	+	.	0	6	2932211_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2932211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_88273501_88298501_317C;SPAN=1343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:37 GQ:9.8 PL:[9.8, 0.0, 79.1] SR:6 DR:0 LR:-9.782 LO:12.99);ALT=T[chr6:88273848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	88273997	+	chr6	88299628	+	.	10	0	2932406_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2932406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:88273997(+)-6:88299628(-)__6_88298001_88323001D;SPAN=25631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:0 DR:10 LR:-22.44 LO:23.91);ALT=T[chr6:88299628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	88521541	+	chr6	88519332	+	.	4	2	2932795_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCAACTTG;MAPQ=60;MATEID=2932795_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_88518501_88543501_298C;SPAN=2209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:77 GQ:4.2 PL:[0.0, 4.2, 194.7] SR:2 DR:4 LR:4.356 LO:8.718);ALT=]chr6:88521541]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	89326733	-	chr18	77406999	+	.	6	22	6686820_1	72.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=TGTAATCCCAGCACTTTGGGAGGCC;MAPQ=31;MATEID=6686820_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_18_77395501_77420501_89C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:21 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:22 DR:6 LR:-72.62 LO:72.62);ALT=[chr18:77406999[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	89791155	+	chr6	89793470	+	.	18	82	2935964_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2935964_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_89768001_89793001_205C;SPAN=2315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:38 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:82 DR:18 LR:-267.4 LO:267.4);ALT=T[chr6:89793470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	89864623	+	chr6	89868044	+	.	3	5	2936131_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=2936131_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_89866001_89891001_226C;SPAN=3421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:38 GQ:12.8 PL:[12.8, 0.0, 78.8] SR:5 DR:3 LR:-12.81 LO:15.58);ALT=T[chr6:89868044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90039677	+	chr6	90042805	+	.	10	11	2936599_1	41.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=2936599_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_90037501_90062501_361C;SPAN=3128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:80 GQ:41 PL:[41.0, 0.0, 153.2] SR:11 DR:10 LR:-41.05 LO:44.68);ALT=C[chr6:90042805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90042926	+	chr6	90045020	+	.	4	3	2936604_1	1.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=2936604_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAA;SCTG=c_6_90037501_90062501_361C;SPAN=2094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:80 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:3 DR:4 LR:-1.433 LO:13.15);ALT=T[chr6:90045020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90048029	+	chr6	90052042	+	TACTCCACGAAGGCTGCCAAGTTTCAGGATGATGGCCTGAGATGCTCAAACAGATTTTCTTGCCCACTTCAAATCGACCATTAG	0	12	2936620_1	23.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TACTCCACGAAGGCTGCCAAGTTTCAGGATGATGGCCTGAGATGCTCAAACAGATTTTCTTGCCCACTTCAAATCGACCATTAG;MAPQ=60;MATEID=2936620_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_90037501_90062501_154C;SPAN=4013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:12 DR:0 LR:-22.81 LO:27.0);ALT=A[chr6:90052042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90048263	+	chr6	90052042	+	.	5	4	2936621_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=2936621_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_6_90037501_90062501_154C;SPAN=3779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:58 GQ:14 PL:[14.0, 0.0, 126.2] SR:4 DR:5 LR:-14.0 LO:19.3);ALT=C[chr6:90052042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90052176	+	chr6	90062258	+	CTAAAGGCTGCGCATGGTAATGATCTGTTGGATCTTTCAATTCTGCCGCTTCTTTCATTAAACGTTTAACAG	13	68	2936632_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTAAAGGCTGCGCATGGTAATGATCTGTTGGATCTTTCAATTCTGCCGCTTCTTTCATTAAACGTTTAACAG;MAPQ=60;MATEID=2936632_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_90037501_90062501_2C;SPAN=10082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:90 GQ:11.9 PL:[206.6, 0.0, 11.9] SR:68 DR:13 LR:-217.1 LO:217.1);ALT=T[chr6:90062258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	90053524	+	chr6	90062344	+	.	29	0	2936635_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2936635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:90053524(+)-6:90062344(-)__6_90037501_90062501D;SPAN=8820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:82 GQ:73.7 PL:[73.7, 0.0, 123.2] SR:0 DR:29 LR:-73.51 LO:74.26);ALT=A[chr6:90062344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	101315916	+	chr6	101328937	+	.	0	10	2960221_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2960221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_101307501_101332501_202C;SPAN=13021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:10 DR:0 LR:-8.085 LO:19.77);ALT=T[chr6:101328937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55518500	+	chr6	101337435	+	.	18	0	5750195_1	48.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5750195_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:101337435(-)-14:55518500(+)__14_55517001_55542001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:39 GQ:45.5 PL:[48.8, 0.0, 45.5] SR:0 DR:18 LR:-48.86 LO:48.86);ALT=]chr14:55518500]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	102283809	+	chr8	107556938	+	.	34	0	4012507_1	98.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4012507_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:102283809(+)-8:107556938(-)__8_107555001_107580001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:52 GQ:25.7 PL:[98.3, 0.0, 25.7] SR:0 DR:34 LR:-100.3 LO:100.3);ALT=T[chr8:107556938[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	106764142	+	chr6	106773401	+	.	10	4	2972352_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2972352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_106771001_106796001_418C;SPAN=9259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:53 GQ:22.1 PL:[22.1, 0.0, 104.6] SR:4 DR:10 LR:-21.95 LO:25.13);ALT=C[chr6:106773401[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	107307807	+	chr8	105231728	+	CCATGATCAGTGGCCATG	32	57	2973824_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;INSERTION=CCATGATCAGTGGCCATG;MAPQ=60;MATEID=2973824_2;MATENM=1;NM=1;NUMPARTS=3;SCTG=c_6_107285501_107310501_193C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:42 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:57 DR:32 LR:-201.3 LO:201.3);ALT=C[chr8:105231728[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	105231899	+	chr6	107307808	+	CCATGATCAGTGGCCATG	32	38	4006369_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AC;INSERTION=CCATGATCAGTGGCCATG;MAPQ=60;MATEID=4006369_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_8_105227501_105252501_237C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:53 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:38 DR:32 LR:-178.2 LO:178.2);ALT=]chr8:105231899]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr22	39710816	+	chr6	108326050	+	.	10	0	7299320_1	14.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=7299320_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:108326050(-)-22:39710816(+)__22_39690001_39715001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:0 DR:10 LR:-14.86 LO:21.25);ALT=]chr22:39710816]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	108533458	+	chr6	108535701	+	.	6	6	2977329_1	32.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=2977329_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_108535001_108560001_88C;SPAN=2243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:25 GQ:26.3 PL:[32.9, 0.0, 26.3] SR:6 DR:6 LR:-32.86 LO:32.86);ALT=C[chr6:108535701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	108533460	+	chr6	108544153	+	.	4	3	2977330_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=2977330_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_108535001_108560001_71C;SPAN=10693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:46 GQ:10.7 PL:[10.7, 0.0, 99.8] SR:3 DR:4 LR:-10.64 LO:14.94);ALT=T[chr6:108544153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	108535828	+	chr6	108544152	+	.	4	42	2977333_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=2977333_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_108535001_108560001_195C;SPAN=8324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:96 GQ:99 PL:[122.6, 0.0, 109.4] SR:42 DR:4 LR:-122.6 LO:122.6);ALT=T[chr6:108544152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	108535875	+	chr6	108581963	+	.	16	0	2977548_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2977548_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:108535875(+)-6:108581963(-)__6_108559501_108584501D;SPAN=46088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:60 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:0 DR:16 LR:-36.56 LO:38.57);ALT=A[chr6:108581963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	108544251	+	chr6	108581964	+	.	72	99	2977550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=2977550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_108559501_108584501_115C;SPAN=37713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:62 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:99 DR:72 LR:-406.0 LO:406.0);ALT=T[chr6:108581964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109169755	+	chr6	109175424	+	.	12	0	2978975_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2978975_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:109169755(+)-6:109175424(-)__6_109172001_109197001D;SPAN=5669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=T[chr6:109175424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109322740	+	chr6	109330681	+	.	11	0	2979402_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2979402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:109322740(+)-6:109330681(-)__6_109319001_109344001D;SPAN=7941;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:0 DR:11 LR:-13.82 LO:22.76);ALT=A[chr6:109330681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109323583	+	chr6	109330635	+	.	9	0	2979408_1	12.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=2979408_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:109323583(+)-6:109330635(-)__6_109319001_109344001D;SPAN=7052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=A[chr6:109330635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109699176	+	chr6	109700782	+	.	0	17	2980156_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=2980156_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_109686501_109711501_84C;SPAN=1606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:74 GQ:36.2 PL:[36.2, 0.0, 141.8] SR:17 DR:0 LR:-36.07 LO:39.69);ALT=T[chr6:109700782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109700869	+	chr6	109703407	+	.	0	28	2980159_1	73.0	.	EVDNC=ASSMB;HOMSEQ=CTGG;MAPQ=60;MATEID=2980159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_109686501_109711501_322C;SPAN=2538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:72 GQ:73.1 PL:[73.1, 0.0, 99.5] SR:28 DR:0 LR:-72.92 LO:73.18);ALT=G[chr6:109703407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	109803292	+	chr6	109804305	+	.	10	0	2980631_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2980631_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:109803292(+)-6:109804305(-)__6_109784501_109809501D;SPAN=1013;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-13.77 LO:20.98);ALT=G[chr6:109804305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110012704	+	chr6	110036281	+	.	0	7	2981079_1	12.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2981079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110005001_110030001_193C;SPAN=23577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:38 GQ:12.8 PL:[12.8, 0.0, 78.8] SR:7 DR:0 LR:-12.81 LO:15.58);ALT=T[chr6:110036281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	146184521	+	chr6	110181755	+	.	6	6	2981671_1	25.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=GGTTGGGGTACTTGCCCCTCCCCTAGAAAAGCAGGACTTGCC;MAPQ=28;MATEID=2981671_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_6_110176501_110201501_316C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:54 GQ:25.1 PL:[25.1, 0.0, 104.3] SR:6 DR:6 LR:-24.98 LO:27.82);ALT=]chr8:146184521]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	110501837	+	chr6	110514383	+	.	0	11	2982157_1	14.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=2982157_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110495001_110520001_336C;SPAN=12546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:80 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:11 DR:0 LR:-14.64 LO:22.95);ALT=G[chr6:110514383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110514471	+	chr6	110522759	+	.	0	17	2982182_1	45.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2982182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110495001_110520001_277C;SPAN=8288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:17 DR:0 LR:-45.01 LO:45.06);ALT=G[chr6:110522759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110522892	+	chr6	110528708	+	.	0	10	2982235_1	12.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=2982235_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110519501_110544501_79C;SPAN=5816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:76 GQ:12.5 PL:[12.5, 0.0, 170.9] SR:10 DR:0 LR:-12.42 LO:20.66);ALT=T[chr6:110528708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110528794	+	chr6	110530285	+	.	2	8	2982243_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=2982243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110519501_110544501_56C;SPAN=1491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:8 DR:2 LR:-10.2 LO:18.38);ALT=T[chr6:110530285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110778201	+	chr6	110797724	+	.	10	0	2982858_1	26.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2982858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:110778201(+)-6:110797724(-)__6_110789001_110814001D;SPAN=19523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:0 DR:10 LR:-26.24 LO:26.3);ALT=A[chr6:110797724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	110796866	+	chr6	110800510	+	.	2	5	2982878_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=2982878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_110789001_110814001_150C;SPAN=3644;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:72 GQ:3.8 PL:[3.8, 0.0, 168.8] SR:5 DR:2 LR:-3.6 LO:13.48);ALT=G[chr6:110800510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	111280048	+	chrX	106374932	+	.	52	0	7492079_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7492079_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:111280048(+)-23:106374932(-)__23_106354501_106379501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:26 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=A[chrX:106374932[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	111303351	+	chr6	111306208	+	.	8	0	2984544_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2984544_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:111303351(+)-6:111306208(-)__6_111279001_111304001D;SPAN=2857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=A[chr6:111306208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	111303364	+	chr20	34340812	+	.	8	0	6992386_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6992386_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:111303364(+)-20:34340812(-)__20_34324501_34349501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:0 DR:8 LR:-14.49 LO:17.76);ALT=G[chr20:34340812[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	113730685	+	chr19	58938759	-	.	2	5	2990307_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAAGAAA;MAPQ=60;MATEID=2990307_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_113729001_113754001_124C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:19 GQ:14.6 PL:[14.6, 0.0, 31.1] SR:5 DR:2 LR:-14.66 LO:15.0);ALT=A]chr19:58938759];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	113730691	-	chr19	58938657	+	.	9	0	6880456_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6880456_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:113730691(-)-19:58938657(-)__19_58922501_58947501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:30 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.58 LO:22.25);ALT=[chr19:58938657[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	114262253	+	chr6	114264515	+	CTTTGGTATCTGTTTTTTCACCACTGTTGTCCTTGGATTTATCTTCTTCCTTAACGT	12	15	2991701_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTTTGGTATCTGTTTTTTCACCACTGTTGTCCTTGGATTTATCTTCTTCCTTAACGT;MAPQ=60;MATEID=2991701_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_114243501_114268501_60C;SPAN=2262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:85 GQ:56.3 PL:[56.3, 0.0, 148.7] SR:15 DR:12 LR:-56.2 LO:58.56);ALT=C[chr6:114264515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	114270425	+	chr6	114274440	+	.	3	4	2991580_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=2991580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_114268001_114293001_253C;SPAN=4015;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:60 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:4 DR:3 LR:-6.852 LO:14.07);ALT=C[chr6:114274440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	114281183	+	chr6	114292017	+	.	12	22	2991620_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TCACC;MAPQ=60;MATEID=2991620_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_6_114268001_114293001_320C;SPAN=10834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:87 GQ:62.3 PL:[62.3, 0.0, 148.1] SR:22 DR:12 LR:-62.26 LO:64.22);ALT=C[chr6:114292017[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	116368767	+	chr9	6360629	-	TAGCTACAAAATTAGCCAGGCATGGTGTCACATGCTTGT	4	66	2995894_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;INSERTION=TAGCTACAAAATTAGCCAGGCATGGTGTCACATGCTTGT;MAPQ=60;MATEID=2995894_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_6_116350501_116375501_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:25 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:66 DR:4 LR:-194.7 LO:194.7);ALT=T]chr9:6360629];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	116750908	+	chr6	116751911	-	.	8	0	2996701_1	3.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=2996701_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:116750908(+)-6:116751911(+)__6_116742501_116767501D;SPAN=1003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=G]chr6:116751911];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	116774807	+	chr7	26241470	-	.	27	0	3217813_1	79.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=3217813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:116774807(+)-7:26241470(+)__7_26239501_26264501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:26 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:0 DR:27 LR:-79.22 LO:79.22);ALT=C]chr7:26241470];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	116892818	+	chr6	116895219	+	.	15	15	2997031_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2997031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_116889501_116914501_39C;SPAN=2401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:88 GQ:52.1 PL:[52.1, 0.0, 161.0] SR:15 DR:15 LR:-52.08 LO:55.21);ALT=G[chr6:116895219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	116892818	+	chr6	116901455	+	.	9	32	2997032_1	94.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=2997032_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_116889501_116914501_260C;SPAN=8637;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:90 GQ:94.4 PL:[94.4, 0.0, 124.1] SR:32 DR:9 LR:-94.45 LO:94.67);ALT=G[chr6:116901455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	116892818	+	chr12	77151016	+	.	20	12	5254544_1	93.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGAGTCCATCTACCCTGACTCCTTCACAG;MAPQ=60;MATEID=5254544_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_12_77150501_77175501_56C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:44 GQ:11.3 PL:[93.8, 0.0, 11.3] SR:12 DR:20 LR:-97.22 LO:97.22);ALT=G[chr12:77151016[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr6	116895334	+	chr6	116901456	+	.	0	14	2997041_1	23.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2997041_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_116889501_116914501_334C;SPAN=6122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:14 DR:0 LR:-23.73 LO:30.57);ALT=G[chr6:116901456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	119013928	+	chr6	119011719	+	.	20	15	3001674_1	73.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=3001674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_118996501_119021501_44C;SPAN=2209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:84 GQ:73.1 PL:[73.1, 0.0, 129.2] SR:15 DR:20 LR:-72.97 LO:73.87);ALT=]chr6:119013928]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr6	119012288	+	chr6	119013928	+	TACATTGTCA	0	22	3001678_1	45.0	.	EVDNC=ASSMB;INSERTION=TACATTGTCA;MAPQ=60;MATEID=3001678_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_118996501_119021501_255C;SPAN=1640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:100 GQ:45.5 PL:[45.5, 0.0, 197.3] SR:22 DR:0 LR:-45.53 LO:50.89);ALT=A[chr6:119013928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	131057569	-	chr9	94148177	+	.	27	52	3028014_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3028014_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_131050501_131075501_19C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:29 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:52 DR:27 LR:-208.0 LO:208.0);ALT=[chr9:94148177[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	131678470	-	chr22	31751841	+	.	11	0	7267931_1	23.0	.	DISC_MAPQ=11;EVDNC=DSCRD;IMPRECISE;MAPQ=11;MATEID=7267931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:131678470(-)-22:31751841(-)__22_31727501_31752501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:47 GQ:23.6 PL:[23.6, 0.0, 89.6] SR:0 DR:11 LR:-23.58 LO:25.79);ALT=[chr22:31751841[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	136710657	+	chr6	136742839	+	AGCTGTTTCTCCCGTTCCTCACGTCGCTCCCGGGCCAGCCGCTGCCGGTCATCAACACGTAACACAGGCGGAGGGT	2	13	3041000_1	33.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=AGCTGTTTCTCCCGTTCCTCACGTCGCTCCCGGGCCAGCCGCTGCCGGTCATCAACACGTAACACAGGCGGAGGGT;MAPQ=60;MATEID=3041000_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_136710001_136735001_247C;SPAN=32182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:46 GQ:33.8 PL:[33.8, 0.0, 76.7] SR:13 DR:2 LR:-33.75 LO:34.71);ALT=T[chr6:136742839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	137105413	+	chr6	137106552	+	.	9	6	3041830_1	12.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=38;MATEID=3041830_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_137102001_137127001_22C;SPAN=1139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:77 GQ:12.2 PL:[12.2, 0.0, 173.9] SR:6 DR:9 LR:-12.15 LO:20.6);ALT=G[chr6:137106552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	137143934	+	chr6	137146351	+	.	0	12	3042118_1	21.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3042118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_137126501_137151501_346C;SPAN=2417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:12 DR:0 LR:-21.73 LO:26.64);ALT=G[chr6:137146351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	137528220	+	chr6	137540379	+	.	9	0	3043011_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3043011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:137528220(+)-6:137540379(-)__6_137518501_137543501D;SPAN=12159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:71 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:0 DR:9 LR:-10.47 LO:18.44);ALT=A[chr6:137540379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	138725734	+	chr6	138727106	+	CCCGGAAGTTATGAGATCCGACACTATGGACCAGCCAAGTGGGTCAGCACGTCCGTGGAGTCTATGGACTGGGATTCAGCCATCCAGACGGGCTTTACGAAACTGAACAGCTACATTCAAGGCAAAAACGAGAA	4	36	3045533_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCCGGAAGTTATGAGATCCGACACTATGGACCAGCCAAGTGGGTCAGCACGTCCGTGGAGTCTATGGACTGGGATTCAGCCATCCAGACGGGCTTTACGAAACTGAACAGCTACATTCAAGGCAAAAACGAGAA;MAPQ=60;MATEID=3045533_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_6_138719001_138744001_36C;SPAN=1372;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:80 GQ:90.5 PL:[103.7, 0.0, 90.5] SR:36 DR:4 LR:-103.8 LO:103.8);ALT=G[chr6:138727106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	138726463	+	chr6	138734015	+	.	14	0	3045536_1	25.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3045536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:138726463(+)-6:138734015(-)__6_138719001_138744001D;SPAN=7552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:76 GQ:25.7 PL:[25.7, 0.0, 157.7] SR:0 DR:14 LR:-25.62 LO:31.17);ALT=C[chr6:138734015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	138727290	+	chr6	138734016	+	.	11	27	3045539_1	91.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=3045539_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_138719001_138744001_35C;SPAN=6726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:88 GQ:91.7 PL:[91.7, 0.0, 121.4] SR:27 DR:11 LR:-91.69 LO:91.93);ALT=T[chr6:138734016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	138774059	-	chr15	23717166	+	GTATATTATC	12	21	5901300_1	80.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=GTATATTATC;MAPQ=60;MATEID=5901300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_23716001_23741001_452C;SPAN=-1;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:68 GQ:80.6 PL:[80.6, 0.0, 83.9] SR:21 DR:12 LR:-80.61 LO:80.61);ALT=[chr15:23717166[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	138774182	+	chr15	23712619	-	.	18	34	5902474_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TG;MAPQ=60;MATEID=5902474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_23691501_23716501_789C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:84 GQ:83 PL:[119.3, 0.0, 83.0] SR:34 DR:18 LR:-119.5 LO:119.5);ALT=G]chr15:23712619];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	139095007	+	chr6	139097213	+	.	23	0	3046770_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3046770_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:139095007(+)-6:139097213(-)__6_139086501_139111501D;SPAN=2206;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:93 GQ:50.9 PL:[50.9, 0.0, 173.0] SR:0 DR:23 LR:-50.73 LO:54.56);ALT=G[chr6:139097213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	139097415	+	chr6	139100957	+	.	5	8	3046774_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3046774_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_139086501_139111501_59C;SPAN=3542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:70 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:8 DR:5 LR:-17.35 LO:23.65);ALT=G[chr6:139100957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	95384452	+	chr6	139294720	+	.	5	20	3047211_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3047211_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_139282501_139307501_316C;SPAN=-1;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:20 DR:5 LR:-65.7 LO:65.7);ALT=]chr14:95384452]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr6	139350013	+	chr6	139355290	+	.	31	40	3047348_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3047348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_139331501_139356501_335C;SPAN=5277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:96 GQ:76.4 PL:[155.6, 0.0, 76.4] SR:40 DR:31 LR:-157.0 LO:157.0);ALT=G[chr6:139355290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	139355358	+	chr6	139363856	+	.	0	105	3047233_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3047233_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_139356001_139381001_139C;SPAN=8498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:62 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:105 DR:0 LR:-310.3 LO:310.3);ALT=A[chr6:139363856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	149433459	+	chr20	16718037	-	.	12	0	6938924_1	27.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6938924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:149433459(+)-20:16718037(+)__20_16709001_16734001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=T]chr20:16718037];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	149433833	+	chr20	16710782	-	.	33	0	6938925_1	92.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=6938925_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:149433833(+)-20:16710782(+)__20_16709001_16734001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:62 GQ:56 PL:[92.3, 0.0, 56.0] SR:0 DR:33 LR:-92.54 LO:92.54);ALT=A]chr20:16710782];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr6	149862723	+	chr6	149867072	+	.	12	3	3070758_1	28.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3070758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_149866501_149891501_186C;SPAN=4349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:42 GQ:28.4 PL:[28.4, 0.0, 71.3] SR:3 DR:12 LR:-28.23 LO:29.36);ALT=C[chr6:149867072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	149887671	+	chr6	149893417	+	.	10	8	3070890_1	36.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACAGG;MAPQ=60;MATEID=3070890_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_149891001_149916001_7C;SPAN=5746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:23 GQ:17 PL:[36.8, 0.0, 17.0] SR:8 DR:10 LR:-36.98 LO:36.98);ALT=G[chr6:149893417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	150071092	+	chr6	150092298	+	.	0	20	3072002_1	53.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3072002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_150087001_150112001_450C;SPAN=21206;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:45 GQ:53.9 PL:[53.9, 0.0, 53.9] SR:20 DR:0 LR:-53.83 LO:53.83);ALT=A[chr6:150092298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	150092404	+	chr6	150111089	+	TTCCAAGCAACAATCAGTGCTCCACACAT	0	10	3072021_1	11.0	.	EVDNC=ASSMB;INSERTION=TTCCAAGCAACAATCAGTGCTCCACACAT;MAPQ=60;MATEID=3072021_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_150087001_150112001_23C;SPAN=18685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:0 LR:-11.34 LO:20.42);ALT=T[chr6:150111089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	154620006	+	chr6	154621505	+	.	123	77	3082933_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GGAAGCTGAGGCAGGAG;MAPQ=60;MATEID=3082933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_154595001_154620001_361C;SPAN=1499;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:19 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:77 DR:123 LR:-452.2 LO:452.2);ALT=G[chr6:154621505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	154871426	-	chr6	154872453	+	.	11	0	3083442_1	15.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3083442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:154871426(-)-6:154872453(-)__6_154864501_154889501D;SPAN=1027;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:78 GQ:15.2 PL:[15.2, 0.0, 173.6] SR:0 DR:11 LR:-15.18 LO:23.09);ALT=[chr6:154872453[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	157699920	+	chr6	157703237	+	.	47	18	3090020_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCTCCCAGGTTCAAGCGATTCTCCTGCCTCAGCCTCCTGAGTAGCTGGGA;MAPQ=60;MATEID=3090020_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_6_157682001_157707001_3C;SPAN=3317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:38 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:18 DR:47 LR:-171.6 LO:171.6);ALT=A[chr6:157703237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	157739968	+	chr6	157744479	+	.	11	0	3090783_1	15.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=3090783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:157739968(+)-6:157744479(-)__6_157731001_157756001D;SPAN=4511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:0 DR:11 LR:-15.45 LO:23.15);ALT=A[chr6:157744479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	157744475	-	chr12	63396370	+	.	12	0	5220685_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5220685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:157744475(-)-12:63396370(-)__12_63381501_63406501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:47 GQ:26.9 PL:[26.9, 0.0, 86.3] SR:0 DR:12 LR:-26.88 LO:28.66);ALT=[chr12:63396370[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	158589482	+	chr6	158613006	+	.	45	0	3092858_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3092858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:158589482(+)-6:158613006(-)__6_158613001_158638001D;SPAN=23524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:36 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=G[chr6:158613006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	158864107	+	chr6	158865208	-	.	3	2	3093638_1	0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=GGAGGCGGAGGTTGCAGTGAGCCAAGATTGC;MAPQ=60;MATEID=3093638_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_6_158858001_158883001_99C;SPAN=1101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:2 DR:3 LR:6.574 LO:6.671);ALT=C]chr6:158865208];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	159058953	+	chr6	159065712	+	.	11	0	3094182_1	13.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3094182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:159058953(+)-6:159065712(-)__6_159054001_159079001D;SPAN=6759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:85 GQ:13.4 PL:[13.4, 0.0, 191.6] SR:0 DR:11 LR:-13.28 LO:22.64);ALT=C[chr6:159065712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159208238	+	chr6	159210318	+	.	0	13	3095247_1	23.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=3095247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_159201001_159226001_209C;SPAN=2080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:74 GQ:23 PL:[23.0, 0.0, 155.0] SR:13 DR:0 LR:-22.86 LO:28.64);ALT=G[chr6:159210318[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159208277	+	chr6	159240342	+	.	9	0	3095248_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3095248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:159208277(+)-6:159240342(-)__6_159201001_159226001D;SPAN=32065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.31 LO:22.09);ALT=A[chr6:159240342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159210403	+	chr6	159239114	+	.	0	7	3095259_1	13.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3095259_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_159201001_159226001_102C;SPAN=28711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:35 GQ:13.7 PL:[13.7, 0.0, 69.8] SR:7 DR:0 LR:-13.62 LO:15.86);ALT=T[chr6:159239114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159210437	+	chr6	159240345	+	.	9	0	3095260_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3095260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:159210437(+)-6:159240345(-)__6_159201001_159226001D;SPAN=29908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=T[chr6:159240345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	159968217	+	chr6	159970838	+	.	57	26	3096791_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGTACCACATTTTTTA;MAPQ=60;MATEID=3096791_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_159960501_159985501_195C;SPAN=2621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:59 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:26 DR:57 LR:-217.9 LO:217.9);ALT=A[chr6:159970838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	160183160	+	chr6	160188034	+	.	8	0	3097388_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3097388_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:160183160(+)-6:160188034(-)__6_160181001_160206001D;SPAN=4874;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-2.025 LO:15.08);ALT=C[chr6:160188034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	160184086	+	chr6	160188035	+	.	0	14	3097392_1	17.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3097392_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_160181001_160206001_121C;SPAN=3949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:106 GQ:17.6 PL:[17.6, 0.0, 238.7] SR:14 DR:0 LR:-17.5 LO:28.95);ALT=G[chr6:160188035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	160209176	+	chr6	160210437	+	.	8	29	3097174_1	83.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3097174_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_160205501_160230501_102C;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:95 GQ:83.3 PL:[83.3, 0.0, 146.0] SR:29 DR:8 LR:-83.2 LO:84.17);ALT=C[chr6:160210437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	160211615	+	chr6	160218316	+	.	11	0	3097185_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3097185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:160211615(+)-6:160218316(-)__6_160205501_160230501D;SPAN=6701;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:79 GQ:14.9 PL:[14.9, 0.0, 176.6] SR:0 DR:11 LR:-14.91 LO:23.02);ALT=C[chr6:160218316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	160212160	+	chr6	160218317	+	.	5	17	3097188_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3097188_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_160205501_160230501_206C;SPAN=6157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:78 GQ:48.2 PL:[48.2, 0.0, 140.6] SR:17 DR:5 LR:-48.19 LO:50.73);ALT=T[chr6:160218317[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	151134	+	chr7	160558	+	TGGCG	70	49	3125958_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=TGGCG;MAPQ=60;MATEID=3125958_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_147001_172001_320C;SPAN=9424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:77 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:49 DR:70 LR:-293.8 LO:293.8);ALT=A[chr7:160558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	220952	+	chr7	222061	+	.	21	0	3125799_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3125799_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:220952(+)-7:222061(-)__7_220501_245501D;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:80 GQ:47.6 PL:[47.6, 0.0, 146.6] SR:0 DR:21 LR:-47.65 LO:50.45);ALT=T[chr7:222061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	303019	+	chr7	304019	+	.	10	0	3126240_1	0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=3126240_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:303019(+)-7:304019(-)__7_294001_319001D;SPAN=1000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:165 GQ:11.5 PL:[0.0, 11.5, 422.5] SR:0 DR:10 LR:11.69 LO:17.13);ALT=A[chr7:304019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	916441	+	chr7	925690	+	.	0	15	3128617_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CAGGTAC;MAPQ=60;MATEID=3128617_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_906501_931501_80C;SPAN=9249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:103 GQ:21.8 PL:[21.8, 0.0, 226.4] SR:15 DR:0 LR:-21.61 LO:31.71);ALT=C[chr7:925690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1037442	+	chr7	1040104	+	.	0	7	3129237_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3129237_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1029001_1054001_269C;SPAN=2662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:7 DR:0 LR:1.818 LO:12.7);ALT=T[chr7:1040104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1040189	+	chr7	1049586	+	.	0	11	3129244_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3129244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1029001_1054001_208C;SPAN=9397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:96 GQ:10.4 PL:[10.4, 0.0, 221.6] SR:11 DR:0 LR:-10.3 LO:22.02);ALT=T[chr7:1049586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1049801	+	chr7	1067894	+	.	30	0	3129276_1	83.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3129276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:1049801(+)-7:1067894(-)__7_1029001_1054001D;SPAN=18093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:56 GQ:50.9 PL:[83.9, 0.0, 50.9] SR:0 DR:30 LR:-84.26 LO:84.26);ALT=A[chr7:1067894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1167020	+	chr7	1177823	+	.	11	0	3129858_1	24.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3129858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:1167020(+)-7:1177823(-)__7_1176001_1201001D;SPAN=10803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:43 GQ:24.8 PL:[24.8, 0.0, 77.6] SR:0 DR:11 LR:-24.66 LO:26.28);ALT=A[chr7:1177823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1185078	+	chr7	1187655	+	.	57	20	3129900_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CACTCTTAAGTTTT;MAPQ=60;MATEID=3129900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1176001_1201001_348C;SPAN=2577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:67 DP:1556 GQ:99 PL:[0.0, 199.9, 4179.0] SR:20 DR:57 LR:200.4 LO:104.6);ALT=T[chr7:1187655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1192862	+	chr7	1195089	+	.	3	4	3129933_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3129933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1176001_1201001_346C;SPAN=2227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:4 DR:3 LR:2.902 LO:12.57);ALT=T[chr7:1195089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1197939	+	chr7	1199706	+	.	23	0	3129960_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3129960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:1197939(+)-7:1199706(-)__7_1176001_1201001D;SPAN=1767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:111 GQ:46.1 PL:[46.1, 0.0, 221.0] SR:0 DR:23 LR:-45.85 LO:52.53);ALT=C[chr7:1199706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	1607488	+	chr7	1608760	+	.	0	14	3131294_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3131294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_1592501_1617501_260C;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:113 GQ:15.8 PL:[15.8, 0.0, 256.7] SR:14 DR:0 LR:-15.6 LO:28.53);ALT=T[chr7:1608760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2281944	+	chr7	2289489	+	.	12	0	3133578_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3133578_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2281944(+)-7:2289489(-)__7_2278501_2303501D;SPAN=7545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:119 GQ:7.4 PL:[7.4, 0.0, 281.3] SR:0 DR:12 LR:-7.372 LO:23.32);ALT=G[chr7:2289489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2281977	+	chr7	2284197	+	.	15	0	3133579_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3133579_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2281977(+)-7:2284197(-)__7_2278501_2303501D;SPAN=2220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:150 GQ:8.9 PL:[8.9, 0.0, 355.4] SR:0 DR:15 LR:-8.876 LO:29.09);ALT=C[chr7:2284197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2284362	+	chr7	2289490	+	.	67	97	3133587_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3133587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_2278501_2303501_64C;SPAN=5128;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:156 GQ:28.9 PL:[435.7, 28.9, 0.0] SR:97 DR:67 LR:-440.4 LO:440.4);ALT=G[chr7:2289490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2294806	+	chr7	2296509	+	.	2	7	3133627_1	0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3133627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_2278501_2303501_317C;SPAN=1703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:7 DR:2 LR:-0.6702 LO:14.89);ALT=T[chr7:2296509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2317940	+	chr7	2353962	+	.	19	0	3134176_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3134176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2317940(+)-7:2353962(-)__7_2352001_2377001D;SPAN=36022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:61 GQ:46.4 PL:[46.4, 0.0, 99.2] SR:0 DR:19 LR:-46.19 LO:47.34);ALT=T[chr7:2353962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2415165	+	chr7	2416583	+	.	3	5	3134009_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=3134009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_2401001_2426001_234C;SPAN=1418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:90 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:5 DR:3 LR:1.276 LO:12.77);ALT=G[chr7:2416583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2443333	+	chr7	2472194	+	.	22	0	3134403_1	59.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3134403_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2443333(+)-7:2472194(-)__7_2450001_2475001D;SPAN=28861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:50 GQ:59 PL:[59.0, 0.0, 62.3] SR:0 DR:22 LR:-59.08 LO:59.08);ALT=C[chr7:2472194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2587114	+	chr7	2593939	+	.	0	7	3135097_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3135097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_2572501_2597501_251C;SPAN=6825;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:112 GQ:6.9 PL:[0.0, 6.9, 283.8] SR:7 DR:0 LR:7.237 LO:12.09);ALT=T[chr7:2593939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	2875361	+	chr20	52831836	+	.	28	0	7062885_1	78.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=7062885_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:2875361(+)-20:52831836(-)__20_52822001_52847001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:53 GQ:48.5 PL:[78.2, 0.0, 48.5] SR:0 DR:28 LR:-78.38 LO:78.38);ALT=T[chr20:52831836[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	4081265	+	chr7	4082297	+	.	60	47	3140500_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3140500_2;MATENM=2;NM=2;NUMPARTS=2;SCTG=c_7_4067001_4092001_137C;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:65 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:47 DR:60 LR:-241.0 LO:241.0);ALT=C[chr7:4082297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	5013792	+	chr7	5015932	+	.	9	1	3144557_1	6.0	.	DISC_MAPQ=41;EVDNC=ASDIS;MAPQ=60;MATEID=3144557_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_4998001_5023001_119C;SPAN=2140;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:1 DR:9 LR:-6.73 LO:19.53);ALT=A[chr7:5015932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	5230126	+	chr7	5239207	+	.	0	9	3145249_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=50;MATEID=3145249_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_5218501_5243501_208C;SPAN=9081;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:99 GQ:2.9 PL:[2.9, 0.0, 237.2] SR:9 DR:0 LR:-2.887 LO:17.06);ALT=T[chr7:5239207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	5267843	+	chr7	5269238	+	.	0	4	3145596_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3145596_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_5267501_5292501_277C;SPAN=1395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:123 GQ:19.8 PL:[0.0, 19.8, 336.6] SR:4 DR:0 LR:20.12 LO:5.753);ALT=G[chr7:5269238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	5831459	+	chr19	8538236	+	.	22	35	6718686_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TCGGGAGGCTGAGGCAG;MAPQ=60;MATEID=6718686_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_19_8526001_8551001_346C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:32 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:35 DR:22 LR:-155.1 LO:155.1);ALT=G[chr19:8538236[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	6049072	+	chr7	6054774	+	.	9	0	3149962_1	11.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3149962_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:6049072(+)-7:6054774(-)__7_6027001_6052001D;SPAN=5702;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=G[chr7:6054774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6084294	+	chr7	6085700	+	.	0	5	3150027_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3150027_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6076001_6101001_48C;SPAN=1406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:85 GQ:6.3 PL:[0.0, 6.3, 217.8] SR:5 DR:0 LR:6.524 LO:8.497);ALT=T[chr7:6085700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6094336	+	chr7	6098597	+	.	12	12	3150079_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3150079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6076001_6101001_446C;SPAN=4261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:126 GQ:22.1 PL:[22.1, 0.0, 282.8] SR:12 DR:12 LR:-21.98 LO:35.32);ALT=C[chr7:6098597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6485736	+	chr7	6487377	+	.	0	8	3151852_1	0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=3151852_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6468001_6493001_348C;SPAN=1641;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:8 DR:0 LR:-0.1283 LO:14.81);ALT=C[chr7:6487377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6509387	+	chr7	6513813	+	.	0	17	3152128_1	21.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3152128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6492501_6517501_400C;SPAN=4426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:129 GQ:21.2 PL:[21.2, 0.0, 291.8] SR:17 DR:0 LR:-21.17 LO:35.14);ALT=T[chr7:6513813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6509428	+	chr7	6523694	+	.	14	0	3152162_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3152162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:6509428(+)-7:6523694(-)__7_6517001_6542001D;SPAN=14266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:61 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:0 DR:14 LR:-29.69 LO:32.68);ALT=C[chr7:6523694[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6513916	+	chr7	6523596	+	.	0	58	3152163_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=3152163_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6517001_6542001_137C;SPAN=9680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:50 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:58 DR:0 LR:-171.6 LO:171.6);ALT=C[chr7:6523596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	6618351	+	chr7	6620186	+	.	2	10	3152504_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3152504_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_6615001_6640001_313C;SPAN=1835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:107 GQ:10.7 PL:[10.7, 0.0, 248.3] SR:10 DR:2 LR:-10.62 LO:23.9);ALT=T[chr7:6620186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	7583516	+	chr7	10708427	-	.	21	117	3166635_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3166635_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_10706501_10731501_20C;SPAN=3124911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:119 DP:67 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:117 DR:21 LR:-353.2 LO:353.2);ALT=G]chr7:10708427];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	7677628	+	chr7	7680003	+	.	22	0	3156873_1	45.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=3156873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:7677628(+)-7:7680003(-)__7_7668501_7693501D;SPAN=2375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:102 GQ:45.2 PL:[45.2, 0.0, 200.3] SR:0 DR:22 LR:-44.99 LO:50.68);ALT=T[chr7:7680003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	8463551	+	chr7	8465542	+	.	61	26	3159575_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=3159575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_8452501_8477501_231C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:67 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:26 DR:61 LR:-214.6 LO:214.6);ALT=A[chr7:8465542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	9634650	+	chr7	9635978	+	.	123	69	3163237_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGAAAAGAGACTACTG;MAPQ=60;MATEID=3163237_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_9628501_9653501_19C;SPAN=1328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:152 DP:44 GQ:40.9 PL:[448.9, 40.9, 0.0] SR:69 DR:123 LR:-448.9 LO:448.9);ALT=G[chr7:9635978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	10491065	-	chr11	122932781	+	.	91	0	5033453_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5033453_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:10491065(-)-11:122932781(-)__11_122916501_122941501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:91 DP:165 GQ:99 PL:[255.8, 0.0, 143.6] SR:0 DR:91 LR:-257.3 LO:257.3);ALT=[chr11:122932781[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	11014572	+	chr7	11021996	+	.	0	35	3167568_1	83.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=3167568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_11000501_11025501_182C;SPAN=7424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:119 GQ:83.3 PL:[83.3, 0.0, 205.4] SR:35 DR:0 LR:-83.3 LO:86.15);ALT=G[chr7:11021996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	19738352	+	chr7	19739695	+	.	0	13	3194931_1	14.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=3194931_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_19722501_19747501_365C;SPAN=1343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:104 GQ:14.9 PL:[14.9, 0.0, 236.0] SR:13 DR:0 LR:-14.74 LO:26.55);ALT=T[chr7:19739695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	19744545	+	chr7	19748386	+	.	10	10	3194947_1	37.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3194947_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_19722501_19747501_232C;SPAN=3841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:45 GQ:37.4 PL:[37.4, 0.0, 70.4] SR:10 DR:10 LR:-37.32 LO:37.92);ALT=T[chr7:19748386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	20369409	+	chr7	20371290	+	.	9	0	3196581_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3196581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:20369409(+)-7:20371290(-)__7_20359501_20384501D;SPAN=1881;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:0 DR:9 LR:-2.075 LO:16.94);ALT=G[chr7:20371290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	20707288	-	chr12	120357808	+	TTTGCCCTGCCTCT	28	55	5364021_1	99.0	.	DISC_MAPQ=10;EVDNC=ASDIS;INSERTION=TTTGCCCTGCCTCT;MAPQ=2;MATEID=5364021_2;MATENM=0;NM=23;NUMPARTS=2;SCTG=c_12_120344001_120369001_147C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:24 GQ:21 PL:[231.0, 21.0, 0.0] SR:55 DR:28 LR:-231.1 LO:231.1);ALT=[chr12:120357808[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	26230749	+	chr7	26232115	+	.	0	9	3217619_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=3217619_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26215001_26240001_46C;SPAN=1366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:149 GQ:10.6 PL:[0.0, 10.6, 382.8] SR:9 DR:0 LR:10.66 LO:15.4);ALT=C[chr7:26232115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26233316	+	chr7	26235465	+	.	13	50	3217638_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=3217638_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26215001_26240001_244C;SPAN=2149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:139 GQ:99 PL:[163.7, 0.0, 173.6] SR:50 DR:13 LR:-163.7 LO:163.7);ALT=T[chr7:26235465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26233316	+	chr7	26236021	+	CCAGGTCCTCCTCCATACCCATTATAGCCATCCCCAAATCCACGTCCACTGCCATATCCAT	43	75	3217639_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCAGGTCCTCCTCCATACCCATTATAGCCATCCCCAAATCCACGTCCACTGCCATATCCAT;MAPQ=60;MATEID=3217639_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26215001_26240001_244C;SPAN=2705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:131 GQ:8.7 PL:[333.3, 8.7, 0.0] SR:75 DR:43 LR:-346.1 LO:346.1);ALT=T[chr7:26236021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26237488	+	chr7	26240192	+	.	82	19	3217816_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3217816_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26239501_26264501_355C;SPAN=2704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:101 DP:135 GQ:29.6 PL:[296.9, 0.0, 29.6] SR:19 DR:82 LR:-309.4 LO:309.4);ALT=T[chr7:26240192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26241365	-	chr15	40854180	+	.	23	54	5931745_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;MAPQ=60;MATEID=5931745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40841501_40866501_163C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:33 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:54 DR:23 LR:-201.3 LO:201.3);ALT=[chr15:40854180[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	26241446	+	chr7	26245987	+	AATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA	33	97	3217824_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=GGCTCTGCCTCTTCAACTTTTTTACTCTTTCCATTCTGTTTTTTTCCCATTTTTTGCAATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA;INSERTION=AATGTAGTTTTGTTGGAGGCCATTTTTTATTGCAGACTTGAAGAGCTATTA;MAPQ=60;MATEID=3217824_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26239501_26264501_0C;SECONDARY;SPAN=4541;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:101 GQ:33.3 PL:[366.3, 33.3, 0.0] SR:97 DR:33 LR:-366.4 LO:366.4);ALT=A[chr7:26245987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26241497	+	chr7	26248008	+	.	11	0	3217826_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3217826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:26241497(+)-7:26248008(-)__7_26239501_26264501D;SPAN=6511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:82 GQ:14.3 PL:[14.3, 0.0, 182.6] SR:0 DR:11 LR:-14.1 LO:22.83);ALT=T[chr7:26248008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26245986	-	chr15	40854179	+	.	11	0	5931748_1	27.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=5931748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:26245986(-)-15:40854179(-)__15_40841501_40866501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:33 GQ:27.5 PL:[27.5, 0.0, 50.6] SR:0 DR:11 LR:-27.37 LO:27.81);ALT=[chr15:40854179[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	26246137	+	chr7	26248026	+	.	16	0	3217860_1	26.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=3217860_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:26246137(+)-7:26248026(-)__7_26239501_26264501D;SPAN=1889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:99 GQ:26 PL:[26.0, 0.0, 214.1] SR:0 DR:16 LR:-25.99 LO:34.61);ALT=A[chr7:26248026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26331706	+	chr7	26400593	+	ATTGATCGTGTCCTGTGCTGAAGATGTTTCCGGAACAACAGAAAG	12	14	3218505_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTGATCGTGTCCTGTGCTGAAGATGTTTCCGGAACAACAGAAAG;MAPQ=60;MATEID=3218505_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26386501_26411501_104C;SPAN=68887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:45 GQ:47.3 PL:[47.3, 0.0, 60.5] SR:14 DR:12 LR:-47.23 LO:47.34);ALT=C[chr7:26400593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26400681	+	chr7	26404155	+	.	0	7	3218566_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3218566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26386501_26411501_86C;SPAN=3474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:109 GQ:6.3 PL:[0.0, 6.3, 277.2] SR:7 DR:0 LR:6.424 LO:12.17);ALT=T[chr7:26404155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26404255	+	chr7	26411441	+	ACAACTGCCAGAACTTCCATCTAAAAACCTGTTTTTCAACATGAACAATCGCCAGCACGTGGATCAGCGTCGCCAGGGTCTGGAAGATTTCCTCAGAAA	0	16	3218576_1	24.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=ACAACTGCCAGAACTTCCATCTAAAAACCTGTTTTTCAACATGAACAATCGCCAGCACGTGGATCAGCGTCGCCAGGGTCTGGAAGATTTCCTCAGAAA;MAPQ=60;MATEID=3218576_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26386501_26411501_281C;SPAN=7186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:104 GQ:24.8 PL:[24.8, 0.0, 226.1] SR:16 DR:0 LR:-24.64 LO:34.24);ALT=T[chr7:26411441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26724469	+	chr7	26729903	+	.	2	4	3219679_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=3219679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26705001_26730001_341C;SPAN=5434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:102 GQ:7.5 PL:[0.0, 7.5, 260.7] SR:4 DR:2 LR:7.828 LO:10.2);ALT=T[chr7:26729903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26778499	+	chr7	26779506	+	.	0	4	3220037_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3220037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26754001_26779001_408C;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:45 GQ:1.1 PL:[1.1, 0.0, 106.7] SR:4 DR:0 LR:-1.012 LO:7.541);ALT=T[chr7:26779506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26883758	+	chr7	26903982	+	TTGTCTTGAAATTCCTGAAGATAGATAGACTTTACATCTTTTATCTTCTTAATAAGGGATTCTCTCTTTTCCTTTGCTTTCTTGGATAAATTTTCTCCTTTCAGTATATCTGCTACAAATGTTTCAACAT	2	27	3220299_1	79.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTGTCTTGAAATTCCTGAAGATAGATAGACTTTACATCTTTTATCTTCTTAATAAGGGATTCTCTCTTTTCCTTTGCTTTCTTGGATAAATTTTCTCCTTTCAGTATATCTGCTACAAATGTTTCAACAT;MAPQ=60;MATEID=3220299_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_26876501_26901501_108C;SPAN=20224;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:47 GQ:33.5 PL:[79.7, 0.0, 33.5] SR:27 DR:2 LR:-80.67 LO:80.67);ALT=T[chr7:26903982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	26894511	+	chr7	26903982	+	.	0	19	3220189_1	51.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3220189_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_26901001_26926001_366C;SPAN=9471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:42 GQ:48.2 PL:[51.5, 0.0, 48.2] SR:19 DR:0 LR:-51.34 LO:51.34);ALT=T[chr7:26903982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27136009	+	chr7	27139396	+	.	0	55	3220952_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=3220952_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27121501_27146501_293C;SPAN=3387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:128 GQ:99 PL:[146.9, 0.0, 163.4] SR:55 DR:0 LR:-146.9 LO:146.9);ALT=T[chr7:27139396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27203460	+	chr7	27204497	+	.	0	15	3221364_1	15.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3221364_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27195001_27220001_115C;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:127 GQ:15.2 PL:[15.2, 0.0, 292.4] SR:15 DR:0 LR:-15.11 LO:30.24);ALT=T[chr7:27204497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27211793	+	chr7	27212967	+	.	0	7	3221391_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=3221391_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27195001_27220001_109C;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:7 DR:0 LR:1.818 LO:12.7);ALT=C[chr7:27212967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27689253	+	chr7	27702317	+	.	0	7	3223270_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=3223270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27685001_27710001_54C;SPAN=13064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:114 GQ:7.5 PL:[0.0, 7.5, 290.4] SR:7 DR:0 LR:7.778 LO:12.03);ALT=C[chr7:27702317[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27779888	+	chr7	27788136	+	.	48	11	3224296_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3224296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27783001_27808001_516C;SPAN=8248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:11 DR:48 LR:-163.7 LO:163.7);ALT=G[chr7:27788136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27779904	+	chr7	27797647	+	.	13	0	3224297_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3224297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:27779904(+)-7:27797647(-)__7_27783001_27808001D;SPAN=17743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:0 DR:13 LR:-30.18 LO:31.58);ALT=G[chr7:27797647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27788307	+	chr7	27797648	+	.	0	28	3224320_1	65.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=3224320_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27783001_27808001_560C;SPAN=9341;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:98 GQ:65.9 PL:[65.9, 0.0, 171.5] SR:28 DR:0 LR:-65.88 LO:68.5);ALT=T[chr7:27797648[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	27797753	+	chr7	27805451	+	.	2	7	3224343_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3224343_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_27783001_27808001_419C;SPAN=7698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:110 GQ:0 PL:[0.0, 0.0, 267.3] SR:7 DR:2 LR:0.0927 LO:16.63);ALT=G[chr7:27805451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	28763949	+	chr7	28843815	+	.	3	3	3227086_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3227086_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_28836501_28861501_101C;SPAN=79866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:80 GQ:8.4 PL:[0.0, 8.4, 211.2] SR:3 DR:3 LR:8.47 LO:6.509);ALT=G[chr7:28843815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	28877819	+	chr7	139205859	-	.	14	0	3227218_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3227218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:28877819(+)-7:139205859(+)__7_28861001_28886001D;SPAN=110328040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:29 GQ:31.7 PL:[38.3, 0.0, 31.7] SR:0 DR:14 LR:-38.39 LO:38.39);ALT=A]chr7:139205859];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	29035500	+	chr7	29070190	+	.	5	13	3227845_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCT;MAPQ=60;MATEID=3227845_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_29057001_29082001_229C;SPAN=34690;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:55 GQ:44.6 PL:[44.6, 0.0, 87.5] SR:13 DR:5 LR:-44.52 LO:45.33);ALT=T[chr7:29070190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	29152440	+	chr7	29160508	+	.	2	5	3228241_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=3228241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_29130501_29155501_37C;SPAN=8068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:36 GQ:10.1 PL:[10.1, 0.0, 76.1] SR:5 DR:2 LR:-10.05 LO:13.07);ALT=T[chr7:29160508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	29160699	+	chr7	29185952	+	.	30	0	3228444_1	82.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3228444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:29160699(+)-7:29185952(-)__7_29179501_29204501D;SPAN=25253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:63 GQ:68.9 PL:[82.1, 0.0, 68.9] SR:0 DR:30 LR:-82.0 LO:82.0);ALT=A[chr7:29185952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	30538557	+	chr7	30544184	+	.	0	7	3233007_1	0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=3233007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_30527001_30552001_316C;SPAN=5627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:131 GQ:12 PL:[0.0, 12.0, 339.9] SR:7 DR:0 LR:12.38 LO:11.6);ALT=G[chr7:30544184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	30540299	+	chr7	30544184	+	.	0	31	3233018_1	65.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=3233018_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_30527001_30552001_107C;SPAN=3885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:135 GQ:65.9 PL:[65.9, 0.0, 260.6] SR:31 DR:0 LR:-65.76 LO:72.38);ALT=T[chr7:30544184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	30634760	+	chr7	30638410	+	.	0	8	3233409_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3233409_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_30625001_30650001_182C;SPAN=3650;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:8 DR:0 LR:3.123 LO:14.39);ALT=G[chr7:30638410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	31315559	+	chr7	31318954	+	.	90	41	3235743_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GGTGGCTCACGCCTGTAATCCCAGCACTTTGG;MAPQ=60;MATEID=3235743_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_7_31311001_31336001_78C;SPAN=3395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:93 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:41 DR:90 LR:-349.9 LO:349.9);ALT=G[chr7:31318954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32390165	+	chr7	32393113	+	.	78	40	3239179_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTGACTAATATAT;MAPQ=60;MATEID=3239179_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_32389001_32414001_54C;SPAN=2948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:38 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:40 DR:78 LR:-290.5 LO:290.5);ALT=T[chr7:32393113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32526950	+	chr7	32529930	+	.	36	0	3239537_1	80.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3239537_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:32526950(+)-7:32529930(-)__7_32511501_32536501D;SPAN=2980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:142 GQ:80.6 PL:[80.6, 0.0, 262.1] SR:0 DR:36 LR:-80.37 LO:85.85);ALT=G[chr7:32529930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32527369	+	chr7	32528861	+	ATATGGTACTGGAAGATGTCACTGAGTT	0	109	3239538_1	99.0	.	EVDNC=ASSMB;INSERTION=ATATGGTACTGGAAGATGTCACTGAGTT;MAPQ=60;MATEID=3239538_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_32511501_32536501_149C;SPAN=1492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:133 GQ:2.7 PL:[326.7, 2.7, 0.0] SR:109 DR:0 LR:-344.1 LO:344.1);ALT=A[chr7:32528861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	32527411	+	chr7	32529930	+	.	53	0	3239539_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3239539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:32527411(+)-7:32529930(-)__7_32511501_32536501D;SPAN=2519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:144 GQ:99 PL:[136.1, 0.0, 212.0] SR:0 DR:53 LR:-135.9 LO:136.9);ALT=A[chr7:32529930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	33075645	+	chr7	33102260	+	.	9	0	3242065_1	15.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3242065_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:33075645(+)-7:33102260(-)__7_33075001_33100001D;SPAN=26615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:0 DR:9 LR:-15.08 LO:19.6);ALT=G[chr7:33102260[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	35658574	+	chr11	122912044	+	.	9	43	5033027_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CACACACACACACACACACACACGCA;MAPQ=60;MATEID=5033027_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_122892001_122917001_226C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:84 GQ:63.2 PL:[139.1, 0.0, 63.2] SR:43 DR:9 LR:-140.5 LO:140.5);ALT=A[chr11:122912044[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	35840930	+	chr7	35872407	+	.	21	0	3251146_1	56.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3251146_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:35840930(+)-7:35872407(-)__7_35819001_35844001D;SPAN=31477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:46 GQ:53.6 PL:[56.9, 0.0, 53.6] SR:0 DR:21 LR:-56.86 LO:56.86);ALT=C[chr7:35872407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	36429653	+	chr7	36435873	+	.	0	7	3253160_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=3253160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_36431501_36456501_391C;SPAN=6220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:58 GQ:7.4 PL:[7.4, 0.0, 132.8] SR:7 DR:0 LR:-7.393 LO:14.18);ALT=G[chr7:36435873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	37354579	+	chr7	37382303	+	.	11	0	3256661_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3256661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:37354579(+)-7:37382303(-)__7_37362501_37387501D;SPAN=27724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:63 GQ:19.4 PL:[19.4, 0.0, 131.6] SR:0 DR:11 LR:-19.24 LO:24.2);ALT=T[chr7:37382303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	37355621	+	chr7	37382318	+	.	8	0	3256663_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3256663_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:37355621(+)-7:37382318(-)__7_37362501_37387501D;SPAN=26697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:0 DR:8 LR:-7.985 LO:16.11);ALT=A[chr7:37382318[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	37382369	+	chr7	37488276	+	.	0	10	3256753_1	22.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3256753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_37485001_37510001_201C;SPAN=105907;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:38 GQ:22.7 PL:[22.7, 0.0, 68.9] SR:10 DR:0 LR:-22.72 LO:24.04);ALT=T[chr7:37488276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	37723507	+	chr7	37725061	+	.	6	5	3257390_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3257390_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_37705501_37730501_382C;SPAN=1554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:477 GQ:99 PL:[0.0, 99.3, 1357.0] SR:5 DR:6 LR:99.52 LO:10.82);ALT=G[chr7:37725061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	37887805	+	chr7	37886731	+	.	18	0	3258031_1	45.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3258031_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:37886731(-)-7:37887805(+)__7_37877001_37902001D;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:51 GQ:45.8 PL:[45.8, 0.0, 75.5] SR:0 DR:18 LR:-45.6 LO:46.07);ALT=]chr7:37887805]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	38218024	+	chr7	38247045	+	.	70	13	3259293_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGGT;MAPQ=60;MATEID=3259293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38195501_38220501_359C;SPAN=29021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:64 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:13 DR:70 LR:-211.3 LO:211.3);ALT=T[chr7:38247045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38299832	+	chr7	38282029	+	.	3	8	3259558_1	13.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=C;MAPQ=57;MATEID=3259558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38293501_38318501_218C;SPAN=17803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:8 DR:3 LR:-13.55 LO:22.7);ALT=]chr7:38299832]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	38289174	+	chr7	38295938	+	.	41	6	3259379_1	99.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3259379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38269001_38294001_169C;SPAN=6764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:63 GQ:16.1 PL:[134.9, 0.0, 16.1] SR:6 DR:41 LR:-139.9 LO:139.9);ALT=C[chr7:38295938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38305280	+	chr7	38315860	+	.	30	37	3259626_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=C;MAPQ=52;MATEID=3259626_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38293501_38318501_23C;SPAN=10580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:129 GQ:99 PL:[146.6, 0.0, 166.4] SR:37 DR:30 LR:-146.6 LO:146.7);ALT=C[chr7:38315860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38381401	+	chr7	38389897	+	.	8	1	3259723_1	2.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3259723_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_7_38367001_38392001_477C;SECONDARY;SPAN=8496;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:1 DR:8 LR:-2.075 LO:16.94);ALT=G[chr7:38389897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38390051	+	chr7	38415156	+	.	24	14	3259775_1	82.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3259775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38367001_38392001_375C;SPAN=25105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:62 GQ:65.9 PL:[82.4, 0.0, 65.9] SR:14 DR:24 LR:-82.3 LO:82.3);ALT=G[chr7:38415156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38390051	+	chr7	38415722	+	.	5	3	3259776_1	6.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3259776_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38367001_38392001_149C;SPAN=25671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:62 GQ:6.5 PL:[6.5, 0.0, 141.8] SR:3 DR:5 LR:-6.31 LO:13.96);ALT=G[chr7:38415722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	38390052	+	chr7	38412964	+	.	15	19	3259777_1	72.0	.	DISC_MAPQ=23;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3259777_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_38367001_38392001_63C;SPAN=22912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:61 GQ:72.8 PL:[72.8, 0.0, 72.8] SR:19 DR:15 LR:-72.6 LO:72.6);ALT=G[chr7:38412964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	39606147	+	chr7	39610105	+	.	0	7	3263820_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3263820_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_39592001_39617001_41C;SPAN=3958;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:109 GQ:6.3 PL:[0.0, 6.3, 277.2] SR:7 DR:0 LR:6.424 LO:12.17);ALT=G[chr7:39610105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	39663424	+	chr7	39729979	+	ATTCTTCTTAATCCTTTGGTGAAAACTGAGACACAAAATGGCTGCAAATAAGCCCAAGGGTCAGAATTCTTTGGCTTTACACAAAGTCATCATGGTGGGCAGTGGTGGCGTGGGCAAGTCAGCTCTGACTCTACAGTTCATGTACGATG	0	21	3264395_1	55.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATTCTTCTTAATCCTTTGGTGAAAACTGAGACACAAAATGGCTGCAAATAAGCCCAAGGGTCAGAATTCTTTGGCTTTACACAAAGTCATCATGGTGGGCAGTGGTGGCGTGGGCAAGTCAGCTCTGACTCTACAGTTCATGTACGATG;MAPQ=60;MATEID=3264395_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_39714501_39739501_21C;SPAN=66555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:53 GQ:55.1 PL:[55.1, 0.0, 71.6] SR:21 DR:0 LR:-54.96 LO:55.11);ALT=G[chr7:39729979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	39663424	+	chr7	39726228	+	.	11	14	3264045_1	55.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3264045_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_39641001_39666001_239C;SPAN=62804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:28 GQ:12.2 PL:[55.1, 0.0, 12.2] SR:14 DR:11 LR:-56.61 LO:56.61);ALT=G[chr7:39726228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	39726380	+	chr7	39729979	+	.	2	7	3264435_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3264435_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_7_39714501_39739501_21C;SPAN=3599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:104 GQ:1.5 PL:[0.0, 1.5, 254.1] SR:7 DR:2 LR:1.768 LO:14.56);ALT=G[chr7:39729979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42964398	+	chr7	42966135	+	.	3	121	3275342_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3275342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_42948501_42973501_166C;SPAN=1737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:146 GQ:16.3 PL:[386.1, 16.3, 0.0] SR:121 DR:3 LR:-396.9 LO:396.9);ALT=T[chr7:42966135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42964437	+	chr7	42971715	+	.	55	0	3275343_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3275343_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:42964437(+)-7:42971715(-)__7_42948501_42973501D;SPAN=7278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:159 GQ:99 PL:[138.5, 0.0, 247.4] SR:0 DR:55 LR:-138.5 LO:140.2);ALT=T[chr7:42971715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42966297	+	chr7	42971716	+	.	133	0	3275350_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=3275350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:42966297(+)-7:42971716(-)__7_42948501_42973501D;SPAN=5419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:152 GQ:31 PL:[429.1, 31.0, 0.0] SR:0 DR:133 LR:-431.5 LO:431.5);ALT=T[chr7:42971716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	42972116	+	chr7	42974553	+	.	9	8	3275378_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3275378_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_42948501_42973501_162C;SPAN=2437;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:8 DR:9 LR:-44.2 LO:44.37);ALT=G[chr7:42974553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	43684998	+	chr7	43687134	+	.	0	17	3277973_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3277973_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_43683501_43708501_63C;SPAN=2136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:120 GQ:23.6 PL:[23.6, 0.0, 267.8] SR:17 DR:0 LR:-23.61 LO:35.71);ALT=T[chr7:43687134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	43687276	+	chr7	43769025	+	.	21	0	3278181_1	52.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3278181_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:43687276(+)-7:43769025(-)__7_43757001_43782001D;SPAN=81749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:63 GQ:52.4 PL:[52.4, 0.0, 98.6] SR:0 DR:21 LR:-52.25 LO:53.09);ALT=T[chr7:43769025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	43906584	+	chr7	43908560	+	.	0	75	3278796_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=3278796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_43904001_43929001_27C;SPAN=1976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:165 GQ:99 PL:[203.0, 0.0, 196.4] SR:75 DR:0 LR:-202.9 LO:202.9);ALT=G[chr7:43908560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	43906631	+	chr7	43908906	+	.	78	0	3278797_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3278797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:43906631(+)-7:43908906(-)__7_43904001_43929001D;SPAN=2275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:119 GQ:63.5 PL:[225.2, 0.0, 63.5] SR:0 DR:78 LR:-230.3 LO:230.3);ALT=C[chr7:43908906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44084393	+	chr7	44092464	+	.	11	0	3280109_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3280109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44084393(+)-7:44092464(-)__7_44075501_44100501D;SPAN=8071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:117 GQ:4.7 PL:[4.7, 0.0, 278.6] SR:0 DR:11 LR:-4.613 LO:21.02);ALT=G[chr7:44092464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44084420	+	chr7	44089823	+	.	16	18	3280110_1	23.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3280110_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CTCTCT;SCTG=c_7_44075501_44100501_437C;SPAN=5403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:125 GQ:23.6 PL:[23.6, 0.0, 200.4] SR:18 DR:16 LR:-23.38 LO:33.17);ALT=G[chr7:44089823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44084420	+	chr7	44091428	+	GCTCTCTTTACCTATGAAGGCAACAGCAATGACATCCGCGTGGCTGGCACAGGG	65	56	3280111_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GCTCTCTTTACCTATGAAGGCAACAGCAATGACATCCGCGTGGCTGGCACAGGG;MAPQ=60;MATEID=3280111_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_7_44075501_44100501_437C;SPAN=7008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:134 GQ:56.3 PL:[267.5, 0.0, 56.3] SR:56 DR:65 LR:-275.0 LO:275.0);ALT=G[chr7:44091428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44092541	+	chr7	44096354	+	.	0	11	3280140_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3280140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_44075501_44100501_19C;SPAN=3813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:137 GQ:0.6 PL:[0.0, 0.6, 333.3] SR:11 DR:0 LR:0.8057 LO:20.23);ALT=G[chr7:44096354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44120518	+	chr7	44121850	+	.	0	12	3279514_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=3279514_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_44100001_44125001_32C;SPAN=1332;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:106 GQ:11 PL:[11.0, 0.0, 245.3] SR:12 DR:0 LR:-10.89 LO:23.95);ALT=G[chr7:44121850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44157664	+	chr7	44161432	+	.	0	10	3279970_1	5.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=3279970_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_7_44149001_44174001_98C;SPAN=3768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:102 GQ:5.6 PL:[5.6, 0.0, 239.9] SR:10 DR:0 LR:-5.376 LO:19.3);ALT=C[chr7:44161432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44646277	+	chr7	44663946	+	.	11	0	3282074_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3282074_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44646277(+)-7:44663946(-)__7_44663501_44688501D;SPAN=17669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:53 GQ:22.1 PL:[22.1, 0.0, 104.6] SR:0 DR:11 LR:-21.95 LO:25.13);ALT=C[chr7:44663946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44875303	+	chr7	44887566	+	.	21	0	3283040_1	53.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=3283040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44875303(+)-7:44887566(-)__7_44859501_44884501D;SPAN=12263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:59 GQ:53.3 PL:[53.3, 0.0, 89.6] SR:0 DR:21 LR:-53.34 LO:53.85);ALT=C[chr7:44887566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	44880622	+	chr7	44887566	+	.	52	0	3283069_1	99.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=3283069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44880622(+)-7:44887566(-)__7_44859501_44884501D;SPAN=6944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:58 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:52 LR:-171.1 LO:171.1);ALT=G[chr7:44887566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93277465	+	chr7	44887593	+	.	73	0	6038799_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6038799_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:44887593(-)-15:93277465(+)__15_93271501_93296501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:92 GQ:5 PL:[216.2, 0.0, 5.0] SR:0 DR:73 LR:-227.9 LO:227.9);ALT=]chr15:93277465]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	45016673	+	chr7	45018464	+	.	45	21	3283667_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=3283667_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_45006501_45031501_206C;SPAN=1791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:119 GQ:99 PL:[139.4, 0.0, 149.3] SR:21 DR:45 LR:-139.4 LO:139.4);ALT=G[chr7:45018464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	45023645	+	chr7	45026122	+	AAGACTGCTTGAACATGAGACTCAAGGAGGGACCTCAGCAGGCCTGGGGTGTTCAGCAACTATTCCTGGCCGGGGCATCTTGCAAAGGAGTTGCTGTGACAGTAAGCTCTTCCACTTTGAGACCGTCACCTCAGCCACGGCTCCC	24	63	3283704_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=AAGACTGCTTGAACATGAGACTCAAGGAGGGACCTCAGCAGGCCTGGGGTGTTCAGCAACTATTCCTGGCCGGGGCATCTTGCAAAGGAGTTGCTGTGACAGTAAGCTCTTCCACTTTGAGACCGTCACCTCAGCCACGGCTCCC;MAPQ=60;MATEID=3283704_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_45006501_45031501_212C;SPAN=2477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:74 DP:122 GQ:82.7 PL:[211.4, 0.0, 82.7] SR:63 DR:24 LR:-214.2 LO:214.2);ALT=A[chr7:45026122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	45024073	+	chr7	45026145	+	.	35	0	3283706_1	83.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3283706_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:45024073(+)-7:45026145(-)__7_45006501_45031501D;SPAN=2072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:119 GQ:83.3 PL:[83.3, 0.0, 205.4] SR:0 DR:35 LR:-83.3 LO:86.15);ALT=C[chr7:45026145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	45119670	+	chr7	45118629	+	.	12	0	3284241_1	11.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=3284241_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:45118629(-)-7:45119670(+)__7_45104501_45129501D;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:103 GQ:11.9 PL:[11.9, 0.0, 236.3] SR:0 DR:12 LR:-11.71 LO:24.11);ALT=]chr7:45119670]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	45148827	+	chr7	45151240	+	.	13	0	3284166_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3284166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:45148827(+)-7:45151240(-)__7_45129001_45154001D;SPAN=2413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:116 GQ:11.6 PL:[11.6, 0.0, 269.0] SR:0 DR:13 LR:-11.49 LO:25.89);ALT=G[chr7:45151240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	47603707	-	chr7	47604840	+	.	8	0	3292797_1	0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=3292797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:47603707(-)-7:47604840(-)__7_47603501_47628501D;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:0 DR:8 LR:-0.6702 LO:14.89);ALT=[chr7:47604840[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	48129962	+	chr7	48134359	+	.	0	9	3295020_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3295020_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_48118001_48143001_181C;SPAN=4397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:151 GQ:10.9 PL:[0.0, 10.9, 386.1] SR:9 DR:0 LR:11.2 LO:15.35);ALT=G[chr7:48134359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	61741164	+	chr7	61739964	+	.	9	0	3334997_1	0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3334997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:61739964(-)-7:61741164(+)__7_61740001_61765001D;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:125 GQ:3.9 PL:[0.0, 3.9, 310.2] SR:0 DR:9 LR:4.157 LO:16.11);ALT=]chr7:61741164]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	61751825	+	chr7	61750825	+	.	12	0	3335070_1	4.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=3335070_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:61750825(-)-7:61751825(+)__7_61740001_61765001D;SPAN=1000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:132 GQ:4.1 PL:[4.1, 0.0, 314.3] SR:0 DR:12 LR:-3.85 LO:22.75);ALT=]chr7:61751825]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	61786098	+	chr7	61780169	+	.	9	0	3334839_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=3334839_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:61780169(-)-7:61786098(+)__7_61764501_61789501D;SPAN=5929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:137 GQ:7.2 PL:[0.0, 7.2, 346.5] SR:0 DR:9 LR:7.408 LO:15.74);ALT=]chr7:61786098]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	61848994	+	chr7	61857679	+	CAAATAT	53	48	3333354_1	99.0	.	DISC_MAPQ=12;EVDNC=ASDIS;INSERTION=CAAATAT;MAPQ=47;MATEID=3333354_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_7_61838001_61863001_89C;SPAN=8685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:144 GQ:93.2 PL:[254.9, 0.0, 93.2] SR:48 DR:53 LR:-258.8 LO:258.8);ALT=C[chr7:61857679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	62002310	+	chr7	62004852	+	.	89	35	3333854_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TTTCTTTTGATAGAACAGTTTTGAAACACTCTTT;MAPQ=60;MATEID=3333854_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_61985001_62010001_172C;SPAN=2542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:26 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:35 DR:89 LR:-326.8 LO:326.8);ALT=T[chr7:62004852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55239304	+	chr7	62079588	+	CAGCTAGAATGAGTACCATG	7	58	3334450_1	99.0	.	DISC_MAPQ=5;EVDNC=TSI_L;HOMSEQ=TGGTGCAATCTCGGCTCACTGCAACCTCTG;INSERTION=CAGCTAGAATGAGTACCATG;MAPQ=60;MATEID=3334450_2;MATENM=0;NM=2;NUMPARTS=3;REPSEQ=TT;SCTG=c_7_62058501_62083501_150C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:48 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:58 DR:7 LR:-178.2 LO:178.2);ALT=]chr20:55239304]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	62354260	+	chr7	62355446	-	.	13	0	3335353_1	36.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3335353_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:62354260(+)-7:62355446(+)__7_62328001_62353001D;SPAN=1186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:13 DP:0 GQ:3.3 PL:[36.3, 3.3, 0.0] SR:0 DR:13 LR:-36.31 LO:36.31);ALT=G]chr7:62355446];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	67427921	+	chr7	63296509	+	.	24	82	3360964_1	99.0	.	DISC_MAPQ=41;EVDNC=TSI_L;MAPQ=60;MATEID=3360964_2;MATENM=3;NM=1;NUMPARTS=3;SCTG=c_7_67424001_67449001_465C;SPAN=4131412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:37 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:82 DR:24 LR:-277.3 LO:277.3);ALT=]chr7:67427921]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	63774532	+	chr7	63796636	+	.	5	4	3342295_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3342295_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_7_63773501_63798501_175C;SECONDARY;SPAN=22104;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:108 GQ:6 PL:[0.0, 6.0, 273.9] SR:4 DR:5 LR:6.153 LO:12.2);ALT=G[chr7:63796636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64315824	+	chr7	64318059	+	.	84	38	3344483_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGAATTTTATTTTATC;MAPQ=60;MATEID=3344483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_64312501_64337501_113C;SPAN=2235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:30 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:38 DR:84 LR:-300.4 LO:300.4);ALT=C[chr7:64318059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64465573	+	chr7	64466919	+	.	0	6	3345326_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=3345326_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_64459501_64484501_103C;SPAN=1346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:116 GQ:11.4 PL:[0.0, 11.4, 303.6] SR:6 DR:0 LR:11.62 LO:9.853);ALT=C[chr7:64466919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	64754604	-	chr7	64755984	+	.	9	0	3346725_1	2.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3346725_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:64754604(-)-7:64755984(-)__7_64753501_64778501D;SPAN=1380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:101 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.346 LO:16.98);ALT=[chr7:64755984[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	65441190	+	chr7	65444385	+	.	3	3	3350671_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=3350671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65439501_65464501_223C;SPAN=3195;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:3 DR:3 LR:5.711 LO:8.577);ALT=C[chr7:65444385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	65445398	+	chr7	65446961	+	.	0	37	3350684_1	92.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3350684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65439501_65464501_118C;SPAN=1563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:112 GQ:92 PL:[92.0, 0.0, 177.8] SR:37 DR:0 LR:-91.79 LO:93.37);ALT=T[chr7:65446961[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	65541080	+	chr7	65546788	+	.	18	12	3351155_1	56.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3351155_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65537501_65562501_312C;SPAN=5708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:108 GQ:56.6 PL:[56.6, 0.0, 205.1] SR:12 DR:18 LR:-56.57 LO:61.32);ALT=G[chr7:65546788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	65579956	+	chr7	65595728	+	.	8	0	3351581_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3351581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:65579956(+)-7:65595728(-)__7_65562001_65587001D;SPAN=15772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=G[chr7:65595728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	65589705	+	chr7	65591966	+	.	42	42	3351273_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=3351273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_65586501_65611501_276C;SPAN=2261;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:74 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:42 DR:42 LR:-217.9 LO:217.9);ALT=C[chr7:65591966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66030576	+	chr7	66258667	-	ACCTGCT	39	29	3353859_1	99.0	.	DISC_MAPQ=32;EVDNC=TSI_L;INSERTION=ACCTGCT;MAPQ=60;MATEID=3353859_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_7_66027501_66052501_45C;SPAN=228091;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:77 GQ:5.6 PL:[180.5, 0.0, 5.6] SR:29 DR:39 LR:-190.3 LO:190.3);ALT=C]chr7:66258667];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	73382119	+	chr7	66193573	+	.	21	52	3386451_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CTCCAC;MAPQ=60;MATEID=3386451_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_73377501_73402501_345C;SPAN=7188546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:60 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:52 DR:21 LR:-208.0 LO:208.0);ALT=]chr7:73382119]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	66258674	-	chr7	75740180	+	.	8	0	3400572_1	12.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3400572_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:66258674(-)-7:75740180(-)__7_75729501_75754501D;SPAN=9481506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=[chr7:75740180[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	66386451	+	chr7	66406834	+	.	0	11	3355223_1	20.0	.	EVDNC=ASSMB;HOMSEQ=GGTG;MAPQ=60;MATEID=3355223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_66395001_66420001_224C;SPAN=20383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:11 DR:0 LR:-20.87 LO:24.74);ALT=G[chr7:66406834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66611102	-	chr7	72130619	+	.	8	0	3356682_1	12.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3356682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:66611102(-)-7:72130619(-)__7_66591001_66616001D;SPAN=5519517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=[chr7:72130619[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	66633029	+	chr7	72109304	-	.	11	0	3356525_1	20.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=3356525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:66633029(+)-7:72109304(+)__7_66615501_66640501D;SPAN=5476275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:61 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-19.78 LO:24.38);ALT=A]chr7:72109304];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	66697505	+	chr7	66699292	+	.	45	18	3356890_1	99.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCCAGCCTGGG;MAPQ=60;MATEID=3356890_2;MATENM=0;NM=2;NUMPARTS=2;REPSEQ=GGG;SCTG=c_7_66689001_66714001_393C;SECONDARY;SPAN=1787;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:80 GQ:21.2 PL:[173.0, 0.0, 21.2] SR:18 DR:45 LR:-180.0 LO:180.0);ALT=G[chr7:66699292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	66764413	+	chr7	66767363	+	.	9	3	3357507_1	7.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=21;MATEID=3357507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_66762501_66787501_349C;SPAN=2950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:96 GQ:7.1 PL:[7.1, 0.0, 224.9] SR:3 DR:9 LR:-7.001 LO:19.58);ALT=T[chr7:66767363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	70420969	+	chr7	70438887	-	.	5	42	3372270_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=3372270_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_7_70437501_70462501_182C;SPAN=17918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:48 GQ:9.6 PL:[135.3, 9.6, 0.0] SR:42 DR:5 LR:-136.3 LO:136.3);ALT=C]chr7:70438887];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	70426185	-	chr7	70438880	+	.	41	43	3372272_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=3372272_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_70437501_70462501_158C;SPAN=12695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:48 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:43 DR:41 LR:-224.5 LO:224.5);ALT=[chr7:70438880[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	70622462	+	chr9	16896157	+	ACGAAACCCCATCTCTACAAAAAATACAAAAATTAGCCAGGCGTGGTG	5	68	4146471_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_L;INSERTION=ACGAAACCCCATCTCTACAAAAAATACAAAAATTAGCCAGGCGTGGTG;MAPQ=60;MATEID=4146471_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_9_16880501_16905501_46C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:8 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:68 DR:5 LR:-214.6 LO:214.6);ALT=G[chr9:16896157[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	71211913	+	chr7	71212956	+	.	51	32	3375663_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAAA;MAPQ=60;MATEID=3375663_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_71197001_71222001_193C;SPAN=1043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:67 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:32 DR:51 LR:-208.0 LO:208.0);ALT=A[chr7:71212956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	71983058	-	chr7	71984269	+	.	8	0	3378425_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=3378425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:71983058(-)-7:71984269(-)__7_71981001_72006001D;SPAN=1211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:108 GQ:2.7 PL:[0.0, 2.7, 267.3] SR:0 DR:8 LR:2.852 LO:14.42);ALT=[chr7:71984269[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	102009660	+	chr7	72355105	+	TATATATATATTTGCTAT	3	7	3380323_1	21.0	.	DISC_MAPQ=5;EVDNC=ASDIS;INSERTION=TATATATATATTTGCTAT;MAPQ=26;MATEID=3380323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_72348501_72373501_301C;SPAN=29654555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:7 DR:3 LR:-21.63 LO:23.53);ALT=]chr7:102009660]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	72966573	+	chr7	72971816	+	.	0	9	3384222_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=3384222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_72961001_72986001_386C;SPAN=5243;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:9 DR:0 LR:-8.577 LO:18.05);ALT=C[chr7:72971816[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73098035	+	chr7	73101146	+	.	16	0	3385188_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3385188_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:73098035(+)-7:73101146(-)__7_73083501_73108501D;SPAN=3111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:136 GQ:16.1 PL:[16.1, 0.0, 313.1] SR:0 DR:16 LR:-15.97 LO:32.22);ALT=C[chr7:73101146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73468108	+	chr8	41187845	+	.	2	16	3834211_1	29.0	.	DISC_MAPQ=11;EVDNC=ASDIS;HOMSEQ=TGGATGGATGGATGGATGGATG;MAPQ=31;MATEID=3834211_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_41184501_41209501_64C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:101 GQ:29 PL:[29.0, 0.0, 213.8] SR:16 DR:2 LR:-28.75 LO:37.11);ALT=G[chr8:41187845[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	73549766	+	chr7	73550967	+	.	34	45	3387402_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTGAGA;MAPQ=60;MATEID=3387402_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_73549001_73574001_217C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:26 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:45 DR:34 LR:-204.7 LO:204.7);ALT=A[chr7:73550967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73624418	+	chr7	73629150	+	.	74	7	3387642_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3387642_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_73622501_73647501_218C;SPAN=4732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:109 GQ:39.8 PL:[224.6, 0.0, 39.8] SR:7 DR:74 LR:-232.0 LO:232.0);ALT=G[chr7:73629150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73624418	+	chr7	73630273	+	.	29	3	3387643_1	68.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=3387643_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_73622501_73647501_178C;SPAN=5855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:124 GQ:68.9 PL:[68.9, 0.0, 230.6] SR:3 DR:29 LR:-68.74 LO:73.71);ALT=G[chr7:73630273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73624431	+	chr7	73634073	+	.	8	0	3387644_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3387644_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:73624431(+)-7:73634073(-)__7_73622501_73647501D;SPAN=9642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:132 GQ:9 PL:[0.0, 9.0, 336.6] SR:0 DR:8 LR:9.354 LO:13.7);ALT=C[chr7:73634073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73624449	+	chr7	73631151	+	.	14	0	3387646_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3387646_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:73624449(+)-7:73631151(-)__7_73622501_73647501D;SPAN=6702;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:138 GQ:8.9 PL:[8.9, 0.0, 325.7] SR:0 DR:14 LR:-8.826 LO:27.24);ALT=C[chr7:73631151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73629270	+	chr7	73630276	+	.	2	13	3387658_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3387658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_73622501_73647501_101C;SPAN=1006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:136 GQ:12.8 PL:[12.8, 0.0, 316.4] SR:13 DR:2 LR:-12.67 LO:29.76);ALT=G[chr7:73630276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73663449	+	chr7	73668600	+	GCAATGATGATGTTGGGCACATTTCCTTCCCTTGCAAAGACCTCTAGCCTGCTCACGGTGTCTTCATTCCCGACAATTTCATTCAGCTTTACTGGCCTATATTTTTCAAC	0	22	3387943_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GCAATGATGATGTTGGGCACATTTCCTTCCCTTGCAAAGACCTCTAGCCTGCTCACGGTGTCTTCATTCCCGACAATTTCATTCAGCTTTACTGGCCTATATTTTTCAAC;MAPQ=60;MATEID=3387943_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_73647001_73672001_169C;SPAN=5151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:128 GQ:38 PL:[38.0, 0.0, 272.3] SR:22 DR:0 LR:-37.94 LO:48.24);ALT=C[chr7:73668600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73664167	+	chr7	73668634	+	.	9	0	3387951_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3387951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:73664167(+)-7:73668634(-)__7_73647001_73672001D;SPAN=4467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:119 GQ:2.4 PL:[0.0, 2.4, 293.7] SR:0 DR:9 LR:2.531 LO:16.31);ALT=A[chr7:73668634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	73666874	+	chr7	73668656	+	.	12	0	3387966_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3387966_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:73666874(+)-7:73668656(-)__7_73647001_73672001D;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:115 GQ:8.6 PL:[8.6, 0.0, 269.3] SR:0 DR:12 LR:-8.456 LO:23.5);ALT=T[chr7:73668656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	74072395	+	chr7	74103457	+	.	0	12	3389840_1	33.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3389840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_74063501_74088501_304C;SPAN=31062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:24 GQ:23.3 PL:[33.2, 0.0, 23.3] SR:12 DR:0 LR:-33.17 LO:33.17);ALT=G[chr7:74103457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	74103561	+	chr7	74105304	+	.	0	12	3389745_1	8.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3389745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_74088001_74113001_324C;SPAN=1743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:117 GQ:8 PL:[8.0, 0.0, 275.3] SR:12 DR:0 LR:-7.914 LO:23.41);ALT=G[chr7:74105304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75221832	+	chr7	75228502	+	.	0	19	3397323_1	30.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3397323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75215001_75240001_12C;SPAN=6670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:118 GQ:30.8 PL:[30.8, 0.0, 255.2] SR:19 DR:0 LR:-30.75 LO:41.07);ALT=G[chr7:75228502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75221878	+	chr7	75268437	+	.	10	0	3397919_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3397919_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:75221878(+)-7:75268437(-)__7_75264001_75289001D;SPAN=46559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:33 GQ:24.2 PL:[24.2, 0.0, 53.9] SR:0 DR:10 LR:-24.07 LO:24.77);ALT=T[chr7:75268437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75363121	+	chr7	75368118	+	.	55	21	3398591_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=3398591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75362001_75387001_343C;SPAN=4997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:137 GQ:99 PL:[174.2, 0.0, 157.7] SR:21 DR:55 LR:-174.2 LO:174.2);ALT=G[chr7:75368118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75651313	+	chr7	75659739	+	CTTCACTCGAAGGGCAGTGATCACATGGCTTTCGTCATACTCCCATTTGGAACGGACAT	3	14	3400337_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTTCACTCGAAGGGCAGTGATCACATGGCTTTCGTCATACTCCCATTTGGAACGGACAT;MAPQ=60;MATEID=3400337_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_7_75656001_75681001_244C;SPAN=8426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:47 GQ:43.4 PL:[43.4, 0.0, 69.8] SR:14 DR:3 LR:-43.38 LO:43.74);ALT=T[chr7:75659739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75658069	+	chr7	75677064	+	.	9	0	3400352_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3400352_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:75658069(+)-7:75677064(-)__7_75656001_75681001D;SPAN=18995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:122 GQ:3 PL:[0.0, 3.0, 300.3] SR:0 DR:9 LR:3.344 LO:16.21);ALT=A[chr7:75677064[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75659849	+	chr7	75677130	+	.	17	11	3400364_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=3400364_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_75656001_75681001_315C;SPAN=17281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:127 GQ:41.6 PL:[41.6, 0.0, 266.0] SR:11 DR:17 LR:-41.52 LO:51.01);ALT=G[chr7:75677130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75677544	+	chr7	75684146	+	.	110	54	3400448_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3400448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75656001_75681001_239C;SPAN=6602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:47 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:54 DR:110 LR:-412.6 LO:412.6);ALT=G[chr7:75684146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75677586	+	chr7	75686725	+	.	24	0	3400451_1	79.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3400451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:75677586(+)-7:75686725(-)__7_75656001_75681001D;SPAN=9139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:27 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:0 DR:24 LR:-78.52 LO:78.52);ALT=G[chr7:75686725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75684317	+	chr7	75686726	+	.	0	66	3399826_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3399826_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75680501_75705501_220C;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:143 GQ:99 PL:[179.3, 0.0, 166.1] SR:66 DR:0 LR:-179.1 LO:179.1);ALT=G[chr7:75686726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75687398	+	chr7	75689690	+	.	4	11	3399839_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=3399839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75680501_75705501_130C;SPAN=2292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:114 GQ:12.2 PL:[12.2, 0.0, 263.0] SR:11 DR:4 LR:-12.03 LO:25.99);ALT=T[chr7:75689690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75689817	+	chr7	75693654	+	GTTTGGATCCAGCTCGAGTCAACGTCCCTGTCATTGGTGGCCATGCTGGGAAGACCATCATCCCCCTGATCTCT	0	12	3399849_1	7.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=GTTTGGATCCAGCTCGAGTCAACGTCCCTGTCATTGGTGGCCATGCTGGGAAGACCATCATCCCCCTGATCTCT;MAPQ=60;MATEID=3399849_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_75680501_75705501_206C;SPAN=3837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:121 GQ:7.1 PL:[7.1, 0.0, 284.3] SR:12 DR:0 LR:-6.83 LO:23.22);ALT=G[chr7:75693654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75689817	+	chr7	75692831	+	.	4	7	3399848_1	1.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=3399848_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_7_75680501_75705501_206C;SPAN=3014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:117 GQ:1.4 PL:[1.4, 0.0, 281.9] SR:7 DR:4 LR:-1.312 LO:18.67);ALT=G[chr7:75692831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75694271	+	chr7	75695596	+	.	5	20	3399872_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3399872_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75680501_75705501_355C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:111 GQ:39.5 PL:[39.5, 0.0, 227.6] SR:20 DR:5 LR:-39.25 LO:47.02);ALT=G[chr7:75695596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	75959550	+	chr7	75988035	+	.	6	11	3401578_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAC;MAPQ=60;MATEID=3401578_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_75950001_75975001_286C;SPAN=28485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:49 GQ:32.9 PL:[32.9, 0.0, 85.7] SR:11 DR:6 LR:-32.94 LO:34.25);ALT=C[chr7:75988035[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	76903688	+	chr7	76906830	+	.	0	7	3406444_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CCTGT;MAPQ=60;MATEID=3406444_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_76881001_76906001_65C;SPAN=3142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:7 DR:0 LR:-9.832 LO:14.73);ALT=T[chr7:76906830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	77423767	+	chr7	77427624	+	.	13	0	3408190_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3408190_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:77423767(+)-7:77427624(-)__7_77420001_77445001D;SPAN=3857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:121 GQ:10.4 PL:[10.4, 0.0, 281.0] SR:0 DR:13 LR:-10.13 LO:25.64);ALT=T[chr7:77427624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	77428283	+	chr7	77522922	+	.	8	0	3409027_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3409027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:77428283(+)-7:77522922(-)__7_77518001_77543001D;SPAN=94639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=C[chr7:77522922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	77428288	+	chr7	77469537	+	.	11	13	3408765_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3408765_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_77469001_77494001_197C;SPAN=41249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:43 GQ:41.3 PL:[41.3, 0.0, 61.1] SR:13 DR:11 LR:-41.17 LO:41.42);ALT=G[chr7:77469537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	77981839	+	chr7	78082249	+	A	25	13	3411044_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=3411044_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_78081501_78106501_76C;SPAN=100410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:31 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:13 DR:25 LR:-89.12 LO:89.12);ALT=C[chr7:78082249[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	78124664	-	chr7	78125927	+	GC	3	3	3411025_1	0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=GC;MAPQ=50;MATEID=3411025_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_78106001_78131001_213C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:99 GQ:10.2 PL:[0.0, 10.2, 260.7] SR:3 DR:3 LR:10.32 LO:8.158);ALT=[chr7:78125927[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	78190207	+	chr7	78257685	+	.	25	16	3411274_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=3411274_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_78253001_78278001_116C;SPAN=67478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:31 GQ:9 PL:[99.0, 9.0, 0.0] SR:16 DR:25 LR:-99.02 LO:99.02);ALT=C[chr7:78257685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80268062	+	chr7	80275402	+	.	61	22	3417511_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3417511_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_80262001_80287001_273C;SPAN=7340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:134 GQ:86 PL:[237.8, 0.0, 86.0] SR:22 DR:61 LR:-241.5 LO:241.5);ALT=G[chr7:80275402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80276176	+	chr7	80285854	+	.	8	11	3417545_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3417545_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_7_80262001_80287001_212C;SPAN=9678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:116 GQ:18.2 PL:[18.2, 0.0, 262.4] SR:11 DR:8 LR:-18.09 LO:30.87);ALT=G[chr7:80285854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80286016	+	chr7	80290377	+	.	22	12	3417376_1	65.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3417376_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_80286501_80311501_318C;SPAN=4361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:75 GQ:65.6 PL:[65.6, 0.0, 115.1] SR:12 DR:22 LR:-65.51 LO:66.29);ALT=G[chr7:80290377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80290527	+	chr7	80292306	+	.	0	29	3417612_1	85.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3417612_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_80262001_80287001_337C;SPAN=1779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:0 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:29 DR:0 LR:-85.82 LO:85.82);ALT=G[chr7:80292306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80290527	+	chr7	80293722	+	CTGCATCCCATATCTATCAAAATCAATTTGTTCAAATGATCCTCAATTCACTTATTAACAAGTCAAAATCTTCTATGTTCCAAGTCAGAACTTTGAGAGAACTGTTATGGGGCTATAGGGATCCATTTTTGAGTTTGGTTCCGTACCCTGTTACTACCACAGTTGGTCTGTTTTATCCT	2	35	3417393_1	90.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTGCATCCCATATCTATCAAAATCAATTTGTTCAAATGATCCTCAATTCACTTATTAACAAGTCAAAATCTTCTATGTTCCAAGTCAGAACTTTGAGAGAACTGTTATGGGGCTATAGGGATCCATTTTTGAGTTTGGTTCCGTACCCTGTTACTACCACAGTTGGTCTGTTTTATCCT;MAPQ=60;MATEID=3417393_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_80286501_80311501_62C;SPAN=3195;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:116 GQ:90.8 PL:[90.8, 0.0, 189.8] SR:35 DR:2 LR:-90.71 LO:92.67);ALT=G[chr7:80293722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80292485	+	chr7	80293722	+	.	5	5	3417398_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3417398_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ACAACA;SCTG=c_7_80286501_80311501_62C;SPAN=1237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:101 GQ:0.9 PL:[0.0, 0.9, 182.0] SR:5 DR:5 LR:1.343 LO:12.42);ALT=T[chr7:80293722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80293814	+	chr7	80299265	+	AATCTGTCCTATTGGGAAAGTCACTGCGACATGATTAATGGT	2	22	3417405_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACAG;INSERTION=AATCTGTCCTATTGGGAAAGTCACTGCGACATGATTAATGGT;MAPQ=60;MATEID=3417405_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_80286501_80311501_245C;SPAN=5451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:124 GQ:45.8 PL:[45.8, 0.0, 253.7] SR:22 DR:2 LR:-45.63 LO:54.01);ALT=G[chr7:80299265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80301407	+	chr7	80303296	+	.	12	0	3417441_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3417441_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:80301407(+)-7:80303296(-)__7_80286501_80311501D;SPAN=1889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:110 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:0 DR:12 LR:-9.81 LO:23.75);ALT=A[chr7:80303296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	80303463	+	chr7	80305700	+	.	11	7	3417448_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3417448_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_80286501_80311501_267C;SPAN=2237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:117 GQ:17.9 PL:[17.9, 0.0, 265.4] SR:7 DR:11 LR:-17.82 LO:30.81);ALT=A[chr7:80305700[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	81789164	+	chr10	60902930	-	.	84	47	3422222_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=3422222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_81781001_81806001_162C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:43 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:47 DR:84 LR:-326.8 LO:326.8);ALT=T]chr10:60902930];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	83929121	+	chr22	24077834	-	.	9	70	3429035_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3429035_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_83912501_83937501_4C;SECONDARY;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:28 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:70 DR:9 LR:-217.9 LO:217.9);ALT=A]chr22:24077834];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	83929122	-	chr22	24077747	+	.	17	61	3429037_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GATCACCTGAGGTCAGGAGTTTGAGACCAGCCTG;MAPQ=8;MATEID=3429037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_83912501_83937501_78C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:27 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:61 DR:17 LR:-227.8 LO:227.8);ALT=[chr22:24077747[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	86954760	+	chr7	86970839	+	.	0	16	3437623_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3437623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_86950501_86975501_295C;SPAN=16079;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:109 GQ:23.3 PL:[23.3, 0.0, 241.1] SR:16 DR:0 LR:-23.29 LO:33.88);ALT=T[chr7:86970839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	86971002	+	chr7	86974619	+	.	0	11	3437676_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3437676_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_86950501_86975501_312C;SPAN=3617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:137 GQ:0.6 PL:[0.0, 0.6, 333.3] SR:11 DR:0 LR:0.8057 LO:20.23);ALT=T[chr7:86974619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	86971003	+	chr7	86974357	+	.	0	10	3437677_1	2.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=3437677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_86950501_86975501_194C;SPAN=3354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:115 GQ:2 PL:[2.0, 0.0, 275.9] SR:10 DR:0 LR:-1.854 LO:18.75);ALT=G[chr7:86974357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	87835819	+	chr7	87837822	+	.	3	40	3440459_1	54.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=3440459_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAGTAAGT;SCTG=c_7_87832501_87857501_13C;SPAN=2003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:112 GQ:54.1 PL:[54.1, 0.0, 86.0] SR:40 DR:3 LR:-53.66 LO:54.34);ALT=A[chr7:87837822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	87835819	+	chr7	87838654	+	ATCATCATATGGGAAATTCACAACACCTTGCTGAGCAGTATCCCGTCTTCGAAAGCTGT	5	66	3440460_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTGTAA;INSERTION=ATCATCATATGGGAAATTCACAACACCTTGCTGAGCAGTATCCCGTCTTCGAAAGCTGT;MAPQ=60;MATEID=3440460_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_87832501_87857501_13C;SPAN=2835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:119 GQ:89.9 PL:[198.8, 0.0, 89.9] SR:66 DR:5 LR:-201.1 LO:201.1);ALT=A[chr7:87838654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	87839500	+	chr7	87849290	+	.	17	0	3440477_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3440477_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:87839500(+)-7:87849290(-)__7_87832501_87857501D;SPAN=9790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:109 GQ:26.6 PL:[26.6, 0.0, 237.8] SR:0 DR:17 LR:-26.59 LO:36.49);ALT=A[chr7:87849290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	87840296	+	chr7	87849291	+	.	10	0	3440483_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3440483_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:87840296(+)-7:87849291(-)__7_87832501_87857501D;SPAN=8995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=C[chr7:87849291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	89810409	+	chr7	89812600	+	.	81	81	3446317_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=3446317_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_89792501_89817501_168C;SPAN=2191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:37 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:81 DR:81 LR:-399.4 LO:399.4);ALT=C[chr7:89812600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	89976116	+	chr7	89982126	+	.	8	0	3447064_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3447064_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:89976116(+)-7:89982126(-)__7_89964001_89989001D;SPAN=6010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=C[chr7:89982126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98923627	+	chr7	98930945	+	.	8	7	3477630_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=3477630_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98906501_98931501_22C;SPAN=7318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:98 GQ:13.1 PL:[13.1, 0.0, 224.3] SR:7 DR:8 LR:-13.06 LO:24.39);ALT=G[chr7:98930945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98923660	+	chr7	98935803	+	.	15	0	3477689_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3477689_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:98923660(+)-7:98935803(-)__7_98931001_98956001D;SPAN=12143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:59 GQ:33.5 PL:[33.5, 0.0, 109.4] SR:0 DR:15 LR:-33.53 LO:35.79);ALT=G[chr7:98935803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98972405	+	chr7	98983323	+	.	95	27	3478075_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3478075_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98980001_99005001_174C;SPAN=10918;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:72 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:27 DR:95 LR:-280.6 LO:280.6);ALT=G[chr7:98983323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98975079	+	chr7	98983321	+	.	0	18	3477895_1	45.0	.	EVDNC=ASSMB;HOMSEQ=ACAGG;MAPQ=60;MATEID=3477895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98955501_98980501_80C;SPAN=8242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:50 GQ:45.8 PL:[45.8, 0.0, 75.5] SR:18 DR:0 LR:-45.87 LO:46.27);ALT=G[chr7:98983321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98985890	+	chr7	98987527	+	.	4	11	3478106_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGGGT;MAPQ=60;MATEID=3478106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98980001_99005001_36C;SPAN=1637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:113 GQ:15.8 PL:[15.8, 0.0, 256.7] SR:11 DR:4 LR:-15.6 LO:28.53);ALT=T[chr7:98987527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98988877	+	chr7	98990293	+	.	14	7	3478121_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3478121_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98980001_99005001_63C;SPAN=1416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:98 GQ:36.2 PL:[36.2, 0.0, 201.2] SR:7 DR:14 LR:-36.17 LO:42.77);ALT=G[chr7:98990293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98990499	+	chr7	98991649	+	.	0	34	3478127_1	82.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=3478127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_98980001_99005001_129C;SPAN=1150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:111 GQ:82.4 PL:[82.4, 0.0, 184.7] SR:34 DR:0 LR:-82.16 LO:84.42);ALT=G[chr7:98991649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98990544	+	chr7	98992071	+	.	13	0	3478128_1	10.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3478128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:98990544(+)-7:98992071(-)__7_98980001_99005001D;SPAN=1527;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:119 GQ:10.7 PL:[10.7, 0.0, 278.0] SR:0 DR:13 LR:-10.67 LO:25.74);ALT=G[chr7:98992071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	98998093	+	chr7	99006157	+	.	8	0	3478311_1	11.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=3478311_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:98998093(+)-7:99006157(-)__7_99004501_99029501D;SPAN=8064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=A[chr7:99006157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99002622	+	chr7	99006157	+	.	10	0	3478313_1	17.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=3478313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99002622(+)-7:99006157(-)__7_99004501_99029501D;SPAN=3535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=T[chr7:99006157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99006156	-	chr12	119632708	+	.	41	0	5361551_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5361551_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99006156(-)-12:119632708(-)__12_119609001_119634001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:41 LR:-132.0 LO:132.0);ALT=[chr12:119632708[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	99006678	+	chr7	99008684	+	.	37	0	3478319_1	95.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3478319_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99006678(+)-7:99008684(-)__7_99004501_99029501D;SPAN=2006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:98 GQ:95.6 PL:[95.6, 0.0, 141.8] SR:0 DR:37 LR:-95.59 LO:96.09);ALT=A[chr7:99008684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99008809	+	chr7	99013759	+	.	0	14	3478335_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=3478335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_99004501_99029501_289C;SPAN=4950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:97 GQ:20 PL:[20.0, 0.0, 214.7] SR:14 DR:0 LR:-19.93 LO:29.53);ALT=G[chr7:99013759[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99015219	+	chr7	99017013	+	.	2	52	3478368_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3478368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_99004501_99029501_371C;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:132 GQ:99 PL:[139.4, 0.0, 179.0] SR:52 DR:2 LR:-139.2 LO:139.5);ALT=G[chr7:99017013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99040900	+	chr12	56194345	+	.	0	36	5201921_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CACATCAACAGTTTTTT;MAPQ=60;MATEID=5201921_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_56178501_56203501_90C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:47 GQ:7.1 PL:[106.1, 0.0, 7.1] SR:36 DR:0 LR:-111.1 LO:111.1);ALT=T[chr12:56194345[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	99041062	+	chr12	56211447	+	.	51	0	5202108_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5202108_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99041062(+)-12:56211447(-)__12_56203001_56228001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:68 GQ:14.6 PL:[149.9, 0.0, 14.6] SR:0 DR:51 LR:-156.4 LO:156.4);ALT=A[chr12:56211447[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	99056010	+	chr7	99063733	+	.	13	0	3478462_1	6.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=3478462_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99056010(+)-7:99063733(-)__7_99053501_99078501D;SPAN=7723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:136 GQ:6.2 PL:[6.2, 0.0, 323.0] SR:0 DR:13 LR:-6.067 LO:24.94);ALT=T[chr7:99063733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99056908	+	chr7	99063733	+	.	31	0	3478463_1	67.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=3478463_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99056908(+)-7:99063733(-)__7_99053501_99078501D;SPAN=6825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:128 GQ:67.7 PL:[67.7, 0.0, 242.6] SR:0 DR:31 LR:-67.65 LO:73.21);ALT=A[chr7:99063733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99057820	+	chr7	99063733	+	.	11	0	3478467_1	1.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=3478467_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99057820(+)-7:99063733(-)__7_99053501_99078501D;SPAN=5913;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:129 GQ:1.4 PL:[1.4, 0.0, 311.6] SR:0 DR:11 LR:-1.362 LO:20.53);ALT=A[chr7:99063733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99156563	+	chr7	99158154	+	.	20	0	3478700_1	36.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3478700_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99156563(+)-7:99158154(-)__7_99151501_99176501D;SPAN=1591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:109 GQ:36.5 PL:[36.5, 0.0, 227.9] SR:0 DR:20 LR:-36.49 LO:44.49);ALT=C[chr7:99158154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99274420	-	chr7	99275557	+	.	8	0	3479306_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3479306_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99274420(-)-7:99275557(-)__7_99249501_99274501D;SPAN=1137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=[chr7:99275557[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	99613350	+	chr7	99621041	+	.	17	2	3480634_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3480634_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_99617001_99642001_476C;SPAN=7691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:59 GQ:40.1 PL:[40.1, 0.0, 102.8] SR:2 DR:17 LR:-40.13 LO:41.66);ALT=G[chr7:99621041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99697418	+	chr7	99698897	+	.	33	0	3480936_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3480936_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99697418(+)-7:99698897(-)__7_99690501_99715501D;SPAN=1479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:87 GQ:85.4 PL:[85.4, 0.0, 125.0] SR:0 DR:33 LR:-85.36 LO:85.79);ALT=A[chr7:99698897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99697741	+	chr7	99698918	+	.	13	0	3480939_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3480939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99697741(+)-7:99698918(-)__7_99690501_99715501D;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=A[chr7:99698918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99746760	+	chr7	99751020	+	.	122	0	3481465_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3481465_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99746760(+)-7:99751020(-)__7_99739501_99764501D;SPAN=4260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:149 GQ:0.6 PL:[363.0, 0.6, 0.0] SR:0 DR:122 LR:-385.1 LO:385.1);ALT=G[chr7:99751020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99747202	+	chr7	99751022	+	.	29	54	3481467_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3481467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_99739501_99764501_296C;SPAN=3820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:177 GQ:99 PL:[206.3, 0.0, 222.8] SR:54 DR:29 LR:-206.2 LO:206.3);ALT=G[chr7:99751022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99747240	+	chr7	99751488	+	.	31	0	3481468_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3481468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99747240(+)-7:99751488(-)__7_99739501_99764501D;SPAN=4248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:164 GQ:58.1 PL:[58.1, 0.0, 338.6] SR:0 DR:31 LR:-57.9 LO:69.4);ALT=A[chr7:99751488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99928173	+	chr7	99930065	+	.	0	29	3482937_1	67.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=17;MATEID=3482937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_99911001_99936001_175C;SPAN=1892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:104 GQ:67.7 PL:[67.7, 0.0, 183.2] SR:29 DR:0 LR:-67.55 LO:70.58);ALT=C[chr7:99930065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	99930229	+	chr7	99933460	+	.	35	0	3482947_1	86.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=3482947_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:99930229(+)-7:99933460(-)__7_99911001_99936001D;SPAN=3231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:106 GQ:86.9 PL:[86.9, 0.0, 169.4] SR:0 DR:35 LR:-86.82 LO:88.31);ALT=A[chr7:99933460[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100271547	+	chr7	100273797	+	.	91	13	3484111_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3484111_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_100254001_100279001_52C;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:97 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:13 DR:91 LR:-287.2 LO:287.2);ALT=G[chr7:100273797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100271594	+	chr7	100274156	+	.	25	0	3484112_1	53.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=3484112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100271594(+)-7:100274156(-)__7_100254001_100279001D;SPAN=2562;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:108 GQ:53.3 PL:[53.3, 0.0, 208.4] SR:0 DR:25 LR:-53.27 LO:58.47);ALT=C[chr7:100274156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100327586	+	chr7	100340717	+	.	26	25	3484159_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GCTCACTGCAACCT;MAPQ=9;MATEID=3484159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_100327501_100352501_182C;SPAN=13131;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:69 GQ:37.4 PL:[129.8, 0.0, 37.4] SR:25 DR:26 LR:-132.7 LO:132.7);ALT=T[chr7:100340717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100479864	+	chr7	100481690	+	.	0	7	3484875_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=3484875_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_100474501_100499501_229C;SPAN=1826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:111 GQ:6.6 PL:[0.0, 6.6, 280.5] SR:7 DR:0 LR:6.966 LO:12.11);ALT=T[chr7:100481690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100533453	+	chr7	100536238	+	.	60	45	3485291_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAGGTTGCAGTGAG;MAPQ=60;MATEID=3485291_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_7_100523501_100548501_71C;SPAN=2785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:87 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:45 DR:60 LR:-256.6 LO:256.6);ALT=G[chr7:100536238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100676566	+	chr7	100677773	+	.	2	11	3485723_1	8.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACTGCTGAAGGTACCAGCATGCCAACCTCAACT;MAPQ=60;MATEID=3485723_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_100670501_100695501_335C;SPAN=1207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:126 GQ:8.9 PL:[8.9, 0.0, 296.0] SR:11 DR:2 LR:-8.777 LO:25.39);ALT=T[chr7:100677773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100797841	+	chr7	100799892	+	.	14	0	3486189_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3486189_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100797841(+)-7:100799892(-)__7_100793001_100818001D;SPAN=2051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:96 GQ:20.3 PL:[20.3, 0.0, 211.7] SR:0 DR:14 LR:-20.21 LO:29.6);ALT=T[chr7:100799892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100797847	+	chr7	100800655	+	.	8	0	3486190_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3486190_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100797847(+)-7:100800655(-)__7_100793001_100818001D;SPAN=2808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:96 GQ:0.5 PL:[0.5, 0.0, 231.5] SR:0 DR:8 LR:-0.3992 LO:14.85);ALT=G[chr7:100800655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100861545	+	chr7	100865880	+	.	51	0	3486487_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3486487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100861545(+)-7:100865880(-)__7_100842001_100867001D;SPAN=4335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:109 GQ:99 PL:[138.8, 0.0, 125.6] SR:0 DR:51 LR:-138.9 LO:138.9);ALT=C[chr7:100865880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100861549	+	chr7	100866756	+	.	33	0	3487180_1	91.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3487180_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100861549(+)-7:100866756(-)__7_100866501_100891501D;SPAN=5207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=G[chr7:100866756[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100883578	+	chr7	100888240	+	.	18	0	3487260_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3487260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:100883578(+)-7:100888240(-)__7_100866501_100891501D;SPAN=4662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:119 GQ:27.2 PL:[27.2, 0.0, 261.5] SR:0 DR:18 LR:-27.18 LO:38.37);ALT=G[chr7:100888240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	100884188	+	chr7	100888241	+	CTCGAGCAGCACGATGCCTTTACGGATGTCATCATTGTACTTGCTCCGCACCAGGCACCAGGCGTACTCAAACTGCGTGCTCTTGGACACCGAGCCTGCTGCCTTCTCAGACTGAAATTTCTTTTCAAACTT	37	101	3487264_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTCGAGCAGCACGATGCCTTTACGGATGTCATCATTGTACTTGCTCCGCACCAGGCACCAGGCGTACTCAAACTGCGTGCTCTTGGACACCGAGCCTGCTGCCTTCTCAGACTGAAATTTCTTTTCAAACTT;MAPQ=60;MATEID=3487264_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_100866501_100891501_246C;SPAN=4053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:138 GQ:2.3 PL:[332.3, 0.0, 2.3] SR:101 DR:37 LR:-352.4 LO:352.4);ALT=C[chr7:100888241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101001266	+	chr7	101003796	+	.	50	28	3489005_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCAATTTTTGTATTTTT;MAPQ=38;MATEID=3489005_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_7_100989001_101014001_394C;SPAN=2530;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:56 GQ:21 PL:[231.0, 21.0, 0.0] SR:28 DR:50 LR:-231.1 LO:231.1);ALT=T[chr7:101003796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101059188	+	chr7	101060267	+	.	45	36	3488111_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CCCGCCTCAGCCTCCCAAAGTGCTGGGATTA;MAPQ=60;MATEID=3488111_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_7_101038001_101063001_241C;SPAN=1079;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:72 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:36 DR:45 LR:-211.3 LO:211.3);ALT=A[chr7:101060267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101459373	+	chr7	101559392	+	.	36	9	3490506_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=3490506_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_101552501_101577501_190C;SPAN=100019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:9 DR:36 LR:-118.8 LO:118.8);ALT=G[chr7:101559392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	101724546	+	chr7	101727700	-	.	15	23	3491343_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=3491343_2;MATENM=3;NM=0;NUMPARTS=3;REPSEQ=TATA;SCTG=c_7_101724001_101749001_333C;SPAN=3154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:54 GQ:28.4 PL:[101.0, 0.0, 28.4] SR:23 DR:15 LR:-103.0 LO:103.0);ALT=T]chr7:101727700];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	101724546	+	chr7	101728039	+	ATATATTGTCTTCAAGGGCATATGGACAATTCAAGAAAACTTCAAAAAAATTTCTAGAGCTAATACGTGAGCATTAAGAGGTCACCTATATTATTATTATATAAACATTACATAATATAAAATATATATTTATATATATTTTATTATTTGTTAAAATGTAAAA	8	45	3491344_1	99.0	.	DISC_MAPQ=52;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=ATATATTGTCTTCAAGGGCATATGGACAATTCAAGAAAACTTCAAAAAAATTTCTAGAGCTAATACGTGAGCATTAAGAGGTCACCTATATTATTATTATATAAACATTACATAATATAAAATATATATTTATATATATTTTATTATTTGTTAAAATGTAAAA;MAPQ=60;MATEID=3491344_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_101724001_101749001_333C;SPAN=3493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:84 GQ:63.2 PL:[139.1, 0.0, 63.2] SR:45 DR:8 LR:-140.5 LO:140.5);ALT=T[chr7:101728039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102036985	+	chr7	102038066	+	.	0	5	3493347_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=3493347_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_102018001_102043001_85C;SPAN=1081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:111 GQ:13.2 PL:[0.0, 13.2, 293.7] SR:5 DR:0 LR:13.57 LO:7.905);ALT=G[chr7:102038066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102074149	+	chr7	102079389	+	.	20	0	3492409_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3492409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:102074149(+)-7:102079389(-)__7_102067001_102092001D;SPAN=5240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:92 GQ:41.3 PL:[41.3, 0.0, 179.9] SR:0 DR:20 LR:-41.1 LO:46.15);ALT=T[chr7:102079389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102076780	+	chr7	102079390	+	.	0	10	3492421_1	3.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3492421_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_102067001_102092001_240C;SPAN=2610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:109 GQ:3.5 PL:[3.5, 0.0, 260.9] SR:10 DR:0 LR:-3.479 LO:19.0);ALT=G[chr7:102079390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102937986	+	chr7	102939888	+	.	9	0	3496863_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3496863_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:102937986(+)-7:102939888(-)__7_102924501_102949501D;SPAN=1902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:112 GQ:0.3 PL:[0.0, 0.3, 270.6] SR:0 DR:9 LR:0.6346 LO:16.56);ALT=T[chr7:102939888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102938005	+	chr7	102939014	+	.	24	6	3496864_1	51.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3496864_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_102924501_102949501_79C;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:128 GQ:51.2 PL:[51.2, 0.0, 259.1] SR:6 DR:24 LR:-51.15 LO:59.12);ALT=G[chr7:102939014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102963242	+	chr7	102966990	+	ATTCTGCTTTTTCTTTTTCTTCTTCATCTAAATAAGAAAATTCTCTCCAAGAATCAAAATTATACCAGAAAGAATAAAATATATCTACATCTTCAAATGATGAATTCATATCACCAAGTTTAGGAACATTTTTTTTATTTGACCAT	0	13	3497102_1	14.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATTCTGCTTTTTCTTTTTCTTCTTCATCTAAATAAGAAAATTCTCTCCAAGAATCAAAATTATACCAGAAAGAATAAAATATATCTACATCTTCAAATGATGAATTCATATCACCAAGTTTAGGAACATTTTTTTTATTTGACCAT;MAPQ=60;MATEID=3497102_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_102949001_102974001_78C;SPAN=3748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:106 GQ:14.3 PL:[14.3, 0.0, 242.0] SR:13 DR:0 LR:-14.2 LO:26.43);ALT=C[chr7:102966990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102965012	+	chr7	102966990	+	.	2	8	3497112_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=3497112_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AA;SCTG=c_7_102949001_102974001_78C;SPAN=1978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:8 DR:2 LR:-4.292 LO:19.12);ALT=G[chr7:102966990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102982402	+	chr7	102985006	+	.	25	33	3497496_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3497496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_102973501_102998501_221C;SPAN=2604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:143 GQ:99 PL:[116.6, 0.0, 228.8] SR:33 DR:25 LR:-116.4 LO:118.5);ALT=C[chr7:102985006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	102989065	-	chr14	50053034	+	.	29	0	5735648_1	0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=5735648_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:102989065(-)-14:50053034(-)__14_50029001_50054001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:29 DP:1186 GQ:99 PL:[0.0, 225.2, 3330.0] SR:0 DR:29 LR:225.6 LO:38.11);ALT=[chr14:50053034[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	104612302	+	chr7	104485067	+	.	57	37	3503166_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3503166_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104590501_104615501_205C;SPAN=127235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:82 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:37 DR:57 LR:-244.3 LO:244.3);ALT=]chr7:104612302]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr7	104654983	+	chr7	104681282	+	.	0	34	3502681_1	96.0	.	EVDNC=ASSMB;HOMSEQ=ACAGG;MAPQ=60;MATEID=3502681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104639501_104664501_128C;SPAN=26299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:59 GQ:46.7 PL:[96.2, 0.0, 46.7] SR:34 DR:0 LR:-97.17 LO:97.17);ALT=G[chr7:104681282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104678647	+	chr7	104681285	+	.	3	13	3502959_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3502959_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_7_104664001_104689001_288C;SPAN=2638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:134 GQ:10.1 PL:[10.1, 0.0, 313.7] SR:13 DR:3 LR:-9.91 LO:27.43);ALT=G[chr7:104681285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104702726	+	chr7	104703797	+	.	2	3	3503452_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3503452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104688501_104713501_305C;SPAN=1071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:112 GQ:13.5 PL:[0.0, 13.5, 297.0] SR:3 DR:2 LR:13.84 LO:7.886);ALT=G[chr7:104703797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104715280	+	chr7	104717414	+	.	9	0	3503717_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3503717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:104715280(+)-7:104717414(-)__7_104713001_104738001D;SPAN=2134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:0 DR:9 LR:-3.158 LO:17.1);ALT=T[chr7:104717414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104717880	+	chr7	104722133	+	ACCATACCCTTTTGTGTTATTCTACTCTAAATTTCATGGGCTAGAAATGTGTGTTGATGCAAGGACTTTTGGGAATGAGGCTCGATTCATCAGGCGGTCTTGTACACCCAATGCAG	0	19	3503729_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=ACCATACCCTTTTGTGTTATTCTACTCTAAATTTCATGGGCTAGAAATGTGTGTTGATGCAAGGACTTTTGGGAATGAGGCTCGATTCATCAGGCGGTCTTGTACACCCAATGCAG;MAPQ=60;MATEID=3503729_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_104713001_104738001_337C;SPAN=4253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:90 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:19 DR:0 LR:-38.34 LO:43.57);ALT=G[chr7:104722133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104717880	+	chr7	104719291	+	.	0	4	3503728_1	0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3503728_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_7_104713001_104738001_337C;SPAN=1411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:88 GQ:10.5 PL:[0.0, 10.5, 234.3] SR:4 DR:0 LR:10.64 LO:6.34);ALT=G[chr7:104719291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104719412	+	chr7	104722133	+	.	3	15	3503732_1	25.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=3503732_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_104713001_104738001_337C;SPAN=2721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:114 GQ:25.4 PL:[25.4, 0.0, 249.8] SR:15 DR:3 LR:-25.23 LO:36.13);ALT=T[chr7:104722133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104722244	+	chr7	104730455	+	.	0	9	3503743_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3503743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104713001_104738001_309C;SPAN=8211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:115 GQ:1.2 PL:[0.0, 1.2, 280.5] SR:9 DR:0 LR:1.447 LO:16.45);ALT=G[chr7:104730455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104787108	+	chr7	104800952	+	.	0	10	3503601_1	1.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=3503601_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_104786501_104811501_60C;SPAN=13844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:118 GQ:1.1 PL:[1.1, 0.0, 284.9] SR:10 DR:0 LR:-1.041 LO:18.64);ALT=G[chr7:104800952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	104844269	+	chr7	105029259	+	.	13	0	3504625_1	36.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3504625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:104844269(+)-7:105029259(-)__7_105007001_105032001D;SPAN=184990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:23 GQ:17 PL:[36.8, 0.0, 17.0] SR:0 DR:13 LR:-36.98 LO:36.98);ALT=A[chr7:105029259[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105148992	+	chr7	105162497	+	.	0	7	3505650_1	9.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=3505650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105154001_105179001_114C;SPAN=13505;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:51 GQ:9.5 PL:[9.5, 0.0, 111.8] SR:7 DR:0 LR:-9.29 LO:14.6);ALT=C[chr7:105162497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105732386	+	chr7	105733395	+	.	6	14	3507949_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3507949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105717501_105742501_203C;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:120 GQ:30.2 PL:[30.2, 0.0, 261.2] SR:14 DR:6 LR:-30.21 LO:40.92);ALT=C[chr7:105733395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105733583	+	chr7	105738135	+	.	7	10	3507953_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3507953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105717501_105742501_313C;SPAN=4552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:105 GQ:14.6 PL:[14.6, 0.0, 239.0] SR:10 DR:7 LR:-14.47 LO:26.49);ALT=C[chr7:105738135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105738345	+	chr7	105739602	+	.	0	25	3507976_1	53.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=3507976_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105717501_105742501_107C;SPAN=1257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:106 GQ:53.9 PL:[53.9, 0.0, 202.4] SR:25 DR:0 LR:-53.81 LO:58.7);ALT=T[chr7:105739602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105738390	+	chr7	105752585	+	.	20	0	3507977_1	53.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=3507977_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:105738390(+)-7:105752585(-)__7_105717501_105742501D;SPAN=14195;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:46 GQ:53.6 PL:[53.6, 0.0, 56.9] SR:0 DR:20 LR:-53.56 LO:53.57);ALT=G[chr7:105752585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	105739729	+	chr7	105752586	+	.	76	44	3507980_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3507980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_105717501_105742501_365C;SPAN=12857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:68 GQ:24 PL:[264.0, 24.0, 0.0] SR:44 DR:76 LR:-264.1 LO:264.1);ALT=C[chr7:105752586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	104432708	+	chr7	105766146	+	.	10	0	4004219_1	22.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=4004219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:105766146(-)-8:104432708(+)__8_104419001_104444001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:41 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-21.9 LO:23.65);ALT=]chr8:104432708]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	109232059	+	chr7	109235968	+	.	18	30	3519366_1	99.0	.	DISC_MAPQ=2;EVDNC=ASDIS;HOMSEQ=A;MAPQ=33;MATEID=3519366_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_109221001_109246001_209C;SPAN=3909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:88 GQ:81.8 PL:[131.3, 0.0, 81.8] SR:30 DR:18 LR:-131.9 LO:131.9);ALT=A[chr7:109235968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54832698	+	chr7	109235968	+	.	5	18	6867054_1	43.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=6867054_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54831001_54856001_58C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:60 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:18 DR:5 LR:-43.16 LO:44.49);ALT=]chr19:54832698]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	125264220	+	chr12	74014367	+	ATTATA	49	58	3568962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTATA;MAPQ=60;MATEID=3568962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_125244001_125269001_225C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:61 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:58 DR:49 LR:-254.2 LO:254.2);ALT=C[chr12:74014367[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	125746123	+	chr7	126166901	+	T	47	38	3570834_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=3570834_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_126150501_126175501_101C;SPAN=420778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:63 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:38 DR:47 LR:-211.3 LO:211.3);ALT=A[chr7:126166901[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	126045889	+	chr7	126051448	+	.	50	53	3570696_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAC;MAPQ=60;MATEID=3570696_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_7_126028001_126053001_151C;SPAN=5559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:25 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:53 DR:50 LR:-257.5 LO:257.5);ALT=C[chr7:126051448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	126098488	-	chr7	126167441	+	.	39	48	3570835_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAT;MAPQ=60;MATEID=3570835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_126150501_126175501_371C;SPAN=68953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:72 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:48 DR:39 LR:-234.4 LO:234.4);ALT=[chr7:126167441[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	127292505	+	chr7	127316821	+	.	2	5	3576151_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3576151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_127277501_127302501_488C;SPAN=24316;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:106 GQ:12 PL:[0.0, 12.0, 280.5] SR:5 DR:2 LR:12.21 LO:8.007);ALT=G[chr7:127316821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	127292507	+	chr7	127326666	+	.	9	15	3576726_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=3576726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_127302001_127327001_571C;SPAN=34159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:86 GQ:32.9 PL:[32.9, 0.0, 174.8] SR:15 DR:9 LR:-32.82 LO:38.43);ALT=T[chr7:127326666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	127979847	+	chr7	127983729	+	.	0	14	3579721_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=3579721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_127963501_127988501_341C;SPAN=3882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:14 DP:189 GQ:4.9 PL:[0.0, 4.9, 468.7] SR:14 DR:0 LR:4.991 LO:25.24);ALT=T[chr7:127983729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128096078	+	chr7	128097253	+	.	35	12	3580607_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3580607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_128086001_128111001_215C;SPAN=1175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:173 GQ:75.5 PL:[75.5, 0.0, 342.8] SR:12 DR:35 LR:-75.27 LO:85.08);ALT=G[chr7:128097253[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128379508	+	chr7	128388634	+	.	10	0	3582404_1	5.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3582404_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128379508(+)-7:128388634(-)__7_128355501_128380501D;SPAN=9126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:101 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.647 LO:19.35);ALT=C[chr7:128388634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128503047	+	chr12	48478956	+	.	40	0	3583351_1	97.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3583351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128503047(+)-12:48478956(-)__7_128502501_128527501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:128 GQ:97.4 PL:[97.4, 0.0, 212.9] SR:0 DR:40 LR:-97.36 LO:99.74);ALT=A[chr12:48478956[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	128503128	+	chr7	128505428	+	.	56	0	3583352_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3583352_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128503128(+)-7:128505428(-)__7_128502501_128527501D;SPAN=2300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:173 GQ:99 PL:[138.2, 0.0, 280.1] SR:0 DR:56 LR:-138.0 LO:140.7);ALT=C[chr7:128505428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128578155	+	chr7	128582120	+	.	38	0	3584032_1	86.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3584032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:128578155(+)-7:128582120(-)__7_128576001_128601001D;SPAN=3965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:146 GQ:86 PL:[86.0, 0.0, 267.5] SR:0 DR:38 LR:-85.88 LO:91.13);ALT=C[chr7:128582120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128582331	+	chr7	128585897	+	.	5	8	3584045_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3584045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_128576001_128601001_338C;SPAN=3566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:13 DP:168 GQ:2.5 PL:[0.0, 2.5, 412.6] SR:8 DR:5 LR:2.602 LO:23.69);ALT=G[chr7:128585897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	128658212	+	chr7	128694703	+	.	0	7	3584652_1	0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=3584652_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_128649501_128674501_266C;SPAN=36491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.547 LO:12.74);ALT=C[chr7:128694703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	129050411	+	chr9	116037593	+	.	33	0	3586964_1	91.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=3586964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:129050411(+)-9:116037593(-)__7_129041501_129066501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:66 GQ:68 PL:[91.1, 0.0, 68.0] SR:0 DR:33 LR:-91.21 LO:91.21);ALT=T[chr9:116037593[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	130061874	+	chr7	130080778	+	.	10	0	3593682_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3593682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:130061874(+)-7:130080778(-)__7_130070501_130095501D;SPAN=18904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=G[chr7:130080778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	130132181	+	chr7	130135206	+	.	6	29	3593934_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3593934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_130119501_130144501_130C;SPAN=3025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:159 GQ:59.3 PL:[59.3, 0.0, 326.6] SR:29 DR:6 LR:-59.25 LO:69.87);ALT=G[chr7:130135206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	130629208	+	chr7	130630479	+	.	0	4	3596213_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=3596213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_130609501_130634501_24C;SPAN=1271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:179 GQ:35.2 PL:[0.0, 35.2, 505.0] SR:4 DR:0 LR:35.29 LO:5.101);ALT=T[chr7:130630479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	130630595	+	chr7	130645881	+	.	20	7	3596222_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=3596222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_130609501_130634501_167C;SPAN=15286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:94 GQ:50.6 PL:[50.6, 0.0, 176.0] SR:7 DR:20 LR:-50.46 LO:54.43);ALT=C[chr7:130645881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45984207	+	chr7	131164309	+	.	9	40	3599195_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GGCGTGGTGGCTCATGCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=25;MATEID=3599195_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_7_131148501_131173501_193C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:81 GQ:67.4 PL:[126.8, 0.0, 67.4] SR:40 DR:9 LR:-127.5 LO:127.5);ALT=]chr11:45984207]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr7	131459651	-	chr7	131461419	+	.	9	0	3601077_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3601077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:131459651(-)-7:131461419(-)__7_131442501_131467501D;SPAN=1768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:135 GQ:6.6 PL:[0.0, 6.6, 339.9] SR:0 DR:9 LR:6.866 LO:15.8);ALT=[chr7:131461419[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	132720594	+	chr11	62341303	+	.	12	0	3607492_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=3607492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:132720594(+)-11:62341303(-)__7_132716501_132741501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:209 GQ:16.9 PL:[0.0, 16.9, 541.3] SR:0 DR:12 LR:17.01 LO:20.26);ALT=G[chr11:62341303[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	132937932	+	chr7	132959732	+	.	10	0	3608616_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3608616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:132937932(+)-7:132959732(-)__7_132937001_132962001D;SPAN=21800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:183 GQ:16.3 PL:[0.0, 16.3, 475.3] SR:0 DR:10 LR:16.57 LO:16.67);ALT=C[chr7:132959732[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	133785003	+	chr7	133798330	+	.	129	68	3612727_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TGC;MAPQ=60;MATEID=3612727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_133794501_133819501_217C;SPAN=13327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:161 DP:77 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:68 DR:129 LR:-475.3 LO:475.3);ALT=C[chr7:133798330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	134136507	+	chr7	134143749	+	.	17	9	3614795_1	41.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3614795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_134113001_134138001_259C;SPAN=7242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:81 GQ:41 PL:[41.0, 0.0, 153.2] SR:9 DR:17 LR:-40.77 LO:44.56);ALT=T[chr7:134143749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	134506355	+	chr7	134520910	-	.	8	21	3616672_1	52.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTGAGA;MAPQ=60;MATEID=3616672_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_7_134505001_134530001_147C;SPAN=14555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:135 GQ:52.7 PL:[52.7, 0.0, 273.8] SR:21 DR:8 LR:-52.55 LO:61.19);ALT=A]chr7:134520910];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	135347372	+	chr7	135358838	+	.	62	0	3621458_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3621458_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:135347372(+)-7:135358838(-)__7_135338001_135363001D;SPAN=11466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:189 GQ:99 PL:[153.5, 0.0, 305.3] SR:0 DR:62 LR:-153.5 LO:156.2);ALT=G[chr7:135358838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135614762	+	chr7	135636264	+	TTGACAGAAGCAATTTCACACAGGAAACATGACCCTCATAGACAGCAGACAGAAGAGGAGTAATATGATGTTTATCTGGAG	2	44	3622787_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTGACAGAAGCAATTTCACACAGGAAACATGACCCTCATAGACAGCAGACAGAAGAGGAGTAATATGATGTTTATCTGGAG;MAPQ=60;MATEID=3622787_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_135632001_135657001_223C;SPAN=21502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:64 GQ:22.4 PL:[131.3, 0.0, 22.4] SR:44 DR:2 LR:-135.4 LO:135.4);ALT=T[chr7:135636264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135614762	+	chr7	135635346	+	.	2	35	3623216_1	97.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=3623216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_135607501_135632501_368C;SPAN=20584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:92 GQ:97.4 PL:[97.4, 0.0, 123.8] SR:35 DR:2 LR:-97.21 LO:97.42);ALT=T[chr7:135635346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	135636380	+	chr7	135661776	+	.	0	41	3623309_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=3623309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_135656501_135681501_21C;SPAN=25396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:118 GQ:99 PL:[103.4, 0.0, 182.6] SR:41 DR:0 LR:-103.4 LO:104.6);ALT=T[chr7:135661776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	136792551	-	chr7	136793794	+	.	8	0	3628661_1	0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=3628661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:136792551(-)-7:136793794(-)__7_136783501_136808501D;SPAN=1243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:145 GQ:12.6 PL:[0.0, 12.6, 376.2] SR:0 DR:8 LR:12.88 LO:13.37);ALT=[chr7:136793794[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	137613141	+	chr7	137620615	+	.	32	0	3632445_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3632445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:137613141(+)-7:137620615(-)__7_137616501_137641501D;SPAN=7474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:61 GQ:56.3 PL:[89.3, 0.0, 56.3] SR:0 DR:32 LR:-89.43 LO:89.43);ALT=G[chr7:137620615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	138474601	-	chr10	101990953	+	.	10	0	3638842_1	14.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3638842_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:138474601(-)-10:101990953(-)__7_138474001_138499001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-14.05 LO:21.05);ALT=[chr10:101990953[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	139026270	+	chr7	139030246	+	.	46	32	3641275_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=3641275_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139013001_139038001_355C;SPAN=3976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:177 GQ:99 PL:[160.1, 0.0, 269.0] SR:32 DR:46 LR:-160.0 LO:161.5);ALT=T[chr7:139030246[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139090534	+	chr7	139091918	+	.	7	9	3642248_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3642248_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139086501_139111501_281C;SPAN=1384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:153 GQ:8.3 PL:[8.3, 0.0, 361.4] SR:9 DR:7 LR:-8.064 LO:28.95);ALT=G[chr7:139091918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139218974	-	chr14	69864948	+	.	85	8	3642952_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CATCGCGCCAAACTCT;MAPQ=32;MATEID=3642952_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_7_139209001_139234001_457C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:83 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:8 DR:85 LR:-267.4 LO:267.4);ALT=[chr14:69864948[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr7	139529281	+	chr7	139572033	+	.	0	34	3645082_1	88.0	.	EVDNC=ASSMB;HOMSEQ=GGTA;MAPQ=60;MATEID=3645082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139552001_139577001_30C;SPAN=42752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:88 GQ:88.4 PL:[88.4, 0.0, 124.7] SR:34 DR:0 LR:-88.39 LO:88.74);ALT=A[chr7:139572033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139572128	+	chr7	139611023	+	GTTTTTGGGAAAGCCAAATGGAGCTCAGAAAGCTGTATGGACCTCTGTGTG	3	17	3645184_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GGTA;INSERTION=GTTTTTGGGAAAGCCAAATGGAGCTCAGAAAGCTGTATGGACCTCTGTGTG;MAPQ=60;MATEID=3645184_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_139552001_139577001_543C;SPAN=38895;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:85 GQ:43.1 PL:[43.1, 0.0, 161.9] SR:17 DR:3 LR:-42.99 LO:46.94);ALT=G[chr7:139611023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139655439	+	chr7	139657432	+	.	9	0	3645248_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3645248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:139655439(+)-7:139657432(-)__7_139650001_139675001D;SPAN=1993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:154 GQ:11.8 PL:[0.0, 11.8, 396.0] SR:0 DR:9 LR:12.01 LO:15.27);ALT=G[chr7:139657432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139657563	+	chr7	139661716	+	.	9	2	3645258_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3645258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139650001_139675001_296C;SPAN=4153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:150 GQ:4.3 PL:[0.0, 4.3, 372.9] SR:2 DR:9 LR:4.328 LO:19.78);ALT=G[chr7:139661716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139715662	+	chr7	139717469	+	.	2	2	3645457_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3645457_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139699001_139724001_131C;SPAN=1807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:181 GQ:35.5 PL:[0.0, 35.5, 508.3] SR:2 DR:2 LR:35.83 LO:5.082);ALT=T[chr7:139717469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	139717635	+	chr7	139719823	+	.	0	25	3645472_1	40.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=3645472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_139699001_139724001_149C;SPAN=2188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:157 GQ:40.1 PL:[40.1, 0.0, 340.4] SR:25 DR:0 LR:-39.99 LO:53.91);ALT=T[chr7:139719823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140171814	+	chr7	140178957	+	.	13	12	3648456_1	25.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=TACCTG;MAPQ=60;MATEID=3648456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_140164501_140189501_336C;SPAN=7143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:137 GQ:25.7 PL:[25.7, 0.0, 306.2] SR:12 DR:13 LR:-25.6 LO:39.73);ALT=G[chr7:140178957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140396642	+	chr7	140402666	+	.	0	65	3650447_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3650447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_140385001_140410001_282C;SPAN=6024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:226 GQ:99 PL:[153.4, 0.0, 394.4] SR:65 DR:0 LR:-153.3 LO:159.2);ALT=A[chr7:140402666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140397040	+	chr7	140404658	+	.	18	0	3650449_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3650449_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:140397040(+)-7:140404658(-)__7_140385001_140410001D;SPAN=7618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:18 DP:220 GQ:0.1 PL:[0.0, 0.1, 534.7] SR:0 DR:18 LR:0.1854 LO:33.26);ALT=G[chr7:140404658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140397086	+	chr7	140402665	+	.	69	0	3650450_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3650450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:140397086(+)-7:140402665(-)__7_140385001_140410001D;SPAN=5579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:209 GQ:99 PL:[171.2, 0.0, 336.2] SR:0 DR:69 LR:-171.1 LO:174.1);ALT=T[chr7:140402665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140402811	+	chr7	140406363	+	GTCACTTTCCGTATCCTGATCCTTCCCAGTGGACAGATGAAGAATTAGGTATCCCTCCTGATGATGAAGACTGAAGGTGTAGACTCAGCCTCACTCTGTACAA	4	105	3650473_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GTCACTTTCCGTATCCTGATCCTTCCCAGTGGACAGATGAAGAATTAGGTATCCCTCCTGATGATGAAGACTGAAGGTGTAGACTCAGCCTCACTCTGTACAA;MAPQ=60;MATEID=3650473_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_140385001_140410001_60C;SPAN=3552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:108 DP:220 GQ:99 PL:[296.9, 0.0, 237.5] SR:105 DR:4 LR:-297.3 LO:297.3);ALT=G[chr7:140406363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140402811	+	chr7	140404659	+	.	0	66	3650472_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3650472_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_7_140385001_140410001_60C;SPAN=1848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:264 GQ:99 PL:[146.5, 0.0, 493.1] SR:66 DR:0 LR:-146.3 LO:156.9);ALT=G[chr7:140404659[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140404764	+	chr7	140406363	+	.	2	27	3650484_1	53.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3650484_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_140385001_140410001_60C;SPAN=1599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:157 GQ:53.3 PL:[53.3, 0.0, 327.2] SR:27 DR:2 LR:-53.19 LO:64.6);ALT=G[chr7:140406363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140706338	+	chr7	140710219	+	.	0	20	3651960_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=3651960_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_140703501_140728501_318C;SPAN=3881;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:157 GQ:23.6 PL:[23.6, 0.0, 356.9] SR:20 DR:0 LR:-23.49 LO:41.02);ALT=G[chr7:140710219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140710461	+	chr7	140714350	+	.	10	3	3651987_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=57;MATEID=3651987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_140703501_140728501_507C;SPAN=3889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:155 GQ:1 PL:[1.0, 0.0, 374.0] SR:3 DR:10 LR:-0.9197 LO:24.17);ALT=C[chr7:140714350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	140710474	+	chr7	140714709	+	.	33	0	3651988_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3651988_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:140710474(+)-7:140714709(-)__7_140703501_140728501D;SPAN=4235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:188 GQ:58 PL:[58.0, 0.0, 398.0] SR:0 DR:33 LR:-58.0 LO:72.7);ALT=G[chr7:140714709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	141438434	+	chr7	141441965	+	.	24	0	3655417_1	58.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3655417_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:141438434(+)-7:141441965(-)__7_141414001_141439001D;SPAN=3531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:78 GQ:58.1 PL:[58.1, 0.0, 130.7] SR:0 DR:24 LR:-58.09 LO:59.65);ALT=C[chr7:141441965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	141438993	+	chr7	141443361	+	CTTCGTCAGTTTGTAAGACATGAGTCCGAAACAACTACCAGTTTGGTTCTTGAAAGAT	7	84	3655575_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=AGGTA;INSERTION=CTTCGTCAGTTTGTAAGACATGAGTCCGAAACAACTACCAGTTTGGTTCTTGAAAGAT;MAPQ=60;MATEID=3655575_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_141438501_141463501_402C;SPAN=4368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:192 GQ:99 PL:[245.3, 0.0, 218.9] SR:84 DR:7 LR:-245.1 LO:245.1);ALT=A[chr7:141443361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	141438993	+	chr7	141441967	+	.	2	28	3655574_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGTA;MAPQ=60;MATEID=3655574_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_7_141438501_141463501_402C;SPAN=2974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:174 GQ:52 PL:[52.0, 0.0, 368.9] SR:28 DR:2 LR:-51.89 LO:65.83);ALT=A[chr7:141441967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	141443505	+	chr7	141445295	+	TGTCAGTCAAAAGACAACATGGCACAGAATATCAGTATTCCGGCCAGGCCTCAGAGACGTGGCATATCAATATGTGAAAAAGG	3	102	3655594_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=TGTCAGTCAAAAGACAACATGGCACAGAATATCAGTATTCCGGCCAGGCCTCAGAGACGTGGCATATCAATATGTGAAAAAGG;MAPQ=60;MATEID=3655594_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_7_141438501_141463501_420C;SPAN=1790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:103 DP:183 GQ:99 PL:[290.6, 0.0, 152.0] SR:102 DR:3 LR:-292.7 LO:292.7);ALT=A[chr7:141445295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	141445384	+	chr7	141450110	+	.	0	54	3655605_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3655605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_141438501_141463501_406C;SPAN=4726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:151 GQ:99 PL:[137.6, 0.0, 226.7] SR:54 DR:0 LR:-137.3 LO:138.6);ALT=G[chr7:141450110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142359260	-	chr7	142362014	+	.	15	74	3659623_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CTT;MAPQ=60;MATEID=3659623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_142345001_142370001_98C;SPAN=2754;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:139 GQ:99 PL:[223.1, 0.0, 114.2] SR:74 DR:15 LR:-225.0 LO:225.0);ALT=[chr7:142362014[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	142553147	+	chr7	142558808	+	.	0	7	3660542_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=3660542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_142541001_142566001_328C;SPAN=5661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:147 GQ:16.6 PL:[0.0, 16.6, 389.4] SR:7 DR:0 LR:16.72 LO:11.24);ALT=G[chr7:142558808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142824847	+	chr7	142893908	+	.	109	47	3661916_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TTAAA;MAPQ=60;MATEID=3661916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_142884001_142909001_275C;SPAN=69061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:54 GQ:36 PL:[396.0, 36.0, 0.0] SR:47 DR:109 LR:-396.1 LO:396.1);ALT=A[chr7:142893908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142962185	+	chr7	142965184	+	AATGAAGACATCACCGAGCCGCAGAGCATCCTGGCGGCTGCAGAGAAGGCTGGTATGTCTGCAGAACAAGCCCAGGGACTTCTGGAAAAGATCGCAACGCCAAAGGTGAAGAACCAGCTCAAGGAGACCACTGAGGCAGCCTGCAGATACGGA	0	37	3662452_1	77.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATGAAGACATCACCGAGCCGCAGAGCATCCTGGCGGCTGCAGAGAAGGCTGGTATGTCTGCAGAACAAGCCCAGGGACTTCTGGAAAAGATCGCAACGCCAAAGGTGAAGAACCAGCTCAAGGAGACCACTGAGGCAGCCTGCAGATACGGA;MAPQ=60;MATEID=3662452_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_7_142957501_142982501_239C;SPAN=2999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:164 GQ:77.9 PL:[77.9, 0.0, 318.8] SR:37 DR:0 LR:-77.71 LO:86.06);ALT=G[chr7:142965184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	142962390	+	chr7	142964709	+	.	9	20	3662453_1	41.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3662453_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_7_142957501_142982501_239C;SPAN=2319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:164 GQ:41.6 PL:[41.6, 0.0, 355.1] SR:20 DR:9 LR:-41.39 LO:56.01);ALT=G[chr7:142964709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	143086085	+	chr7	143087668	+	.	13	0	3663056_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3663056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:143086085(+)-7:143087668(-)__7_143080001_143105001D;SPAN=1583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:13 DP:228 GQ:18.7 PL:[0.0, 18.7, 590.8] SR:0 DR:13 LR:18.86 LO:21.91);ALT=G[chr7:143087668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	149731143	+	chr7	149735125	+	.	21	0	3688733_1	52.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=3688733_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:149731143(+)-7:149735125(-)__7_149719501_149744501D;SPAN=3982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:63 GQ:52.4 PL:[52.4, 0.0, 98.6] SR:0 DR:21 LR:-52.25 LO:53.09);ALT=C[chr7:149735125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	149734015	+	chr7	153757489	-	.	8	0	3688749_1	21.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=3688749_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:149734015(+)-7:153757489(+)__7_149719501_149744501D;SPAN=4023474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:18 GQ:21.5 PL:[21.5, 0.0, 21.5] SR:0 DR:8 LR:-21.53 LO:21.53);ALT=T]chr7:153757489];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	149847642	+	chr7	149849129	+	.	23	43	3689303_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;MAPQ=0;MATEID=3689303_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=CC;SCTG=c_7_149842001_149867001_377C;SECONDARY;SPAN=1487;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:87 GQ:39.2 PL:[171.2, 0.0, 39.2] SR:43 DR:23 LR:-175.8 LO:175.8);ALT=A[chr7:149849129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150066015	+	chr7	150068314	+	.	9	0	3689770_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3689770_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:150066015(+)-7:150068314(-)__7_150062501_150087501D;SPAN=2299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=A[chr7:150068314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150130917	+	chr7	150132117	+	.	0	16	3690306_1	23.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3690306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_150111501_150136501_194C;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:111 GQ:23 PL:[23.0, 0.0, 244.1] SR:16 DR:0 LR:-22.74 LO:33.74);ALT=G[chr7:150132117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150382887	+	chr7	150389401	+	.	15	0	3690995_1	20.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3690995_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:150382887(+)-7:150389401(-)__7_150381001_150406001D;SPAN=6514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:109 GQ:20 PL:[20.0, 0.0, 244.4] SR:0 DR:15 LR:-19.98 LO:31.31);ALT=T[chr7:150389401[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150413784	+	chr7	150417134	+	.	9	0	3691092_1	2.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3691092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:150413784(+)-7:150417134(-)__7_150405501_150430501D;SPAN=3350;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:0 DR:9 LR:-2.075 LO:16.94);ALT=C[chr7:150417134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150725700	+	chr7	150730689	+	.	8	4	3692102_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGTA;MAPQ=60;MATEID=3692102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_150724001_150749001_68C;SPAN=4989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:109 GQ:0.2 PL:[0.2, 0.0, 264.2] SR:4 DR:8 LR:-0.1782 LO:16.67);ALT=A[chr7:150730689[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	150746657	+	chr15	84810725	+	.	44	33	3692179_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=3692179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_150724001_150749001_17C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:31 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:33 DR:44 LR:-191.4 LO:191.4);ALT=C[chr15:84810725[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr7	150922077	+	chr7	150923391	+	.	0	9	3692549_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=3692549_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_150920001_150945001_4C;SPAN=1314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:9 DR:0 LR:-15.89 LO:19.85);ALT=G[chr7:150923391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	151038981	+	chr7	151046156	+	.	20	0	3692742_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3692742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:151038981(+)-7:151046156(-)__7_151042501_151067501D;SPAN=7175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:32 GQ:17.9 PL:[57.5, 0.0, 17.9] SR:0 DR:20 LR:-58.32 LO:58.32);ALT=G[chr7:151046156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	151042553	+	chr7	151046157	+	.	5	10	3692658_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=3692658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_151018001_151043001_72C;SPAN=3604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:23 GQ:17 PL:[36.8, 0.0, 17.0] SR:10 DR:5 LR:-36.98 LO:36.98);ALT=G[chr7:151046157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	151483628	+	chr7	151573591	+	.	0	7	3693665_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=3693665_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_151557001_151582001_272C;SPAN=89963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:21 GQ:17.6 PL:[17.6, 0.0, 30.8] SR:7 DR:0 LR:-17.42 LO:17.7);ALT=C[chr7:151573591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	152131009	+	chr22	17084686	-	.	16	0	7205705_1	33.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=7205705_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:152131009(+)-22:17084686(+)__22_17076501_17101501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:70 GQ:33.8 PL:[33.8, 0.0, 136.1] SR:0 DR:16 LR:-33.85 LO:37.32);ALT=T]chr22:17084686];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	152281703	+	chr7	152284306	+	.	43	38	3695637_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=CACATGTTTTA;MAPQ=60;MATEID=3695637_2;MATENM=2;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_7_152267501_152292501_263C;SPAN=2603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:37 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:38 DR:43 LR:-194.7 LO:194.7);ALT=A[chr7:152284306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	152574767	+	chr7	152760110	-	.	22	18	3696721_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAA;MAPQ=60;MATEID=3696721_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_7_152757501_152782501_91C;SPAN=185343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:24 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:18 DR:22 LR:-105.6 LO:105.6);ALT=T]chr7:152760110];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr7	152574806	+	chr7	152580428	+	.	15	0	3696274_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3696274_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:152574806(+)-7:152580428(-)__7_152561501_152586501D;SPAN=5622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:10 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=A[chr7:152580428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr7	152580431	-	chr7	152759969	+	.	24	0	3696722_1	71.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=3696722_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:152580431(-)-7:152759969(-)__7_152757501_152782501D;SPAN=179538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:30 GQ:1.7 PL:[71.0, 0.0, 1.7] SR:0 DR:24 LR:-75.13 LO:75.13);ALT=[chr7:152759969[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr7	152975471	+	chr9	94389041	-	.	10	0	3697078_1	7.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=3697078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:152975471(+)-9:94389041(+)__7_152953501_152978501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:0 DR:10 LR:-7.543 LO:19.68);ALT=A]chr9:94389041];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr7	154391983	+	chr7	154399731	+	.	24	0	3699278_1	69.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CCAGGCTGGAGTACAGTGGCACAATCTCAGCTCACTGCAAGCTCTGCCTCCCGGGTTCAAGCAATTCTCCTGCCTCAGCCTCCCAAGTAGCTGGGATTACAGGCA;MAPQ=60;MATEID=3699278_2;MATENM=5;NM=6;NUMPARTS=2;SCTG=c_7_154374501_154399501_110C;SPAN=7748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:0 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=A[chr7:154399731[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11098997	-	chr18	22222390	+	.	19	30	6563296_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=ACTACTGATAA;MAPQ=60;MATEID=6563296_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_22221501_22246501_210C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:41 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:30 DR:19 LR:-141.9 LO:141.9);ALT=[chr18:22222390[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	11245561	+	chr8	11247208	+	.	48	45	3743746_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAG;MAPQ=60;MATEID=3743746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11245501_11270501_317C;SPAN=1647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:66 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:45 DR:48 LR:-208.0 LO:208.0);ALT=G[chr8:11247208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11660440	+	chr8	11667173	+	.	18	4	3744849_1	49.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=3744849_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_8_11637501_11662501_99C;SPAN=6733;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:61 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:4 DR:18 LR:-49.49 LO:50.39);ALT=G[chr8:11667173[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11660441	+	chr8	11666300	+	.	50	23	3745060_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=3745060_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_11662001_11687001_301C;SPAN=5859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:60 GQ:9.6 PL:[165.0, 9.6, 0.0] SR:23 DR:50 LR:-167.9 LO:167.9);ALT=G[chr8:11666300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11683726	+	chr8	11687751	+	.	4	2	3745159_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3745159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11686501_11711501_383C;SPAN=4025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:2 DR:4 LR:-3.23 LO:9.742);ALT=T[chr8:11687751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11687931	+	chr8	11689025	+	.	7	7	3745165_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=3745165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11686501_11711501_217C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:101 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:7 DR:7 LR:-15.55 LO:26.73);ALT=T[chr8:11689025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11689179	+	chr8	11695895	+	.	7	5	3745169_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3745169_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_11686501_11711501_253C;SPAN=6716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:5 DR:7 LR:-7.051 LO:21.42);ALT=G[chr8:11695895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11710989	+	chr8	11725507	+	.	40	6	3745233_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=3745233_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_11686501_11711501_378C;SPAN=14518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:51 GQ:2.9 PL:[118.4, 0.0, 2.9] SR:6 DR:40 LR:-124.4 LO:124.4);ALT=C[chr8:11725507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	11893340	+	chr8	11788246	+	.	24	0	3745495_1	71.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=3745495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:11788246(-)-8:11893340(+)__8_11784501_11809501D;SPAN=105094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:30 GQ:1.7 PL:[71.0, 0.0, 1.7] SR:0 DR:24 LR:-75.13 LO:75.13);ALT=]chr8:11893340]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	12427810	+	chr8	12432836	+	GGAATTTTGTG	36	29	3752489_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;INSERTION=GGAATTTTGTG;MAPQ=60;MATEID=3752489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_12421501_12446501_1306C;SPAN=5026;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:256 GQ:99 PL:[118.9, 0.0, 501.8] SR:29 DR:36 LR:-118.8 LO:132.2);ALT=G[chr8:12432836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	14583503	-	chr8	14585046	+	.	2	3	3755509_1	0	.	DISC_MAPQ=50;EVDNC=ASDIS;MAPQ=60;MATEID=3755509_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_14577501_14602501_96C;SPAN=1543;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:3 DR:2 LR:13.62 LO:6.133);ALT=[chr8:14585046[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	15289364	+	chr13	74314062	-	.	57	70	3757473_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TATGTT;MAPQ=60;MATEID=3757473_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_15288001_15313001_184C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:31 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:70 DR:57 LR:-326.8 LO:326.8);ALT=T]chr13:74314062];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	15289367	-	chr13	74313858	+	.	72	80	3757475_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGGC;MAPQ=60;MATEID=3757475_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_15288001_15313001_68C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:31 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:80 DR:72 LR:-369.7 LO:369.7);ALT=[chr13:74313858[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr19	38178938	+	chr8	28739769	+	.	14	0	6807946_1	36.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6807946_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:28739769(-)-19:38178938(+)__19_38171001_38196001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:37 GQ:36.2 PL:[36.2, 0.0, 52.7] SR:0 DR:14 LR:-36.19 LO:36.38);ALT=]chr19:38178938]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	29921411	+	chr8	29923502	+	.	8	0	3801322_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3801322_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:29921411(+)-8:29923502(-)__8_29914501_29939501D;SPAN=2091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:0 DR:8 LR:-0.6702 LO:14.89);ALT=C[chr8:29923502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29924436	+	chr8	29927157	+	.	9	4	3801336_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=3801336_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_8_29914501_29939501_347C;SPAN=2721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:94 GQ:14.3 PL:[14.3, 0.0, 212.3] SR:4 DR:9 LR:-14.15 LO:24.62);ALT=T[chr8:29927157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29927576	+	chr8	29940363	+	.	33	29	3801846_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=3801846_2;MATENM=0;NM=2;NUMPARTS=3;REPSEQ=GGG;SCTG=c_8_29939001_29964001_338C;SPAN=12787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:139 GQ:99 PL:[120.8, 0.0, 216.5] SR:29 DR:33 LR:-120.8 LO:122.3);ALT=C[chr8:29940363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29931572	+	chr8	29940363	+	.	84	90	3801848_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=3801848_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_29939001_29964001_156C;SPAN=8791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:139 GQ:37.6 PL:[412.6, 37.6, 0.0] SR:90 DR:84 LR:-412.6 LO:412.6);ALT=C[chr8:29940363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29953044	+	chr8	29963261	+	CTTTGATTAGTTTGTCCTTTGGAGGAGCAATCGGACTGATGTTTTTGATGCTTGGATGTGCCCTTCCAATATACAACAAATACTGGCCCCTCTTTGTTCTATTTTTTTACATCCTTTCACCTATTCCATACTGCATAGCAAGAAGATTAGTGGATGATACAGATGCTATGAGTAACGCTTGTAAGGAACTTGCCATCTTTCTTACAACGGGCATTGTCGTGTCAGCTTTTGGACTCCCTATTGTATTTGCCAGAGCACATCT	3	27	3801896_1	71.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTTTGATTAGTTTGTCCTTTGGAGGAGCAATCGGACTGATGTTTTTGATGCTTGGATGTGCCCTTCCAATATACAACAAATACTGGCCCCTCTTTGTTCTATTTTTTTACATCCTTTCACCTATTCCATACTGCATAGCAAGAAGATTAGTGGATGATACAGATGCTATGAGTAACGCTTGTAAGGAACTTGCCATCTTTCTTACAACGGGCATTGTCGTGTCAGCTTTTGGACTCCCTATTGTATTTGCCAGAGCACATCT;MAPQ=60;MATEID=3801896_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_29939001_29964001_123C;SPAN=10217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:76 GQ:71.9 PL:[71.9, 0.0, 111.5] SR:27 DR:3 LR:-71.84 LO:72.33);ALT=G[chr8:29963261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29953044	+	chr8	29959412	+	.	26	11	3801895_1	73.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3801895_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TTT;SCTG=c_8_29939001_29964001_123C;SPAN=6368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:72 GQ:73.1 PL:[73.1, 0.0, 99.5] SR:11 DR:26 LR:-72.92 LO:73.18);ALT=G[chr8:29959412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29953095	+	chr8	29961815	+	.	72	0	3801898_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3801898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:29953095(+)-8:29961815(-)__8_29939001_29964001D;SPAN=8720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:95 GQ:17.3 PL:[212.0, 0.0, 17.3] SR:0 DR:72 LR:-221.5 LO:221.5);ALT=G[chr8:29961815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	29962002	+	chr8	29963261	+	.	5	15	3801935_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=3801935_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_8_29939001_29964001_123C;SPAN=1259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:81 GQ:44.3 PL:[44.3, 0.0, 149.9] SR:15 DR:5 LR:-44.08 LO:47.43);ALT=G[chr8:29963261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	30032706	+	chr8	30034642	+	.	0	7	3801826_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=3801826_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_30012501_30037501_22C;SPAN=1936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.547 LO:12.74);ALT=C[chr8:30034642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7167959	+	chr8	30145402	+	.	35	43	6301911_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=T;MAPQ=60;MATEID=6301911_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_17_7154001_7179001_15C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:50 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:43 DR:35 LR:-201.3 LO:201.3);ALT=]chr17:7167959]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	30145623	+	chr17	7167890	+	.	0	44	6301912_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6301912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_7154001_7179001_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:58 GQ:10.7 PL:[129.5, 0.0, 10.7] SR:44 DR:0 LR:-135.4 LO:135.4);ALT=A[chr17:7167890[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	30567421	+	chr8	30585043	+	TTTTGGGTACACATCCAACAT	0	10	3803881_1	22.0	.	EVDNC=ASSMB;INSERTION=TTTTGGGTACACATCCAACAT;MAPQ=60;MATEID=3803881_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_30551501_30576501_189C;SPAN=17622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:41 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:10 DR:0 LR:-21.9 LO:23.65);ALT=T[chr8:30585043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	30891489	+	chr8	30915887	+	.	3	3	3804790_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3804790_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_30894501_30919501_259C;SPAN=24398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:38 GQ:6.2 PL:[6.2, 0.0, 85.4] SR:3 DR:3 LR:-6.21 LO:10.33);ALT=G[chr8:30915887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	35383204	+	chr17	42143930	+	.	17	0	6404482_1	44.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=6404482_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:35383204(+)-17:42143930(-)__17_42140001_42165001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:42 GQ:44.9 PL:[44.9, 0.0, 54.8] SR:0 DR:17 LR:-44.74 LO:44.82);ALT=C[chr17:42143930[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	37620277	+	chr8	37623798	+	ATCTCCCAGCCATCCAGCCCCGGCTAGTGGCGGTCAGCAAAACCAAACCTGCAGACATGGTGATCGAGGCCTATGGACATGGGCAGCGCACTTTTGGCGAGAACTACGTTCAGGAACTGCTAGAAAAAGCATCAAATCCCAAA	4	23	3823205_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=ATCTCCCAGCCATCCAGCCCCGGCTAGTGGCGGTCAGCAAAACCAAACCTGCAGACATGGTGATCGAGGCCTATGGACATGGGCAGCGCACTTTTGGCGAGAACTACGTTCAGGAACTGCTAGAAAAAGCATCAAATCCCAAA;MAPQ=60;MATEID=3823205_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_8_37607501_37632501_136C;SPAN=3521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:99 GQ:52.4 PL:[52.4, 0.0, 187.7] SR:23 DR:4 LR:-52.4 LO:56.69);ALT=G[chr8:37623798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	37620277	+	chr8	37623043	+	.	23	15	3823204_1	67.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3823204_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TCTC;SCTG=c_8_37607501_37632501_136C;SPAN=2766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:116 GQ:67.7 PL:[67.7, 0.0, 212.9] SR:15 DR:23 LR:-67.6 LO:71.85);ALT=G[chr8:37623043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	37888239	+	chr8	37917421	+	CCAGGATCATCTATGACCGGAAATTCCTGATGGAGTGTCGGAACTCACCTGTGACCAAAACACCCCCAAGGGATCTGCCCACCATTCCGGGGGTCACCAGCCCTTCCAGTGATGAGCCCCCCATGGAAGCCAGCCAGAGCCACCTGCGCAATAGCCCAGAAGATAAGCGGGCGGGC	0	85	3824403_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGTGA;INSERTION=CCAGGATCATCTATGACCGGAAATTCCTGATGGAGTGTCGGAACTCACCTGTGACCAAAACACCCCCAAGGGATCTGCCCACCATTCCGGGGGTCACCAGCCCTTCCAGTGATGAGCCCCCCATGGAAGCCAGCCAGAGCCACCTGCGCAATAGCCCAGAAGATAAGCGGGCGGGC;MAPQ=60;MATEID=3824403_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_37901501_37926501_31C;SPAN=29182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:51 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:85 DR:0 LR:-250.9 LO:250.9);ALT=A[chr8:37917421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	37888239	+	chr8	37914597	+	.	69	72	3824402_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGGTA;MAPQ=60;MATEID=3824402_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_37901501_37926501_31C;SPAN=26358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:53 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:72 DR:69 LR:-356.5 LO:356.5);ALT=A[chr8:37914597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	37914782	+	chr8	37917421	+	.	3	8	3824447_1	12.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGTGA;MAPQ=60;MATEID=3824447_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_37901501_37926501_31C;SPAN=2639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:8 DR:3 LR:-12.74 LO:22.52);ALT=A[chr8:37917421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	38027436	+	chr8	38033793	+	AAATTGATCAATGCTTCTTAAAAAGCCTATAAGTGTCCTTCCATCTCGAAGCAGAACCAAGTGCTTTT	0	20	3824673_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AAATTGATCAATGCTTCTTAAAAAGCCTATAAGTGTCCTTCCATCTCGAAGCAGAACCAAGTGCTTTT;MAPQ=60;MATEID=3824673_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_38024001_38049001_397C;SPAN=6357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:85 GQ:43.1 PL:[43.1, 0.0, 161.9] SR:20 DR:0 LR:-42.99 LO:46.94);ALT=C[chr8:38033793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	38029595	+	chr8	38033892	+	.	10	0	3824681_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3824681_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:38029595(+)-8:38033892(-)__8_38024001_38049001D;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:0 DR:10 LR:-7.543 LO:19.68);ALT=T[chr8:38033892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	38089377	+	chr8	38090503	+	.	4	4	3824971_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3824971_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_38073001_38098001_308C;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:79 GQ:1.7 PL:[1.7, 0.0, 189.8] SR:4 DR:4 LR:-1.704 LO:13.19);ALT=G[chr8:38090503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	38758964	+	chr8	38775424	+	.	0	7	3827566_1	13.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3827566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_38734501_38759501_108C;SPAN=16460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:37 GQ:13.1 PL:[13.1, 0.0, 75.8] SR:7 DR:0 LR:-13.08 LO:15.67);ALT=G[chr8:38775424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	39232074	+	chr8	39387229	+	T	46	32	3829053_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=3829053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_39371501_39396501_56C;SPAN=155155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:21 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:32 DR:46 LR:-188.1 LO:188.1);ALT=G[chr8:39387229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	40289707	+	chr8	40296198	+	.	76	59	3832045_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAAAAAATACACAGGA;MAPQ=60;MATEID=3832045_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_8_40278001_40303001_55C;SPAN=6491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:33 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:59 DR:76 LR:-303.7 LO:303.7);ALT=A[chr8:40296198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	40817287	-	chr8	40818561	+	.	12	0	3833122_1	24.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3833122_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:40817287(-)-8:40818561(-)__8_40792501_40817501D;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:57 GQ:24.2 PL:[24.2, 0.0, 113.3] SR:0 DR:12 LR:-24.17 LO:27.5);ALT=[chr8:40818561[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	41348484	+	chr8	41355027	+	.	23	27	3834720_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=3834720_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_41331501_41356501_163C;SPAN=6543;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:100 GQ:99 PL:[108.2, 0.0, 134.6] SR:27 DR:23 LR:-108.2 LO:108.4);ALT=G[chr8:41355027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	41906816	+	chr8	41909440	+	.	8	0	3836536_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3836536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:41906816(+)-8:41909440(-)__8_41895001_41920001D;SPAN=2624;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=T[chr8:41909440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42129724	+	chr8	42146150	+	.	0	8	3837280_1	14.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3837280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_42115501_42140501_382C;SPAN=16426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:8 DR:0 LR:-13.95 LO:17.59);ALT=G[chr8:42146150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42190485	+	chr8	42194353	+	.	95	0	3837614_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CCTGTAATCCCAGCTACTCGGGAGGCTGAGGCAGGAGAATCGCTTGAACCCGGGAGGCAGAGGTTGCAGTGAGCCGAGATCGTGCCATTGCACTCC;MAPQ=60;MATEID=3837614_2;MATENM=2;NM=4;NUMPARTS=2;SCTG=c_8_42189001_42214001_113C;SPAN=3868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:5 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:0 DR:95 LR:-280.6 LO:280.6);ALT=C[chr8:42194353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42249488	+	chr8	42256228	+	.	19	0	3837824_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3837824_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:42249488(+)-8:42256228(-)__8_42238001_42263001D;SPAN=6740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:99 GQ:35.9 PL:[35.9, 0.0, 204.2] SR:0 DR:19 LR:-35.9 LO:42.68);ALT=C[chr8:42256228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42396848	+	chr8	42401612	+	.	15	3	3838186_1	37.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3838186_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_42385001_42410001_330C;SPAN=4764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:70 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:3 DR:15 LR:-37.15 LO:40.17);ALT=C[chr8:42401612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42396882	+	chr8	42403796	+	.	12	0	3838187_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3838187_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:42396882(+)-8:42403796(-)__8_42385001_42410001D;SPAN=6914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:0 DR:12 LR:-24.71 LO:27.71);ALT=C[chr8:42403796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42401750	+	chr8	42403797	+	.	0	13	3838207_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=3838207_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_42385001_42410001_362C;SPAN=2047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:79 GQ:21.5 PL:[21.5, 0.0, 170.0] SR:13 DR:0 LR:-21.51 LO:28.24);ALT=G[chr8:42403797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	42740058	+	chr11	82567909	-	.	11	0	3840295_1	23.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3840295_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:42740058(+)-11:82567909(+)__8_42728001_42753001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:48 GQ:23.3 PL:[23.3, 0.0, 92.6] SR:0 DR:11 LR:-23.31 LO:25.67);ALT=T]chr11:82567909];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	42752331	+	chr8	42761315	+	.	0	14	3840345_1	35.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=3840345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_42728001_42753001_402C;SPAN=8984;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:39 GQ:35.6 PL:[35.6, 0.0, 58.7] SR:14 DR:0 LR:-35.65 LO:35.96);ALT=G[chr8:42761315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	52406453	-	chr11	62899264	+	.	19	19	4884340_1	95.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=GTTCTCTGTATTTCCTGGATTTGAATGTTGGCCTGCCT;MAPQ=60;MATEID=4884340_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_11_62891501_62916501_103C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:19 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:19 DR:19 LR:-95.72 LO:95.72);ALT=[chr11:62899264[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	52773817	+	chr8	52811511	+	.	20	0	3858194_1	52.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=3858194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:52773817(+)-8:52811511(-)__8_52797501_52822501D;SPAN=37694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:52 GQ:52.1 PL:[52.1, 0.0, 71.9] SR:0 DR:20 LR:-51.93 LO:52.15);ALT=A[chr8:52811511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	56675627	+	chr8	56685827	+	.	18	0	3869239_1	38.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=3869239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:56675627(+)-8:56685827(-)__8_56668501_56693501D;SPAN=10200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:77 GQ:38.6 PL:[38.6, 0.0, 147.5] SR:0 DR:18 LR:-38.56 LO:42.19);ALT=C[chr8:56685827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	56792663	+	chr8	56854413	+	.	12	15	3869829_1	56.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=3869829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_56840001_56865001_53C;SPAN=61750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:48 GQ:56.3 PL:[56.3, 0.0, 59.6] SR:15 DR:12 LR:-56.32 LO:56.32);ALT=G[chr8:56854413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	56963762	+	chr14	53174015	-	.	12	0	5744240_1	26.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5744240_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:56963762(+)-14:53174015(+)__14_53165001_53190001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:51 GQ:26 PL:[26.0, 0.0, 95.3] SR:0 DR:12 LR:-25.8 LO:28.16);ALT=G]chr14:53174015];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	57124431	+	chr8	57127154	+	.	9	0	3870879_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3870879_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:57124431(+)-8:57127154(-)__8_57109501_57134501D;SPAN=2723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:94 GQ:4.4 PL:[4.4, 0.0, 222.2] SR:0 DR:9 LR:-4.242 LO:17.27);ALT=C[chr8:57127154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	57124431	+	chr8	57129888	+	.	12	0	3870880_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3870880_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:57124431(+)-8:57129888(-)__8_57109501_57134501D;SPAN=5457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:0 DR:12 LR:-16.31 LO:25.12);ALT=C[chr8:57129888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	57124433	+	chr8	57128950	+	.	18	0	3870881_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3870881_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:57124433(+)-8:57128950(-)__8_57109501_57134501D;SPAN=4517;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:89 GQ:35.3 PL:[35.3, 0.0, 180.5] SR:0 DR:18 LR:-35.31 LO:40.89);ALT=C[chr8:57128950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	57125468	+	chr8	57127155	+	.	3	3	3870887_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3870887_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_57109501_57134501_46C;SPAN=1687;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:70 GQ:0.8 PL:[0.8, 0.0, 169.1] SR:3 DR:3 LR:-0.8413 LO:11.21);ALT=G[chr8:57127155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	58126666	+	chr8	58122281	+	.	7	14	3874007_1	8.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GGAAGGC;MAPQ=60;MATEID=3874007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_58114001_58139001_323C;SPAN=4385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:202 GQ:8.2 PL:[8.2, 0.0, 480.2] SR:14 DR:7 LR:-7.992 LO:36.31);ALT=]chr8:58126666]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	63939825	+	chr8	63948214	+	CATTAATAGATTTGAAAAGTATTTCATAGTCTTTCTCTGTAAGATCCAG	0	11	3888643_1	24.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CATTAATAGATTTGAAAAGTATTTCATAGTCTTTCTCTGTAAGATCCAG;MAPQ=60;MATEID=3888643_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_63945001_63970001_118C;SPAN=8389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:11 DR:0 LR:-24.12 LO:26.03);ALT=C[chr8:63948214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	63948330	+	chr8	63951218	+	.	0	11	3888653_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=3888653_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_63945001_63970001_182C;SPAN=2888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:82 GQ:14.3 PL:[14.3, 0.0, 182.6] SR:11 DR:0 LR:-14.1 LO:22.83);ALT=C[chr8:63951218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	71487243	+	chr8	71495399	+	.	7	5	3909529_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=3909529_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_71491001_71516001_221C;SPAN=8156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:5 DR:7 LR:-26.29 LO:27.14);ALT=G[chr8:71495399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	71510493	+	chr8	71520312	+	TTGCTGGGAGGGTGACATTGTACTGAAGAGTAACAAAAATGATAGAAGCTTTTGCCGTTAT	0	27	3909602_1	78.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTGCTGGGAGGGTGACATTGTACTGAAGAGTAACAAAAATGATAGAAGCTTTTGCCGTTAT;MAPQ=60;MATEID=3909602_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_71515501_71540501_346C;SPAN=9819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:40 GQ:18.8 PL:[78.2, 0.0, 18.8] SR:27 DR:0 LR:-80.33 LO:80.33);ALT=G[chr8:71520312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	71583571	+	chr8	71584644	+	.	84	72	3909790_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATGATCTCATTTTTTT;MAPQ=60;MATEID=3909790_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_71564501_71589501_137C;SPAN=1073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:52 GQ:33 PL:[363.0, 33.0, 0.0] SR:72 DR:84 LR:-363.1 LO:363.1);ALT=T[chr8:71584644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	72214752	+	chr8	72217809	+	.	45	33	3911452_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGCTGA;MAPQ=60;MATEID=3911452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_72201501_72226501_151C;SPAN=3057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:71 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:33 DR:45 LR:-205.9 LO:205.9);ALT=A[chr8:72217809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	73611044	-	chr8	73612655	+	.	8	0	3915126_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=3915126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:73611044(-)-8:73612655(-)__8_73598001_73623001D;SPAN=1611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr8:73612655[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	73787775	+	chr8	73793824	+	.	62	57	3915763_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGCAAATCTT;MAPQ=60;MATEID=3915763_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_73769501_73794501_251C;SPAN=6049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:102 DP:127 GQ:5.3 PL:[302.3, 0.0, 5.3] SR:57 DR:62 LR:-319.7 LO:319.7);ALT=T[chr8:73793824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	74742716	+	chr8	74791042	+	.	13	0	3918423_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3918423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:74742716(+)-8:74791042(-)__8_74774001_74799001D;SPAN=48326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.66 LO:29.98);ALT=G[chr8:74791042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	74868295	+	chr8	74884310	+	.	24	0	3918908_1	66.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=3918908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:74868295(+)-8:74884310(-)__8_74872001_74897001D;SPAN=16015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:46 GQ:43.7 PL:[66.8, 0.0, 43.7] SR:0 DR:24 LR:-66.99 LO:66.99);ALT=G[chr8:74884310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	74884147	-	chr18	4459288	+	.	19	0	3918952_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3918952_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:74884147(-)-18:4459288(-)__8_74872001_74897001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:40 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:0 DR:19 LR:-51.91 LO:51.91);ALT=[chr18:4459288[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	74884310	-	chr15	41849171	+	.	18	0	3918954_1	47.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3918954_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:74884310(-)-15:41849171(-)__8_74872001_74897001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:46 GQ:47 PL:[47.0, 0.0, 63.5] SR:0 DR:18 LR:-46.96 LO:47.11);ALT=[chr15:41849171[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr20	17550857	+	chr8	74896721	+	.	9	10	3918988_1	39.0	.	DISC_MAPQ=7;EVDNC=ASDIS;HOMSEQ=GGCGAAGATGG;MAPQ=21;MATEID=3918988_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_74872001_74897001_59C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:10 DR:9 LR:-39.0 LO:39.93);ALT=]chr20:17550857]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	74903725	+	chr8	74917029	+	.	11	0	3919437_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3919437_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:74903725(+)-8:74917029(-)__8_74896501_74921501D;SPAN=13304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:89 GQ:12.2 PL:[12.2, 0.0, 203.6] SR:0 DR:11 LR:-12.2 LO:22.41);ALT=T[chr8:74917029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	75362871	+	chr8	75367000	+	CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA	34	56	3920406_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTACAATGTAATAACATTGCCAAATAATTATAATGCCAAATATAATGATA;MAPQ=60;MATEID=3920406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_75337501_75362501_106C;SPAN=4129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:0 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:56 DR:34 LR:-208.0 LO:208.0);ALT=A[chr8:75367000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	75516588	+	chr12	53846160	-	.	17	68	5195584_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TCCCCTTTTCCCCTCAGTCGCCTCGCGCCTGCAG;MAPQ=59;MATEID=5195584_2;MATENM=1;NM=3;NUMPARTS=2;SCTG=c_12_53826501_53851501_317C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:128 GQ:64.4 PL:[245.9, 0.0, 64.4] SR:68 DR:17 LR:-251.8 LO:251.8);ALT=A]chr12:53846160];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	80518566	+	chr19	39037385	+	AAAGAAAATGATAAAACAAATGTGATGCAGGGTGCGTCACGTGCCTGTAATCCCAGCACTTTGGGAGGCCGAGGCCAGAGGATCTCTTGAGCCCAGC	0	70	6811710_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=AAAGAAAATGATAAAACAAATGTGATGCAGGGTGCGTCACGTGCCTGTAATCCCAGCACTTTGGGAGGCCGAGGCCAGAGGATCTCTTGAGCCCAGC;MAPQ=60;MATEID=6811710_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_19_39028501_39053501_275C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:28 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:70 DR:0 LR:-208.0 LO:208.0);ALT=G[chr19:39037385[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	80976830	+	chr8	81083658	+	.	6	4	3935022_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=3935022_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_81070501_81095501_255C;SPAN=106828;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:4 DR:6 LR:-16.11 LO:18.33);ALT=T[chr8:81083658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	81133436	+	chr8	81134538	-	.	9	0	3935176_1	5.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=3935176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:81133436(+)-8:81134538(+)__8_81119501_81144501D;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:0 DR:9 LR:-4.784 LO:17.36);ALT=C]chr8:81134538];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	82045018	+	chr8	82046625	+	TTACGT	70	36	3937783_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;INSERTION=TTACGT;MAPQ=60;MATEID=3937783_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_8_82026001_82051001_324C;SPAN=1607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:59 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:36 DR:70 LR:-267.4 LO:267.4);ALT=G[chr8:82046625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	82192863	+	chr11	59549161	-	.	58	0	4874864_1	99.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=4874864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:82192863(+)-11:59549161(+)__11_59535001_59560001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:43 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:58 LR:-171.6 LO:171.6);ALT=G]chr11:59549161];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	82627166	+	chr8	82633462	+	.	10	0	3939612_1	7.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=3939612_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:82627166(+)-8:82633462(-)__8_82614001_82639001D;SPAN=6296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:96 GQ:7.1 PL:[7.1, 0.0, 224.9] SR:0 DR:10 LR:-7.001 LO:19.58);ALT=T[chr8:82633462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	83269755	+	chr8	83295603	+	.	41	27	3941214_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTTATCT;MAPQ=60;MATEID=3941214_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_83251001_83276001_12C;SPAN=25848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:29 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:27 DR:41 LR:-151.8 LO:151.8);ALT=T[chr8:83295603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	97244179	+	chr8	97247739	+	.	28	0	3982351_1	65.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=3982351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:97244179(+)-8:97247739(-)__8_97240501_97265501D;SPAN=3560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:100 GQ:65.3 PL:[65.3, 0.0, 177.5] SR:0 DR:28 LR:-65.34 LO:68.2);ALT=T[chr8:97247739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	97274448	+	chr8	97285524	+	.	0	12	3982290_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=3982290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_97265001_97290001_118C;SPAN=11076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:112 GQ:9.5 PL:[9.5, 0.0, 260.3] SR:12 DR:0 LR:-9.269 LO:23.65);ALT=G[chr8:97285524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	97657630	+	chr8	97797090	+	.	23	8	3983784_1	77.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3983784_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_97779501_97804501_41C;SPAN=139460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:44 GQ:27.8 PL:[77.3, 0.0, 27.8] SR:8 DR:23 LR:-78.37 LO:78.37);ALT=G[chr8:97797090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98657115	+	chr8	98673300	+	.	6	34	3986120_1	98.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=3986120_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_98661501_98686501_44C;SPAN=16185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:49 GQ:19.7 PL:[98.9, 0.0, 19.7] SR:34 DR:6 LR:-101.9 LO:101.9);ALT=A[chr8:98673300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98673401	+	chr8	98698894	+	.	3	8	3986207_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=3986207_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_98686001_98711001_335C;SPAN=25493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:8 DR:3 LR:-18.6 LO:20.81);ALT=G[chr8:98698894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98699835	+	chr8	98703179	+	GATTCTCATCTAAATGTTCAAGTTAGCAACTTTAAATCTGGAAAAGGAGATTCTACACTTCAG	3	13	3986271_1	31.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GATTCTCATCTAAATGTTCAAGTTAGCAACTTTAAATCTGGAAAAGGAGATTCTACACTTCAG;MAPQ=60;MATEID=3986271_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_98686001_98711001_276C;SPAN=3344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:67 GQ:31.4 PL:[31.4, 0.0, 130.4] SR:13 DR:3 LR:-31.36 LO:34.83);ALT=T[chr8:98703179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98703417	+	chr8	98718854	+	GTCTACTGCTGAGCCAGTTTCTCAGTCTACCACTTCTGATTATCAGTGGGATGTTAGCCGTAATCAACCCTATATCGATGATGAATGGTCTGGGTTAA	0	63	3986325_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GTCTACTGCTGAGCCAGTTTCTCAGTCTACCACTTCTGATTATCAGTGGGATGTTAGCCGTAATCAACCCTATATCGATGATGAATGGTCTGGGTTAA;MAPQ=60;MATEID=3986325_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_98710501_98735501_151C;SPAN=15437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:62 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:63 DR:0 LR:-184.8 LO:184.8);ALT=G[chr8:98718854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98703417	+	chr8	98711981	+	.	4	20	3986324_1	65.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3986324_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_8_98710501_98735501_151C;SPAN=8564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:20 DR:4 LR:-65.7 LO:65.7);ALT=G[chr8:98711981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98712080	+	chr8	98718854	+	.	0	40	3986329_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=3986329_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_8_98710501_98735501_151C;SPAN=6774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:101 GQ:99 PL:[104.9, 0.0, 137.9] SR:40 DR:0 LR:-104.7 LO:105.0);ALT=A[chr8:98718854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	98731417	+	chr8	98735105	+	.	0	9	3986397_1	5.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=3986397_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_98710501_98735501_204C;SPAN=3688;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:9 DR:0 LR:-5.326 LO:17.45);ALT=G[chr8:98735105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	99054108	+	chr8	99057733	+	.	9	0	3987710_1	0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=3987710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:99054108(+)-8:99057733(-)__8_99053501_99078501D;SPAN=3625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:796 GQ:99 PL:[0.0, 185.6, 2304.0] SR:0 DR:9 LR:185.9 LO:8.866);ALT=T[chr8:99057733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	99055005	+	chr8	99057170	+	.	0	121	3987717_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=3987717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_99053501_99078501_129C;SPAN=2165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:121 DP:1080 GQ:99 PL:[107.0, 0.0, 2517.0] SR:121 DR:0 LR:-106.8 LO:241.0);ALT=T[chr8:99057170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	99055064	+	chr8	99057733	+	.	34	0	3987718_1	0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=3987718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:99055064(+)-8:99057733(-)__8_99053501_99078501D;SPAN=2669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:34 DP:814 GQ:99 PL:[0.0, 107.9, 2192.0] SR:0 DR:34 LR:108.3 LO:52.63);ALT=G[chr8:99057733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	100890495	+	chr8	100899718	+	.	0	162	3992788_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=35;MATEID=3992788_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_100891001_100916001_276C;SPAN=9223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:162 DP:64 GQ:43.6 PL:[478.6, 43.6, 0.0] SR:162 DR:0 LR:-478.6 LO:478.6);ALT=T[chr8:100899718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	100899897	+	chr8	100905864	+	.	45	0	3992816_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=3992816_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:100899897(+)-8:100905864(-)__8_100891001_100916001D;SPAN=5967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:148 GQ:99 PL:[108.5, 0.0, 250.4] SR:0 DR:45 LR:-108.4 LO:111.6);ALT=G[chr8:100905864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	100904324	+	chr8	100905793	+	.	61	0	3992830_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=3992830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:100904324(+)-8:100905793(-)__8_100891001_100916001D;SPAN=1469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:79 GQ:11.6 PL:[179.9, 0.0, 11.6] SR:0 DR:61 LR:-188.7 LO:188.7);ALT=A[chr8:100905793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101162981	+	chr8	101164049	+	.	46	0	3993692_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=3993692_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101162981(+)-8:101164049(-)__8_101160501_101185501D;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:104 GQ:99 PL:[123.8, 0.0, 127.1] SR:0 DR:46 LR:-123.7 LO:123.7);ALT=C[chr8:101164049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101162989	+	chr8	101165521	+	.	47	0	3993693_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=3993693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101162989(+)-8:101165521(-)__8_101160501_101185501D;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:100 GQ:99 PL:[128.0, 0.0, 114.8] SR:0 DR:47 LR:-128.1 LO:128.1);ALT=G[chr8:101165521[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101164144	+	chr8	101165522	+	.	3	57	3993699_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;MAPQ=60;MATEID=3993699_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_101160501_101185501_0C;SPAN=1378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:101 GQ:71.9 PL:[170.9, 0.0, 71.9] SR:57 DR:3 LR:-172.8 LO:172.8);ALT=T[chr8:101165522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101300497	+	chr8	101322095	+	.	24	10	3994237_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=3994237_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_101307501_101332501_313C;SPAN=21598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:10 DR:24 LR:-99.02 LO:99.02);ALT=T[chr8:101322095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101717290	+	chr8	101718883	+	.	14	0	3995931_1	22.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=3995931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101717290(+)-8:101718883(-)__8_101699501_101724501D;SPAN=1593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:88 GQ:22.4 PL:[22.4, 0.0, 190.7] SR:0 DR:14 LR:-22.37 LO:30.18);ALT=A[chr8:101718883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101719249	+	chr8	101721686	+	.	23	0	3995953_1	47.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=3995953_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101719249(+)-8:101721686(-)__8_101699501_101724501D;SPAN=2437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:105 GQ:47.6 PL:[47.6, 0.0, 206.0] SR:0 DR:23 LR:-47.48 LO:53.16);ALT=A[chr8:101721686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101721988	+	chr8	101724878	+	.	12	0	3995976_1	26.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=3995976_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101721988(+)-8:101724878(-)__8_101699501_101724501D;SPAN=2890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:48 GQ:26.6 PL:[26.6, 0.0, 89.3] SR:0 DR:12 LR:-26.61 LO:28.53);ALT=C[chr8:101724878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101727834	+	chr8	101730312	+	.	8	0	3995494_1	0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=3995494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101727834(+)-8:101730312(-)__8_101724001_101749001D;SPAN=2478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=T[chr8:101730312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101727844	+	chr8	101730007	+	.	8	0	3995495_1	1.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=3995495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101727844(+)-8:101730007(-)__8_101724001_101749001D;SPAN=2163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=A[chr8:101730007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101730118	+	chr8	101733619	+	CGGAGCGTGCTTTGGACACCATGAATTTTGATGTTATAAAGGGCAAGCCAGTACGCATCATGTGGTCTCAGCGTGATCCATCACTTCGCAAAAGTGGAGTAGGCAACATATTCATTAAAAATCTGGACAAATCCATTGATAATAAAGCACTGTATGATACATTTTCTGCTTTTGGTAACATCCTTTCATGTA	2	47	3995507_1	99.0	.	DISC_MAPQ=44;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=CGGAGCGTGCTTTGGACACCATGAATTTTGATGTTATAAAGGGCAAGCCAGTACGCATCATGTGGTCTCAGCGTGATCCATCACTTCGCAAAAGTGGAGTAGGCAACATATTCATTAAAAATCTGGACAAATCCATTGATAATAAAGCACTGTATGATACATTTTCTGCTTTTGGTAACATCCTTTCATGTA;MAPQ=60;MATEID=3995507_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_101724001_101749001_81C;SPAN=3501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:86 GQ:75.8 PL:[131.9, 0.0, 75.8] SR:47 DR:2 LR:-132.6 LO:132.6);ALT=T[chr8:101733619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101730509	+	chr8	101733619	+	.	24	35	3995508_1	99.0	.	DISC_MAPQ=35;EVDNC=TSI_L;HOMSEQ=G;MAPQ=51;MATEID=3995508_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_101724001_101749001_81C;SPAN=3110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:83 GQ:37.1 PL:[162.5, 0.0, 37.1] SR:35 DR:24 LR:-166.6 LO:166.6);ALT=C[chr8:101733619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101905126	+	chr9	100558852	-	.	8	0	4354116_1	16.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=4354116_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101905126(+)-9:100558852(+)__9_100548001_100573001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:37 GQ:16.4 PL:[16.4, 0.0, 72.5] SR:0 DR:8 LR:-16.38 LO:18.44);ALT=A]chr9:100558852];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr8	101961128	+	chr8	101964156	+	.	106	0	3996479_1	99.0	.	DISC_MAPQ=5;EVDNC=DSCRD;IMPRECISE;MAPQ=5;MATEID=3996479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:101961128(+)-8:101964156(-)__8_101944501_101969501D;SPAN=3028;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:96 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:0 DR:106 LR:-313.6 LO:313.6);ALT=T[chr8:101964156[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	101964157	-	chr10	23425817	+	.	31	15	4543359_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCGCCACCACCCACTCCGGACACAG;MAPQ=60;MATEID=4543359_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_23422001_23447001_75C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:54 GQ:18.5 PL:[110.9, 0.0, 18.5] SR:15 DR:31 LR:-114.4 LO:114.4);ALT=[chr10:23425817[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	103664626	+	chr8	103667793	+	.	19	10	4001695_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4001695_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_103659501_103684501_283C;SPAN=3167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:69 GQ:50.6 PL:[50.6, 0.0, 116.6] SR:10 DR:19 LR:-50.63 LO:52.07);ALT=C[chr8:103667793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	103855975	+	chr8	103870241	+	.	3	6	4002488_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4002488_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_103855501_103880501_329C;SPAN=14266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:91 GQ:4.5 PL:[0.0, 4.5, 227.7] SR:6 DR:3 LR:4.848 LO:10.5);ALT=A[chr8:103870241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	104153286	+	chr8	104225146	+	.	3	2	4003688_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4003688_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_104223001_104248001_44C;SPAN=71860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:59 GQ:0.5 PL:[0.5, 0.0, 142.4] SR:2 DR:3 LR:-0.5205 LO:9.318);ALT=G[chr8:104225146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	104414284	+	chr8	104415391	+	.	0	6	4004073_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4004073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_104394501_104419501_305C;SPAN=1107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:97 GQ:6.3 PL:[0.0, 6.3, 247.5] SR:6 DR:0 LR:6.474 LO:10.33);ALT=T[chr8:104415391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	104427766	+	chr8	104432490	+	.	11	0	4004248_1	13.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4004248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:104427766(+)-8:104432490(-)__8_104419001_104444001D;SPAN=4724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:0 DR:11 LR:-13.55 LO:22.7);ALT=A[chr8:104432490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	107008900	-	chr9	15365423	+	.	7	29	4011133_1	92.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=TTCTCCAAGTCCCCACCCAA;MAPQ=15;MATEID=4011133_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_8_106991501_107016501_7C;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:47 GQ:20.3 PL:[92.9, 0.0, 20.3] SR:29 DR:7 LR:-95.43 LO:95.43);ALT=[chr9:15365423[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	108348501	+	chr8	108359166	+	.	0	14	4014565_1	21.0	.	EVDNC=ASSMB;HOMSEQ=GTACCT;MAPQ=60;MATEID=4014565_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_108339001_108364001_51C;SPAN=10665;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:92 GQ:21.5 PL:[21.5, 0.0, 199.7] SR:14 DR:0 LR:-21.29 LO:29.89);ALT=T[chr8:108359166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109226945	+	chr8	109228639	+	.	4	26	4016964_1	70.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=4016964_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_109221001_109246001_190C;SPAN=1694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:95 GQ:70.1 PL:[70.1, 0.0, 159.2] SR:26 DR:4 LR:-69.99 LO:71.95);ALT=C[chr8:109228639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109229689	+	chr8	109240496	+	.	3	6	4016969_1	8.0	.	DISC_MAPQ=41;EVDNC=ASDIS;MAPQ=60;MATEID=4016969_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_109221001_109246001_254C;SPAN=10807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:6 DR:3 LR:-8.035 LO:17.94);ALT=T[chr8:109240496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109252328	+	chr8	109254028	+	.	4	5	4017306_1	3.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4017306_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_109245501_109270501_336C;SPAN=1700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:5 DR:4 LR:-3.429 LO:17.14);ALT=C[chr8:109254028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109252371	+	chr8	109260871	+	.	110	0	4017307_1	99.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=4017307_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:109252371(+)-8:109260871(-)__8_109245501_109270501D;SPAN=8500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:90 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:110 LR:-326.8 LO:326.8);ALT=A[chr8:109260871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109254166	+	chr8	109260881	+	.	143	0	4017313_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=4017313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:109254166(+)-8:109260881(-)__8_109245501_109270501D;SPAN=6715;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:163 GQ:34 PL:[462.1, 34.0, 0.0] SR:0 DR:143 LR:-464.5 LO:464.5);ALT=A[chr8:109260881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	109462165	+	chr8	109465290	+	TTTGGATCATATATGAACAGGTGATGATTGCAGCACTAGACTATGGTCGGGATGACTTGGCATT	0	9	4017708_1	9.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTGGATCATATATGAACAGGTGATGATTGCAGCACTAGACTATGGTCGGGATGACTTGGCATT;MAPQ=60;MATEID=4017708_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_109441501_109466501_144C;SPAN=3125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:9 DR:0 LR:-9.119 LO:18.15);ALT=A[chr8:109465290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110346705	+	chr8	110348356	+	.	31	33	4020045_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4020045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110323501_110348501_3C;SPAN=1651;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:128 GQ:99 PL:[130.4, 0.0, 179.9] SR:33 DR:31 LR:-130.4 LO:130.8);ALT=T[chr8:110348356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110346718	+	chr8	110351547	+	.	31	0	4020047_1	84.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4020047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:110346718(+)-8:110351547(-)__8_110323501_110348501D;SPAN=4829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:66 GQ:74.6 PL:[84.5, 0.0, 74.6] SR:0 DR:31 LR:-84.47 LO:84.47);ALT=T[chr8:110351547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110348433	+	chr8	110351548	+	.	2	77	4020260_1	99.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4020260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110348001_110373001_258C;SPAN=3115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:118 GQ:60.5 PL:[225.5, 0.0, 60.5] SR:77 DR:2 LR:-230.8 LO:230.8);ALT=G[chr8:110351548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110351619	+	chr8	110352715	+	.	0	72	4020273_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AAG;MAPQ=60;MATEID=4020273_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110348001_110373001_152C;SPAN=1096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:111 GQ:59.3 PL:[207.8, 0.0, 59.3] SR:72 DR:0 LR:-212.0 LO:212.0);ALT=G[chr8:110352715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	110352792	+	chr8	110355632	+	.	0	40	4020281_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=41;MATEID=4020281_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_110348001_110373001_79C;SPAN=2840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:100 GQ:99 PL:[104.9, 0.0, 137.9] SR:40 DR:0 LR:-104.9 LO:105.2);ALT=G[chr8:110355632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	112294052	+	chr8	112297140	+	.	108	86	4024740_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4024740_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_112283501_112308501_73C;SPAN=3088;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:155 DP:41 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:86 DR:108 LR:-458.8 LO:458.8);ALT=G[chr8:112297140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	123212527	-	chr8	123213699	+	.	8	0	4053717_1	2.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4053717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:123212527(-)-8:123213699(-)__8_123210501_123235501D;SPAN=1172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=[chr8:123213699[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	123966310	+	chr8	123964494	+	.	12	21	4055926_1	43.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=4055926_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_123945501_123970501_344C;SPAN=1816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:156 GQ:43.7 PL:[43.7, 0.0, 334.1] SR:21 DR:12 LR:-43.56 LO:56.63);ALT=]chr8:123966310]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	123964496	-	chr8	123966232	+	.	5	14	4055927_1	13.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4055927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_123945501_123970501_51C;SPAN=1736;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:168 GQ:13.9 PL:[13.9, 0.0, 393.5] SR:14 DR:5 LR:-13.9 LO:35.47);ALT=[chr8:123966232[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	124251402	+	chr8	124253526	+	.	10	0	4057029_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4057029_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:124251402(+)-8:124253526(-)__8_124239501_124264501D;SPAN=2124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.918 LO:19.39);ALT=A[chr8:124253526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	124263542	+	chr8	124268078	+	.	8	2	4057071_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTG;MAPQ=60;MATEID=4057071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_124239501_124264501_269C;SPAN=4536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:2 DR:8 LR:-19.19 LO:22.57);ALT=G[chr8:124268078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	124327052	+	chr19	21890756	+	.	6	11	4057122_1	48.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=GCCCGGCAGCCGCCCCGTCTGGGAAGTGAGGAGCGTCTCCGCC;MAPQ=60;MATEID=4057122_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_124313001_124338001_93C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:28 GQ:18.8 PL:[48.5, 0.0, 18.8] SR:11 DR:6 LR:-49.21 LO:49.21);ALT=C[chr19:21890756[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	124392917	+	chr8	124408426	+	.	0	9	4057281_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4057281_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_124386501_124411501_64C;SPAN=15509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:91 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:9 DR:0 LR:-5.055 LO:17.41);ALT=C[chr8:124408426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	124874943	+	chr20	21894248	+	.	15	0	6956439_1	41.0	.	DISC_MAPQ=11;EVDNC=DSCRD;IMPRECISE;MAPQ=11;MATEID=6956439_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:124874943(+)-20:21894248(-)__20_21878501_21903501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:29 GQ:28.4 PL:[41.6, 0.0, 28.4] SR:0 DR:15 LR:-41.78 LO:41.78);ALT=C[chr20:21894248[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	125528284	+	chr8	125551265	+	.	15	0	4060914_1	35.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=4060914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:125528284(+)-8:125551265(-)__8_125538001_125563001D;SPAN=22981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:53 GQ:35.3 PL:[35.3, 0.0, 91.4] SR:0 DR:15 LR:-35.16 LO:36.62);ALT=A[chr8:125551265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	125551262	-	chr10	64981924	+	.	45	0	4060953_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4060953_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:125551262(-)-10:64981924(-)__8_125538001_125563001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:0 DR:45 LR:-141.9 LO:141.9);ALT=[chr10:64981924[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	125551528	+	chr8	125555326	+	.	121	37	4060956_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4060956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_125538001_125563001_3C;SPAN=3798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:119 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:37 DR:121 LR:-422.5 LO:422.5);ALT=G[chr8:125555326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	125555522	+	chr8	125559239	+	.	0	43	4060966_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=35;MATEID=4060966_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_125538001_125563001_301C;SPAN=3717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:111 GQ:99 PL:[112.1, 0.0, 155.0] SR:43 DR:0 LR:-111.9 LO:112.3);ALT=T[chr8:125559239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	126104200	+	chr8	126114290	+	.	16	3	4062617_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4062617_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_126101501_126126501_279C;SPAN=10090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:86 GQ:56 PL:[56.0, 0.0, 151.7] SR:3 DR:16 LR:-55.92 LO:58.42);ALT=G[chr8:126114290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	126595129	+	chr8	126601135	+	.	104	46	4064665_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACTCACA;MAPQ=60;MATEID=4064665_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_8_126591501_126616501_153C;SPAN=6006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:156 GQ:19 PL:[415.9, 19.0, 0.0] SR:46 DR:104 LR:-426.4 LO:426.4);ALT=A[chr8:126601135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	127192205	+	chr8	127194572	+	T	47	42	4065851_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=T;MAPQ=60;MATEID=4065851_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_127179501_127204501_144C;SPAN=2367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:60 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:42 DR:47 LR:-224.5 LO:224.5);ALT=C[chr8:127194572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	134878295	+	chr8	135682508	+	.	12	0	4090404_1	24.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=4090404_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:134878295(+)-8:135682508(-)__8_135681001_135706001D;SPAN=804213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:56 GQ:24.5 PL:[24.5, 0.0, 110.3] SR:0 DR:12 LR:-24.44 LO:27.6);ALT=T[chr8:135682508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	135683093	+	chr8	134878854	+	.	9	0	4090405_1	18.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=4090405_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:134878854(-)-8:135683093(+)__8_135681001_135706001D;SPAN=804239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=]chr8:135683093]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	134972222	-	chr18	57070970	+	.	45	0	6641939_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6641939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:134972222(-)-18:57070970(-)__18_57060501_57085501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:33 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=[chr18:57070970[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr8	135082929	+	chr8	135089016	+	.	30	11	4088921_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CATTCTTCAACATTTT;MAPQ=60;MATEID=4088921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_135068501_135093501_317C;SPAN=6087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:36 DP:499 GQ:16.2 PL:[0.0, 16.2, 1244.0] SR:11 DR:30 LR:16.36 LO:64.47);ALT=T[chr8:135089016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	141461511	+	chr8	141467765	+	.	8	0	4106315_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4106315_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:141461511(+)-8:141467765(-)__8_141463001_141488001D;SPAN=6254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=A[chr8:141467765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	141521746	+	chr8	141524467	+	.	0	16	4106502_1	23.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4106502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_141512001_141537001_56C;SPAN=2721;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:108 GQ:23.6 PL:[23.6, 0.0, 238.1] SR:16 DR:0 LR:-23.56 LO:33.95);ALT=G[chr8:141524467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35270594	+	chr8	141735346	+	.	17	88	4107225_1	99.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=4107225_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_141732501_141757501_70C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:73 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:88 DR:17 LR:-267.4 LO:267.4);ALT=]chr20:35270594]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	142402218	+	chr8	142431484	+	.	12	0	4109370_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4109370_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:142402218(+)-8:142431484(-)__8_142418501_142443501D;SPAN=29266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=C[chr8:142431484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	142428118	+	chr8	142431487	+	.	15	3	4109392_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4109392_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_142418501_142443501_117C;SPAN=3369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:70 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:3 DR:15 LR:-30.55 LO:34.51);ALT=G[chr8:142431487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	143304652	+	chr8	143302979	+	.	17	0	4111934_1	22.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=4111934_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:143302979(-)-8:143304652(+)__8_143300501_143325501D;SPAN=1673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:125 GQ:22.4 PL:[22.4, 0.0, 279.8] SR:0 DR:17 LR:-22.25 LO:35.39);ALT=]chr8:143304652]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	143310611	+	chr8	143312472	-	.	9	0	4111992_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4111992_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:143310611(+)-8:143312472(+)__8_143300501_143325501D;SPAN=1861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:117 GQ:1.8 PL:[0.0, 1.8, 287.1] SR:0 DR:9 LR:1.989 LO:16.38);ALT=G]chr8:143312472];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr8	143564804	+	chr8	143563439	+	.	12	0	4112635_1	13.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=4112635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:143563439(-)-8:143564804(+)__8_143545501_143570501D;SPAN=1365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:98 GQ:13.1 PL:[13.1, 0.0, 224.3] SR:0 DR:12 LR:-13.06 LO:24.39);ALT=]chr8:143564804]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr8	144100003	+	chr8	144102299	+	.	57	18	4114262_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4114262_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_8_144084501_144109501_279C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:70 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:18 DR:57 LR:-208.0 LO:208.0);ALT=G[chr8:144102299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144100038	+	chr8	144102800	+	.	13	0	4114264_1	18.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4114264_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144100038(+)-8:144102800(-)__8_144084501_144109501D;SPAN=2762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=C[chr8:144102800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144356972	+	chr8	144358066	+	.	2	5	4114850_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4114850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144354001_144379001_250C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:5 DR:2 LR:-3.059 LO:13.4);ALT=G[chr8:144358066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144411643	+	chr8	144413393	+	.	2	15	4115808_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4115808_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144403001_144428001_220C;SPAN=1750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:107 GQ:23.9 PL:[23.9, 0.0, 235.1] SR:15 DR:2 LR:-23.83 LO:34.02);ALT=T[chr8:144413393[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144411688	+	chr8	144416932	+	.	10	0	4115809_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4115809_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144411688(+)-8:144416932(-)__8_144403001_144428001D;SPAN=5244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:0 DR:10 LR:-7.543 LO:19.68);ALT=C[chr8:144416932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144413511	+	chr8	144416908	+	.	24	10	4115815_1	58.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4115815_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144403001_144428001_239C;SPAN=3397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:103 GQ:58.1 PL:[58.1, 0.0, 190.1] SR:10 DR:24 LR:-57.92 LO:61.95);ALT=T[chr8:144416908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144634067	+	chr8	144636240	+	.	0	47	4116095_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=TGT;MAPQ=60;MATEID=4116095_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_8_144623501_144648501_212C;SPAN=2173;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:74 GQ:42.8 PL:[135.2, 0.0, 42.8] SR:47 DR:0 LR:-137.6 LO:137.6);ALT=T[chr8:144636240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144663501	+	chr8	144668899	+	.	3	52	4116199_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4116199_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144648001_144673001_338C;SPAN=5398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:145 GQ:99 PL:[142.4, 0.0, 208.4] SR:52 DR:3 LR:-142.3 LO:143.0);ALT=G[chr8:144668899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144672283	+	chr8	144679515	+	.	8	0	4115995_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4115995_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144672283(+)-8:144679515(-)__8_144672501_144697501D;SPAN=7232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=G[chr8:144679515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	98558028	+	chr8	144716231	+	.	12	0	6056270_1	28.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=6056270_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144716231(-)-15:98558028(+)__15_98539001_98564001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=]chr15:98558028]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr8	144716350	+	chr15	98558143	+	.	15	0	6056271_1	35.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=6056271_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144716350(+)-15:98558143(-)__15_98539001_98564001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:50 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.97 LO:37.08);ALT=T[chr15:98558143[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr8	144720433	-	chr8	144721457	+	.	9	0	4116236_1	24.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4116236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144720433(-)-8:144721457(-)__8_144721501_144746501D;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:21 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.02 LO:24.03);ALT=[chr8:144721457[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr8	144903899	+	chr8	144911446	+	.	16	0	4116830_1	31.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4116830_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144903899(+)-8:144911446(-)__8_144893001_144918001D;SPAN=7547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:81 GQ:31.1 PL:[31.1, 0.0, 163.1] SR:0 DR:16 LR:-30.87 LO:36.16);ALT=G[chr8:144911446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144904086	+	chr8	144906482	+	.	0	13	4116832_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=4116832_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_144893001_144918001_132C;SPAN=2396;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:86 GQ:19.7 PL:[19.7, 0.0, 188.0] SR:13 DR:0 LR:-19.61 LO:27.71);ALT=G[chr8:144906482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	144904134	+	chr8	144911447	+	.	30	0	4116833_1	77.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4116833_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:144904134(+)-8:144911447(-)__8_144893001_144918001D;SPAN=7313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:79 GQ:77.6 PL:[77.6, 0.0, 113.9] SR:0 DR:30 LR:-77.63 LO:78.01);ALT=A[chr8:144911447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145133802	+	chr8	145134844	+	.	0	10	4117480_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4117480_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_145113501_145138501_63C;SPAN=1042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:103 GQ:5.3 PL:[5.3, 0.0, 242.9] SR:10 DR:0 LR:-5.105 LO:19.26);ALT=G[chr8:145134844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145512987	+	chr8	145514954	+	.	0	8	4118541_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4118541_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_145505501_145530501_97C;SPAN=1967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:8 DR:0 LR:-6.631 LO:15.85);ALT=T[chr8:145514954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145515556	+	chr8	145532591	+	.	0	15	4118686_1	37.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4118686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_145530001_145555001_289C;SPAN=17035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:44 GQ:37.7 PL:[37.7, 0.0, 67.4] SR:15 DR:0 LR:-37.59 LO:38.11);ALT=G[chr8:145532591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145650481	+	chr8	145653869	+	.	13	0	4119064_1	29.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4119064_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145650481(+)-8:145653869(-)__8_145628001_145653001D;SPAN=3388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:50 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:0 DR:13 LR:-29.37 LO:31.17);ALT=A[chr8:145653869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145650481	+	chr8	145652315	+	.	13	0	4119063_1	15.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4119063_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145650481(+)-8:145652315(-)__8_145628001_145653001D;SPAN=1834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:100 GQ:15.8 PL:[15.8, 0.0, 227.0] SR:0 DR:13 LR:-15.82 LO:26.79);ALT=A[chr8:145652315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145651155	+	chr8	145652292	+	TTCTCCCTCTCCCGGGCGTTCTTGTACAACTTCACTTCCTCATACAGCTCCGGCTTGTTCCCAGGGG	0	84	4119068_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TAC;INSERTION=TTCTCCCTCTCCCGGGCGTTCTTGTACAACTTCACTTCCTCATACAGCTCCGGCTTGTTCCCAGGGG;MAPQ=60;MATEID=4119068_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_8_145628001_145653001_92C;SPAN=1137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:100 GQ:7.2 PL:[257.4, 7.2, 0.0] SR:84 DR:0 LR:-267.7 LO:267.7);ALT=C[chr8:145652292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145651208	+	chr8	145653869	+	.	52	0	4119069_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4119069_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145651208(+)-8:145653869(-)__8_145628001_145653001D;SPAN=2661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:29 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=C[chr8:145653869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145651505	+	chr8	145653868	+	.	11	0	4119072_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4119072_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145651505(+)-8:145653868(-)__8_145628001_145653001D;SPAN=2363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:34 GQ:27.2 PL:[27.2, 0.0, 53.6] SR:0 DR:11 LR:-27.1 LO:27.63);ALT=A[chr8:145653868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	145652603	+	chr8	145653869	+	.	9	0	4119077_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4119077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=8:145652603(+)-8:145653869(-)__8_145628001_145653001D;SPAN=1266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:27 GQ:22.4 PL:[22.4, 0.0, 42.2] SR:0 DR:9 LR:-22.39 LO:22.75);ALT=A[chr8:145653869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	146076781	+	chr8	146078223	+	.	11	4	4120238_1	9.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4120238_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_146069001_146094001_227C;SPAN=1442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:4 DR:11 LR:-9.219 LO:21.81);ALT=C[chr8:146078223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr8	146221997	+	chr8	146224989	+	.	2	2	4120804_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTAA;MAPQ=60;MATEID=4120804_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_8_146216001_146241001_197C;SPAN=2992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:2 DR:2 LR:13.62 LO:6.133);ALT=A[chr8:146224989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	4722627	+	chr9	4740937	+	.	18	25	4129213_1	89.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4129213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_4728501_4753501_130C;SPAN=18310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:29 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:25 DR:18 LR:-89.12 LO:89.12);ALT=T[chr9:4740937[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	5361890	+	chr9	5436567	+	GAAGTCGAGCATTCATAAGCATGAACTCCTTTTGATTTTTCATGCTTTCATTCATAGATTTTGAAAATATAAACCCCATTTTG	0	25	4130145_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=GAAGTCGAGCATTCATAAGCATGAACTCCTTTTGATTTTTCATGCTTTCATTCATAGATTTTGAAAATATAAACCCCATTTTG;MAPQ=60;MATEID=4130145_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_5414501_5439501_231C;SPAN=74677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:21 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:25 DR:0 LR:-72.62 LO:72.62);ALT=T[chr9:5436567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	5432036	+	chr9	5437785	+	.	14	0	4130169_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4130169_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:5432036(+)-9:5437785(-)__9_5414501_5439501D;SPAN=5749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:46 GQ:33.8 PL:[33.8, 0.0, 76.7] SR:0 DR:14 LR:-33.75 LO:34.71);ALT=T[chr9:5437785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	5436694	+	chr9	5437786	+	.	13	6	4130172_1	36.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAC;MAPQ=60;MATEID=4130172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_5414501_5439501_160C;SPAN=1092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:6 DR:13 LR:-36.83 LO:38.71);ALT=C[chr9:5437786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	6700570	+	chr9	6710599	+	.	18	0	4132150_1	52.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TTTCACCATGTTGGCTAGGCTGGTCTCAAACTCCTGATCTCAGGTGATCCACCTGCCTCGGCCTCCCAAAGTGCTAGGATTACAGGCATGAG;MAPQ=60;MATEID=4132150_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_9_6688501_6713501_51C;SPAN=10029;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:13 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=G[chr9:6710599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	6758166	+	chr9	6792967	+	.	8	0	4132472_1	19.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4132472_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:6758166(+)-9:6792967(-)__9_6737501_6762501D;SPAN=34801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:27 GQ:19.1 PL:[19.1, 0.0, 45.5] SR:0 DR:8 LR:-19.09 LO:19.72);ALT=T[chr9:6792967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	129647131	+	chr9	10208234	+	.	28	0	4717576_1	82.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4717576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:10208234(-)-10:129647131(+)__10_129629501_129654501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:20 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:0 DR:28 LR:-82.52 LO:82.52);ALT=]chr10:129647131]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	10798394	-	chr20	24867273	+	.	17	0	4137961_1	49.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4137961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:10798394(-)-20:24867273(-)__9_10780001_10805001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:15 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:17 LR:-49.51 LO:49.51);ALT=[chr20:24867273[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	15472750	+	chr9	15474007	+	.	3	6	4144049_1	13.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4144049_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_15459501_15484501_297C;SPAN=1257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:6 DR:3 LR:-13.13 LO:17.35);ALT=T[chr9:15474007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	32315161	+	chrX	55088075	-	.	4	32	7428697_1	95.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ATTCTTTTAGTTATTTTAAAATGTATGATTAAATTATT;MAPQ=60;MATEID=7428697_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_23_55076001_55101001_97C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:25 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:32 DR:4 LR:-95.72 LO:95.72);ALT=T]chrX:55088075];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	32571051	+	chr9	32572877	+	.	0	35	4170481_1	84.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=4170481_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_32560501_32585501_52C;SPAN=1826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:116 GQ:84.2 PL:[84.2, 0.0, 196.4] SR:35 DR:0 LR:-84.11 LO:86.62);ALT=C[chr9:32572877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33025382	+	chr9	33026472	+	.	0	16	4172138_1	30.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4172138_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33001501_33026501_302C;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:82 GQ:30.8 PL:[30.8, 0.0, 166.1] SR:16 DR:0 LR:-30.6 LO:36.07);ALT=G[chr9:33026472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33037117	+	chr9	33038680	+	.	2	5	4172407_1	0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TTACCTT;MAPQ=60;MATEID=4172407_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33026001_33051001_131C;SPAN=1563;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:119 GQ:12.3 PL:[0.0, 12.3, 313.5] SR:5 DR:2 LR:12.43 LO:9.786);ALT=A[chr9:33038680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33073804	+	chr9	33076581	+	.	17	3	4172328_1	42.0	.	DISC_MAPQ=16;EVDNC=ASDIS;MAPQ=60;MATEID=4172328_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33050501_33075501_200C;SPAN=2777;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:3 DR:17 LR:-42.84 LO:43.35);ALT=A[chr9:33076581[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33255308	+	chr9	33256799	+	GAACCTTTTTTACCAAGCCTTTCCTTTTCAATCTACTGTCTTTGAAATTTTCTGGCAGGAT	0	33	4173215_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GAACCTTTTTTACCAAGCCTTTCCTTTTCAATCTACTGTCTTTGAAATTTTCTGGCAGGAT;MAPQ=60;MATEID=4173215_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_33246501_33271501_55C;SPAN=1491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:134 GQ:72.8 PL:[72.8, 0.0, 251.0] SR:33 DR:0 LR:-72.63 LO:78.21);ALT=T[chr9:33256799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33259033	+	chr9	33261085	+	.	0	9	4173231_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4173231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33246501_33271501_307C;SPAN=2052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:9 DR:0 LR:-2.075 LO:16.94);ALT=T[chr9:33261085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33261168	+	chr9	33262699	+	.	4	8	4173238_1	9.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4173238_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33246501_33271501_201C;SPAN=1531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:8 DR:4 LR:-9.169 LO:19.98);ALT=C[chr9:33262699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33262828	+	chr9	33264221	+	.	0	10	4173244_1	3.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4173244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_33246501_33271501_281C;SPAN=1393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:110 GQ:3.2 PL:[3.2, 0.0, 263.9] SR:10 DR:0 LR:-3.208 LO:18.96);ALT=C[chr9:33264221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33265149	+	chr9	33270620	+	.	15	0	4173259_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4173259_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33265149(+)-9:33270620(-)__9_33246501_33271501D;SPAN=5471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:117 GQ:17.9 PL:[17.9, 0.0, 265.4] SR:0 DR:15 LR:-17.82 LO:30.81);ALT=G[chr9:33270620[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	33339520	+	chr15	100798971	+	.	9	0	4173710_1	13.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=4173710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33339520(+)-15:100798971(-)__9_33320001_33345001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:59 GQ:13.7 PL:[13.7, 0.0, 129.2] SR:0 DR:9 LR:-13.72 LO:19.22);ALT=A[chr15:100798971[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	33361658	-	chr9	33362714	+	.	9	0	4173590_1	2.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4173590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33361658(-)-9:33362714(-)__9_33344501_33369501D;SPAN=1056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:100 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.617 LO:17.02);ALT=[chr9:33362714[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	33613971	-	chr9	33796667	+	.	24	0	4174883_1	70.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4174883_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33613971(-)-9:33796667(-)__9_33614001_33639001D;SPAN=182696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:32 GQ:4.7 PL:[70.7, 0.0, 4.7] SR:0 DR:24 LR:-73.59 LO:73.59);ALT=[chr9:33796667[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	33624302	+	chr15	60656730	-	.	8	0	4174915_1	7.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4174915_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33624302(+)-15:60656730(+)__9_33614001_33639001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:0 DR:8 LR:-6.901 LO:15.9);ALT=C]chr15:60656730];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	33625276	+	chr15	60639832	-	.	10	0	4174918_1	14.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=4174918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:33625276(+)-15:60639832(+)__9_33614001_33639001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:0 DR:10 LR:-14.59 LO:21.18);ALT=T]chr15:60639832];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	34125278	+	chr9	34126352	+	.	3	5	4177081_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4177081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_34104001_34129001_43C;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:117 GQ:11.7 PL:[0.0, 11.7, 306.9] SR:5 DR:3 LR:11.89 LO:9.831);ALT=G[chr9:34126352[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34329650	+	chr9	34339018	+	.	8	0	4178022_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4178022_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:34329650(+)-9:34339018(-)__9_34324501_34349501D;SPAN=9368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=C[chr9:34339018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34416144	+	chr9	34417247	-	.	8	0	4178341_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4178341_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:34416144(+)-9:34417247(+)__9_34398001_34423001D;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:0 DR:8 LR:-3.109 LO:15.25);ALT=A]chr9:34417247];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	34616112	+	chr9	34617882	+	.	0	24	4179200_1	50.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4179200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_34594001_34619001_361C;SPAN=1770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:107 GQ:50.3 PL:[50.3, 0.0, 208.7] SR:24 DR:0 LR:-50.24 LO:55.75);ALT=T[chr9:34617882[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34616161	+	chr9	34620362	+	.	11	0	4179201_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4179201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:34616161(+)-9:34620362(-)__9_34594001_34619001D;SPAN=4201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:0 DR:11 LR:-22.49 LO:25.34);ALT=C[chr9:34620362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34618018	+	chr9	34620362	+	.	42	0	4179209_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4179209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:34618018(+)-9:34620362(-)__9_34594001_34619001D;SPAN=2344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:47 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:42 LR:-137.9 LO:137.9);ALT=C[chr9:34620362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	34618759	+	chr9	34620363	+	.	51	25	4179028_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=4179028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_34618501_34643501_268C;SPAN=1604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:115 GQ:99 PL:[163.7, 0.0, 114.2] SR:25 DR:51 LR:-164.0 LO:164.0);ALT=T[chr9:34620363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35065380	+	chr9	35066671	+	.	6	3	4180787_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4180787_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35059501_35084501_415C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:105 GQ:5.1 PL:[0.0, 5.1, 264.0] SR:3 DR:6 LR:5.34 LO:12.29);ALT=T[chr9:35066671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35068359	+	chr9	35072334	+	.	12	9	4180800_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4180800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35059501_35084501_331C;SPAN=3975;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:120 GQ:26.9 PL:[26.9, 0.0, 264.5] SR:9 DR:12 LR:-26.91 LO:38.3);ALT=A[chr9:35072334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35725727	+	chr9	35732069	+	.	51	5	4183288_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCTG;MAPQ=60;MATEID=4183288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35721001_35746001_51C;SPAN=6342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:97 GQ:79.4 PL:[155.3, 0.0, 79.4] SR:5 DR:51 LR:-156.6 LO:156.6);ALT=G[chr9:35732069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	35813784	+	chr9	35814894	+	.	58	20	4183550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=4183550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_35794501_35819501_373C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:133 GQ:99 PL:[191.9, 0.0, 129.2] SR:20 DR:58 LR:-192.3 LO:192.3);ALT=G[chr9:35814894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36037098	+	chr9	36058822	+	CATTGTGTTGTAATCATTCAAAGGATAACCAAATGTGCCGTGATGTATGTGAAC	0	7	4184570_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CATTGTGTTGTAATCATTCAAAGGATAACCAAATGTGCCGTGATGTATGTGAAC;MAPQ=60;MATEID=4184570_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_36039501_36064501_339C;SPAN=21724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:26 GQ:16.1 PL:[16.1, 0.0, 45.8] SR:7 DR:0 LR:-16.06 LO:16.91);ALT=G[chr9:36058822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136823	+	chr9	36162355	+	.	11	0	4185052_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4185052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136823(+)-9:36162355(-)__9_36162001_36187001D;SPAN=25532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:0 DR:11 LR:-23.85 LO:25.91);ALT=C[chr9:36162355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136840	+	chr9	36150864	+	.	15	0	4184926_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4184926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136840(+)-9:36150864(-)__9_36113001_36138001D;SPAN=14024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:40 GQ:38.6 PL:[38.6, 0.0, 58.4] SR:0 DR:15 LR:-38.68 LO:38.9);ALT=G[chr9:36150864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136870	+	chr9	36147778	+	.	31	0	4184927_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4184927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136870(+)-9:36147778(-)__9_36113001_36138001D;SPAN=10908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:36 GQ:6.3 PL:[99.0, 6.3, 0.0] SR:0 DR:31 LR:-99.82 LO:99.82);ALT=G[chr9:36147778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36136870	+	chr9	36148542	+	.	47	0	4184928_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4184928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:36136870(+)-9:36148542(-)__9_36113001_36138001D;SPAN=11672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:36 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:0 DR:47 LR:-138.6 LO:138.6);ALT=G[chr9:36148542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36148648	+	chr9	36150865	+	.	2	47	4184792_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACAGG;MAPQ=60;MATEID=4184792_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_36137501_36162501_405C;SPAN=2217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:131 GQ:99 PL:[123.2, 0.0, 192.5] SR:47 DR:2 LR:-123.0 LO:123.9);ALT=G[chr9:36150865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36150947	+	chr9	36162358	+	.	5	11	4185053_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4185053_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_36162001_36187001_16C;SPAN=11411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:47 GQ:36.8 PL:[36.8, 0.0, 76.4] SR:11 DR:5 LR:-36.78 LO:37.57);ALT=G[chr9:36162358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36191270	+	chr9	36198974	+	ATGCTGTTGATGGAGTAATGAATGGTGAATACTACC	4	33	4184955_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGCTGTTGATGGAGTAATGAATGGTGAATACTACC;MAPQ=60;MATEID=4184955_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_36186501_36211501_296C;SPAN=7704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:96 GQ:89.6 PL:[89.6, 0.0, 142.4] SR:33 DR:4 LR:-89.53 LO:90.21);ALT=G[chr9:36198974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	36362896	+	chr9	36364080	+	.	134	101	4185954_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GCCTCCCAAAGTGCT;MAPQ=0;MATEID=4185954_2;MATENM=1;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_9_36358001_36383001_217C;SECONDARY;SPAN=1184;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:222 DP:39 GQ:59.8 PL:[656.8, 59.8, 0.0] SR:101 DR:134 LR:-656.9 LO:656.9);ALT=T[chr9:36364080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37120674	+	chr9	37126308	+	.	26	0	4188847_1	49.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4188847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:37120674(+)-9:37126308(-)__9_37117501_37142501D;SPAN=5634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:136 GQ:49.1 PL:[49.1, 0.0, 280.1] SR:0 DR:26 LR:-48.98 LO:58.35);ALT=C[chr9:37126308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37422794	+	chr9	37425915	+	.	16	0	4189927_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4189927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:37422794(+)-9:37425915(-)__9_37411501_37436501D;SPAN=3121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:121 GQ:20.3 PL:[20.3, 0.0, 271.1] SR:0 DR:16 LR:-20.03 LO:33.1);ALT=C[chr9:37425915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37422830	+	chr9	37424842	+	.	86	43	4189930_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4189930_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37411501_37436501_296C;SPAN=2012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:109 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:43 DR:86 LR:-326.8 LO:326.8);ALT=A[chr9:37424842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37424973	+	chr9	37426534	+	GGCCAATCTCAAAGTCATCAGCACCATGTCTGTGGGCATCGACCACTTGGCTTTGGATGAAATCAAGAAGC	0	57	4189940_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GGCCAATCTCAAAGTCATCAGCACCATGTCTGTGGGCATCGACCACTTGGCTTTGGATGAAATCAAGAAGC;MAPQ=60;MATEID=4189940_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_37411501_37436501_74C;SPAN=1561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:112 GQ:99 PL:[158.0, 0.0, 111.8] SR:57 DR:0 LR:-158.2 LO:158.2);ALT=G[chr9:37426534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37426651	+	chr9	37428481	+	.	2	6	4189947_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4189947_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37411501_37436501_176C;SPAN=1830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:134 GQ:9.6 PL:[0.0, 9.6, 343.2] SR:6 DR:2 LR:9.896 LO:13.65);ALT=A[chr9:37428481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37428570	+	chr9	37429726	+	.	0	5	4189956_1	0	.	EVDNC=ASSMB;HOMSEQ=TAGG;MAPQ=60;MATEID=4189956_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37411501_37436501_345C;SPAN=1156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:120 GQ:15.9 PL:[0.0, 15.9, 323.4] SR:5 DR:0 LR:16.01 LO:7.734);ALT=G[chr9:37429726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37432135	+	chr9	37436657	+	.	3	14	4190372_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4190372_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37436001_37461001_354C;SPAN=4522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:69 GQ:37.4 PL:[37.4, 0.0, 129.8] SR:14 DR:3 LR:-37.42 LO:40.29);ALT=G[chr9:37436657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37588930	+	chr9	37592307	+	.	58	4	4190789_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4190789_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_37583001_37608001_124C;SPAN=3377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:106 GQ:83.6 PL:[172.7, 0.0, 83.6] SR:4 DR:58 LR:-174.3 LO:174.3);ALT=C[chr9:37592307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	37637304	+	chr11	66036196	-	.	49	0	4894603_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4894603_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:37637304(+)-11:66036196(+)__11_66027501_66052501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:44 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:0 DR:49 LR:-145.2 LO:145.2);ALT=G]chr11:66036196];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	57480279	+	chr9	37885689	+	AGAGAAGT	0	24	4869904_1	66.0	.	EVDNC=ASSMB;INSERTION=AGAGAAGT;MAPQ=60;MATEID=4869904_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_57477001_57502001_194C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:46 GQ:43.7 PL:[66.8, 0.0, 43.7] SR:24 DR:0 LR:-66.99 LO:66.99);ALT=]chr11:57480279]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	38243898	+	chr15	63770026	+	.	31	0	5969671_1	89.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5969671_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:38243898(+)-15:63770026(-)__15_63749001_63774001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:20 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=A[chr15:63770026[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	70578661	+	chr20	33674281	-	.	8	0	6989564_1	14.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6989564_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:70578661(+)-20:33674281(+)__20_33663001_33688001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:0 DR:8 LR:-14.49 LO:17.76);ALT=A]chr20:33674281];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	93564288	+	chr9	93606135	+	.	48	0	4329568_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4329568_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:93564288(+)-9:93606135(-)__9_93590001_93615001D;SPAN=41847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:55 GQ:11.4 PL:[155.1, 11.4, 0.0] SR:0 DR:48 LR:-155.5 LO:155.5);ALT=G[chr9:93606135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	93607877	+	chr9	93624488	+	.	3	3	4329644_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4329644_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_93590001_93615001_379C;SPAN=16611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:47 GQ:0.5 PL:[0.5, 0.0, 112.7] SR:3 DR:3 LR:-0.4706 LO:7.462);ALT=G[chr9:93624488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	94395817	+	chr9	94403299	+	.	51	46	4332069_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=A;MAPQ=60;MATEID=4332069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_94374001_94399001_58C;SPAN=7482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:45 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:46 DR:51 LR:-227.8 LO:227.8);ALT=A[chr9:94403299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95050564	+	chr9	95051583	+	.	0	4	4334243_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4334243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_95035501_95060501_284C;SPAN=1019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:89 GQ:10.8 PL:[0.0, 10.8, 237.6] SR:4 DR:0 LR:10.91 LO:6.32);ALT=T[chr9:95051583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95526452	-	chr9	95527467	+	.	8	0	4336033_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4336033_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:95526452(-)-9:95527467(-)__9_95525501_95550501D;SPAN=1015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:0 DR:8 LR:-11.51 LO:16.91);ALT=[chr9:95527467[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	95726687	+	chr9	95737562	+	.	13	0	4336499_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4336499_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:95726687(+)-9:95737562(-)__9_95721501_95746501D;SPAN=10875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:96 GQ:17 PL:[17.0, 0.0, 215.0] SR:0 DR:13 LR:-16.9 LO:27.04);ALT=T[chr9:95737562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95821113	+	chr9	95838063	+	.	5	5	4336671_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4336671_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_95819501_95844501_139C;SPAN=16950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:72 GQ:3.8 PL:[3.8, 0.0, 168.8] SR:5 DR:5 LR:-3.6 LO:13.48);ALT=G[chr9:95838063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95858634	+	chr9	95869954	+	.	63	21	4337099_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4337099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_95868501_95893501_16C;SPAN=11320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:58 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:21 DR:63 LR:-201.3 LO:201.3);ALT=G[chr9:95869954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95858677	+	chr9	95872847	+	.	28	0	4337101_1	73.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4337101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:95858677(+)-9:95872847(-)__9_95868501_95893501D;SPAN=14170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:69 GQ:73.7 PL:[73.7, 0.0, 93.5] SR:0 DR:28 LR:-73.73 LO:73.87);ALT=G[chr9:95872847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95870109	+	chr9	95872848	+	.	5	7	4337116_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4337116_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_95868501_95893501_37C;SPAN=2739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:116 GQ:5 PL:[5.0, 0.0, 275.6] SR:7 DR:5 LR:-4.884 LO:21.06);ALT=G[chr9:95872848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95873004	+	chr9	95874500	+	.	0	4	4337128_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4337128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_95868501_95893501_180C;SPAN=1496;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:91 GQ:11.1 PL:[0.0, 11.1, 240.9] SR:4 DR:0 LR:11.45 LO:6.281);ALT=G[chr9:95874500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95887345	+	chr9	95896425	+	AAGGAAGATGAGCAGCACCCCCACGCCGATCTGCAGCACAAGGGAGATGGAGATGAGGACCACCAGGGGCACATAGAAGGCGAAGCTGGGGCCCTGTTCCACGACGGCCTTCAGCTGGGACGCGTTGGCCATCAGCAGCGCGATGTCCAGCATGCTCTCGGCTGCGCTCTTCTTGCTGGCGTAATGGTTCACGTTGATGGGCCCGTGCCTCCAGCCCCAGCGGGCCGG	0	18	4337182_1	46.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AAGGAAGATGAGCAGCACCCCCACGCCGATCTGCAGCACAAGGGAGATGGAGATGAGGACCACCAGGGGCACATAGAAGGCGAAGCTGGGGCCCTGTTCCACGACGGCCTTCAGCTGGGACGCGTTGGCCATCAGCAGCGCGATGTCCAGCATGCTCTCGGCTGCGCTCTTCTTGCTGGCGTAATGGTTCACGTTGATGGGCCCGTGCCTCCAGCCCCAGCGGGCCGG;MAPQ=60;MATEID=4337182_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_9_95868501_95893501_130C;SPAN=9080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:48 GQ:46.4 PL:[46.4, 0.0, 69.5] SR:18 DR:0 LR:-46.41 LO:46.68);ALT=C[chr9:95896425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	95888921	+	chr9	95896425	+	.	44	9	4337300_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4337300_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_95893001_95918001_203C;SPAN=7504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:35 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:9 DR:44 LR:-145.2 LO:145.2);ALT=C[chr9:95896425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	99029763	-	chr9	99031131	+	.	8	0	4348163_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4348163_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:99029763(-)-9:99031131(-)__9_99029001_99054001D;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=[chr9:99031131[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	99413779	+	chr9	99417372	+	CAATATGATGGTAGGATGACTGTCCAATCACTATAAGGGTGACATTTGCTTCTTGTAAGAAACTCCTGGGGATTTTGGCCAGATCCTCTACGTATTCCTTGCAGATGTAACACAGGAAATG	0	23	4349865_1	54.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CAATATGATGGTAGGATGACTGTCCAATCACTATAAGGGTGACATTTGCTTCTTGTAAGAAACTCCTGGGGATTTTGGCCAGATCCTCTACGTATTCCTTGCAGATGTAACACAGGAAATG;MAPQ=60;MATEID=4349865_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_9_99396501_99421501_174C;SPAN=3593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:79 GQ:54.5 PL:[54.5, 0.0, 137.0] SR:23 DR:0 LR:-54.52 LO:56.49);ALT=T[chr9:99417372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100396200	+	chr9	100403075	+	.	4	4	4353459_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=4353459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_100376501_100401501_378C;SPAN=6875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:47 GQ:3.8 PL:[3.8, 0.0, 109.4] SR:4 DR:4 LR:-3.772 LO:9.838);ALT=G[chr9:100403075[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100456043	+	chr9	100459402	+	.	0	7	4353704_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4353704_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_100450001_100475001_234C;SPAN=3359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:109 GQ:6.3 PL:[0.0, 6.3, 277.2] SR:7 DR:0 LR:6.424 LO:12.17);ALT=T[chr9:100459402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100760967	+	chr9	100767252	+	.	11	0	4354699_1	11.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=4354699_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:100760967(+)-9:100767252(-)__9_100744001_100769001D;SPAN=6285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:0 DR:11 LR:-10.84 LO:22.13);ALT=A[chr9:100767252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100767244	-	chr15	75614477	+	.	15	0	5990983_1	41.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5990983_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:100767244(-)-15:75614477(-)__15_75607001_75632001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:30 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:0 DR:15 LR:-41.46 LO:41.46);ALT=[chr15:75614477[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	100767435	+	chr9	100773551	+	.	9	39	4354719_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4354719_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_100744001_100769001_245C;SPAN=6116;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:70 GQ:30.5 PL:[139.4, 0.0, 30.5] SR:39 DR:9 LR:-143.4 LO:143.4);ALT=G[chr9:100773551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100773672	+	chr9	100777644	+	TCATCCTCATCCTCATCTTCATCTTCTTCATCAAGTCCAAATTCTTCTT	17	63	4355119_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=TCATCCTCATCCTCATCTTCATCTTCTTCATCAAGTCCAAATTCTTCTT;MAPQ=60;MATEID=4355119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_100768501_100793501_123C;SPAN=3972;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:76 DP:120 GQ:73.1 PL:[218.3, 0.0, 73.1] SR:63 DR:17 LR:-222.4 LO:222.4);ALT=G[chr9:100777644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100774789	+	chr9	100777708	+	.	8	0	4355124_1	0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=4355124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:100774789(+)-9:100777708(-)__9_100768501_100793501D;SPAN=2919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:139 GQ:11.1 PL:[0.0, 11.1, 359.7] SR:0 DR:8 LR:11.25 LO:13.52);ALT=T[chr9:100777708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100799448	-	chr9	100800539	+	.	9	0	4354765_1	0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4354765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:100799448(-)-9:100800539(-)__9_100793001_100818001D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:109 GQ:0.2 PL:[0.2, 0.0, 264.2] SR:0 DR:9 LR:-0.1782 LO:16.67);ALT=[chr9:100800539[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	100819223	+	chr9	100823062	+	.	0	37	4354981_1	87.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4354981_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_9_100817501_100842501_30C;SPAN=3839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:129 GQ:87.2 PL:[87.2, 0.0, 225.8] SR:37 DR:0 LR:-87.19 LO:90.59);ALT=G[chr9:100823062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	100843364	+	chr9	100845126	+	.	0	26	4354876_1	54.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4354876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_100842001_100867001_318C;SPAN=1762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:115 GQ:54.8 PL:[54.8, 0.0, 223.1] SR:26 DR:0 LR:-54.67 LO:60.5);ALT=G[chr9:100845126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32575908	+	chr9	101475196	+	ACACACAGA	14	20	7270977_1	79.0	.	DISC_MAPQ=43;EVDNC=ASDIS;INSERTION=ACACACAGA;MAPQ=57;MATEID=7270977_2;MATENM=1;NM=7;NUMPARTS=2;SCTG=c_22_32560501_32585501_445C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:26 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:20 DR:14 LR:-79.22 LO:79.22);ALT=]chr22:32575908]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr9	101984648	+	chr9	101990179	+	CTGCCGGACAGTGGATCCCGCCGCCCGGGCGGCCACTGCTTTGCTGGGAGAGCGCCCTGAGGATCCCACGTTAGTGCCACTGGGGGTCGGACCAGG	62	146	4358926_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CTGCCGGACAGTGGATCCCGCCGCCCGGGCGGCCACTGCTTTGCTGGGAGAGCGCCCTGAGGATCCCACGTTAGTGCCACTGGGGGTCGGACCAGG;MAPQ=60;MATEID=4358926_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_101969001_101994001_136C;SPAN=5531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:185 DP:150 GQ:49.9 PL:[547.9, 49.9, 0.0] SR:146 DR:62 LR:-547.9 LO:547.9);ALT=G[chr9:101990179[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	102677644	+	chr9	102713340	+	TATCAAAGGTGCAGAATCTGGGACAAGTTGCATGAAGAGCATATCAATGCAGGACGTACAGTTC	0	8	4361003_1	14.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TATCAAAGGTGCAGAATCTGGGACAAGTTGCATGAAGAGCATATCAATGCAGGACGTACAGTTC;MAPQ=60;MATEID=4361003_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_102655001_102680001_181C;SPAN=35696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:8 DR:0 LR:-14.76 LO:17.85);ALT=G[chr9:102713340[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	102769973	+	chr9	102778603	+	.	2	4	4361380_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4361380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_102753001_102778001_99C;SPAN=8630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:45 GQ:7.7 PL:[7.7, 0.0, 100.1] SR:4 DR:2 LR:-7.614 LO:12.43);ALT=T[chr9:102778603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	102822481	+	chr9	102861199	+	.	10	0	4361426_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4361426_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:102822481(+)-9:102861199(-)__9_102851001_102876001D;SPAN=38718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:0 DR:10 LR:-14.86 LO:21.25);ALT=A[chr9:102861199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	103064587	+	chr9	103065914	+	.	0	5	4362174_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4362174_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_103047001_103072001_77C;SPAN=1327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:105 GQ:11.7 PL:[0.0, 11.7, 277.2] SR:5 DR:0 LR:11.94 LO:8.028);ALT=C[chr9:103065914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	105967270	+	chr17	74553940	-	.	99	0	6501910_1	99.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=6501910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:105967270(+)-17:74553940(+)__17_74529001_74554001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:39 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:0 DR:99 LR:-293.8 LO:293.8);ALT=C]chr17:74553940];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr9	106568322	+	chr9	106569729	+	.	45	0	4371896_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4371896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:106568322(+)-9:106569729(-)__9_106550501_106575501D;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:45 LR:-132.0 LO:132.0);ALT=A[chr9:106569729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	107362880	+	chr9	107369022	+	.	12	0	4374444_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4374444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:107362880(+)-9:107369022(-)__9_107359001_107384001D;SPAN=6142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:0 DR:12 LR:-23.36 LO:27.2);ALT=G[chr9:107369022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	107369441	+	chr9	107363217	+	.	14	9	4374448_1	59.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCTAATTTCTTGAAATAAGAAGAAAAATTCTTATTTCCTCCT;MAPQ=60;MATEID=4374448_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_9_107359001_107384001_306C;SPAN=6224;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:61 GQ:59.6 PL:[59.6, 0.0, 86.0] SR:9 DR:14 LR:-59.4 LO:59.71);ALT=]chr9:107369441]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	107369914	+	chr9	107363718	+	.	11	0	4374451_1	5.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=4374451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:107363718(-)-9:107369914(+)__9_107359001_107384001D;SPAN=6196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:113 GQ:5.9 PL:[5.9, 0.0, 266.6] SR:0 DR:11 LR:-5.697 LO:21.19);ALT=]chr9:107369914]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	107510133	+	chr9	107513233	+	.	46	18	4374800_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=4374800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_107506001_107531001_333C;SPAN=3100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:112 GQ:99 PL:[151.4, 0.0, 118.4] SR:18 DR:46 LR:-151.4 LO:151.4);ALT=G[chr9:107513233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	107513447	+	chr9	107515186	+	.	0	11	4374809_1	9.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4374809_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_107506001_107531001_156C;SPAN=1739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:98 GQ:9.8 PL:[9.8, 0.0, 227.6] SR:11 DR:0 LR:-9.76 LO:21.91);ALT=G[chr9:107515186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	108007185	+	chr9	108061499	+	.	0	9	4376734_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4376734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_107996001_108021001_326C;SPAN=54314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:9 DR:0 LR:-20.5 LO:21.66);ALT=G[chr9:108061499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	108457054	+	chr9	108467877	+	.	0	10	4378263_1	21.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4378263_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_108461501_108486501_87C;SPAN=10823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:10 DR:0 LR:-21.63 LO:23.53);ALT=G[chr9:108467877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	109879128	-	chr11	34937799	+	.	10	0	4820940_1	20.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=4820940_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:109879128(-)-11:34937799(-)__11_34937001_34962001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:0 DR:10 LR:-20.28 LO:22.97);ALT=[chr11:34937799[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr9	110018286	+	chr9	110020849	+	.	18	13	4382753_1	53.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=ATAAATCTT;MAPQ=60;MATEID=4382753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_110005001_110030001_54C;SPAN=2563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:143 GQ:53.9 PL:[53.9, 0.0, 291.5] SR:13 DR:18 LR:-53.69 LO:63.17);ALT=T[chr9:110020849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110033387	+	chr9	110035549	-	.	3	3	4382960_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;MAPQ=60;MATEID=4382960_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_110029501_110054501_184C;SPAN=2162;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:91 GQ:7.8 PL:[0.0, 7.8, 234.3] SR:3 DR:3 LR:8.149 LO:8.345);ALT=A]chr9:110035549];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr9	110033454	+	chr9	110035446	+	.	62	22	4382962_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=ATTATTATTATT;MAPQ=60;MATEID=4382962_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_110029501_110054501_364C;SPAN=1992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:66 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:22 DR:62 LR:-227.8 LO:227.8);ALT=T[chr9:110035446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110045978	+	chr9	110062421	+	.	2	3	4383001_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4383001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_110029501_110054501_353C;SPAN=16443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:32 GQ:8 PL:[8.0, 0.0, 67.4] SR:3 DR:2 LR:-7.835 LO:10.74);ALT=T[chr9:110062421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110248211	+	chr9	110249307	+	.	7	3	4383515_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTGT;MAPQ=60;MATEID=4383515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_110225501_110250501_12C;SPAN=1096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:96 GQ:7.1 PL:[7.1, 0.0, 224.9] SR:3 DR:7 LR:-7.001 LO:19.58);ALT=T[chr9:110249307[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	110537535	+	chr9	110540596	+	.	78	34	4384765_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TAAAAATATTTTGTA;MAPQ=60;MATEID=4384765_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_110519501_110544501_1C;SPAN=3061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:53 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:34 DR:78 LR:-283.9 LO:283.9);ALT=A[chr9:110540596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	114731359	-	chr9	114732663	+	.	10	0	4398580_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4398580_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:114731359(-)-9:114732663(-)__9_114709001_114734001D;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:120 GQ:0.5 PL:[0.5, 0.0, 290.9] SR:0 DR:10 LR:-0.4991 LO:18.56);ALT=[chr9:114732663[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	115017546	-	chr9	115018829	+	.	11	0	4399264_1	11.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=4399264_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:115017546(-)-9:115018829(-)__9_115003001_115028001D;SPAN=1283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:91 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:0 DR:11 LR:-11.66 LO:22.29);ALT=[chr9:115018829[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	115060197	+	chr9	115095750	+	.	0	11	4399915_1	21.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4399915_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_115052001_115077001_133C;SPAN=35553;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:11 DR:0 LR:-21.68 LO:25.03);ALT=C[chr9:115095750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	115142495	+	chr9	115166273	+	.	10	0	4400665_1	16.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4400665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:115142495(+)-9:115166273(-)__9_115125501_115150501D;SPAN=23778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:0 DR:10 LR:-16.21 LO:21.62);ALT=G[chr9:115166273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	115166438	+	chr9	115167904	+	.	0	7	4400451_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4400451_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_115150001_115175001_34C;SPAN=1466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:117 GQ:8.4 PL:[0.0, 8.4, 300.3] SR:7 DR:0 LR:8.591 LO:11.95);ALT=A[chr9:115167904[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	115973873	+	chr9	115983471	+	.	4	4	4403746_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4403746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_115958501_115983501_405C;SPAN=9598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:86 GQ:3.3 PL:[0.0, 3.3, 214.5] SR:4 DR:4 LR:3.494 LO:10.65);ALT=C[chr9:115983471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	115983959	+	chr9	115989556	+	.	4	3	4403578_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4403578_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_115983001_116008001_352C;SPAN=5597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:103 GQ:11.1 PL:[0.0, 11.1, 270.6] SR:3 DR:4 LR:11.4 LO:8.071);ALT=G[chr9:115989556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	116112060	+	chr9	116116519	+	.	0	7	4404089_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4404089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_116105501_116130501_202C;SPAN=4459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.547 LO:12.74);ALT=G[chr9:116116519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	116116618	+	chr9	116122786	+	.	3	3	4404106_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4404106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_116105501_116130501_92C;SPAN=6168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:105 GQ:11.7 PL:[0.0, 11.7, 277.2] SR:3 DR:3 LR:11.94 LO:8.028);ALT=G[chr9:116122786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	116155929	+	chr9	116163490	+	.	9	0	4404182_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4404182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:116155929(+)-9:116163490(-)__9_116154501_116179501D;SPAN=7561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:117 GQ:1.8 PL:[0.0, 1.8, 287.1] SR:0 DR:9 LR:1.989 LO:16.38);ALT=G[chr9:116163490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	117099592	+	chr9	117103814	+	.	8	0	4407623_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4407623_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:117099592(+)-9:117103814(-)__9_117085501_117110501D;SPAN=4222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:112 GQ:3.6 PL:[0.0, 3.6, 277.2] SR:0 DR:8 LR:3.936 LO:14.29);ALT=G[chr9:117103814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	117143768	+	chr9	117150201	+	.	11	0	4407972_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4407972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:117143768(+)-9:117150201(-)__9_117134501_117159501D;SPAN=6433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:0 DR:11 LR:-11.39 LO:22.24);ALT=A[chr9:117150201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	117350201	+	chr9	117354832	+	.	87	52	4408633_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4408633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_117330501_117355501_306C;SPAN=4631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:119 DP:185 GQ:99 PL:[342.8, 0.0, 105.2] SR:52 DR:87 LR:-349.6 LO:349.6);ALT=G[chr9:117354832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123637035	+	chr9	123639369	+	.	0	10	4428122_1	9.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4428122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_123627001_123652001_287C;SPAN=2334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:10 DR:0 LR:-9.169 LO:19.98);ALT=C[chr9:123639369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123837325	+	chr9	123850572	+	.	11	0	4428946_1	21.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4428946_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:123837325(+)-9:123850572(-)__9_123847501_123872501D;SPAN=13247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:0 DR:11 LR:-21.68 LO:25.03);ALT=G[chr9:123850572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123837336	+	chr9	123842582	+	.	11	0	4428530_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4428530_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:123837336(+)-9:123842582(-)__9_123823001_123848001D;SPAN=5246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:115 GQ:5.3 PL:[5.3, 0.0, 272.6] SR:0 DR:11 LR:-5.155 LO:21.11);ALT=C[chr9:123842582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123943851	+	chr9	123945588	+	GTTTTTGCACTCGCTTCGAGGAACAATAAG	8	8	4428792_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTTTTTGCACTCGCTTCGAGGAACAATAAG;MAPQ=60;MATEID=4428792_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_123945501_123970501_96C;SPAN=1737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:45 GQ:34.1 PL:[34.1, 0.0, 73.7] SR:8 DR:8 LR:-34.02 LO:34.88);ALT=C[chr9:123945588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123954503	+	chr9	123963917	+	AATAATAATATATTTAAAGATGTAAGAGTAGTTGTATGGTGCAGTTGCCATGGTGGCA	0	35	4428816_1	89.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AATAATAATATATTTAAAGATGTAAGAGTAGTTGTATGGTGCAGTTGCCATGGTGGCA;MAPQ=60;MATEID=4428816_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_123945501_123970501_207C;SPAN=9414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:95 GQ:89.9 PL:[89.9, 0.0, 139.4] SR:35 DR:0 LR:-89.8 LO:90.41);ALT=C[chr9:123963917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	123955743	+	chr9	123964034	+	.	14	0	4428820_1	19.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4428820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:123955743(+)-9:123964034(-)__9_123945501_123970501D;SPAN=8291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:98 GQ:19.7 PL:[19.7, 0.0, 217.7] SR:0 DR:14 LR:-19.66 LO:29.47);ALT=A[chr9:123964034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124030552	+	chr9	124043744	+	.	19	0	4429175_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4429175_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:124030552(+)-9:124043744(-)__9_124043501_124068501D;SPAN=13192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:80 GQ:41 PL:[41.0, 0.0, 153.2] SR:0 DR:19 LR:-41.05 LO:44.68);ALT=G[chr9:124043744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124030552	+	chr9	124064234	+	.	84	0	4429176_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4429176_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:124030552(+)-9:124064234(-)__9_124043501_124068501D;SPAN=33682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:67 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=G[chr9:124064234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124043840	+	chr9	124064239	+	.	33	47	4429179_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4429179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_124043501_124068501_195C;SPAN=20399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:132 GQ:99 PL:[202.1, 0.0, 116.3] SR:47 DR:33 LR:-203.1 LO:203.1);ALT=G[chr9:124064239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124062283	+	chr9	124064240	+	.	14	6	4429246_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4429246_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_124043501_124068501_237C;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:129 GQ:27.8 PL:[27.8, 0.0, 285.2] SR:6 DR:14 LR:-27.77 LO:40.26);ALT=G[chr9:124064240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124081158	+	chr9	124083543	+	.	7	6	4429487_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4429487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_124068001_124093001_52C;SPAN=2385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:119 GQ:2.4 PL:[0.0, 2.4, 293.7] SR:6 DR:7 LR:2.531 LO:16.31);ALT=G[chr9:124083543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124083680	+	chr9	124086831	+	.	3	5	4429499_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4429499_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_9_124068001_124093001_186C;SPAN=3151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:125 GQ:13.8 PL:[0.0, 13.8, 330.0] SR:5 DR:3 LR:14.06 LO:9.655);ALT=G[chr9:124086831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124083680	+	chr9	124088786	+	CAGGGTGCCCAGTCTACCCAGGATGAGGTCGCTGCATCTGCCATCCTGACTGCTCAGCTGGATGAGGAGCTGGGAGGTACCCCTGT	8	11	4429500_1	24.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCAG;INSERTION=CAGGGTGCCCAGTCTACCCAGGATGAGGTCGCTGCATCTGCCATCCTGACTGCTCAGCTGGATGAGGAGCTGGGAGGTACCCCTGT;MAPQ=60;MATEID=4429500_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_124068001_124093001_186C;SPAN=5106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:117 GQ:24.5 PL:[24.5, 0.0, 258.8] SR:11 DR:8 LR:-24.42 LO:35.92);ALT=G[chr9:124088786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124086922	+	chr9	124088786	+	.	2	5	4429510_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCAG;MAPQ=60;MATEID=4429510_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_124068001_124093001_186C;SPAN=1864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:123 GQ:9.9 PL:[0.0, 9.9, 316.8] SR:5 DR:2 LR:10.22 LO:11.79);ALT=G[chr9:124088786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124089760	+	chr9	124091166	+	.	9	8	4429520_1	19.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4429520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_124068001_124093001_257C;SPAN=1406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:110 GQ:19.7 PL:[19.7, 0.0, 247.4] SR:8 DR:9 LR:-19.71 LO:31.24);ALT=G[chr9:124091166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124091628	+	chr9	124094710	+	.	10	0	4429346_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4429346_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:124091628(+)-9:124094710(-)__9_124092501_124117501D;SPAN=3082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:0 DR:10 LR:-14.59 LO:21.18);ALT=G[chr9:124094710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124118457	+	chr9	124132445	+	.	9	0	4429267_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4429267_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:124118457(+)-9:124132445(-)__9_124117001_124142001D;SPAN=13988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:119 GQ:2.4 PL:[0.0, 2.4, 293.7] SR:0 DR:9 LR:2.531 LO:16.31);ALT=A[chr9:124132445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	124914689	+	chr9	124921902	+	.	0	7	4432215_1	0	.	EVDNC=ASSMB;HOMSEQ=TCACCT;MAPQ=60;MATEID=4432215_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_124901001_124926001_81C;SPAN=7213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:108 GQ:6 PL:[0.0, 6.0, 273.9] SR:7 DR:0 LR:6.153 LO:12.2);ALT=T[chr9:124921902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	125023789	+	chr9	125026994	+	.	11	5	4432528_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4432528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_125023501_125048501_26C;SPAN=3205;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:105 GQ:17.9 PL:[17.9, 0.0, 235.7] SR:5 DR:11 LR:-17.77 LO:29.01);ALT=T[chr9:125026994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	125589074	+	chr9	125590750	+	.	6	3	4434058_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4434058_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_125587001_125612001_88C;SPAN=1676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:118 GQ:2.1 PL:[0.0, 2.1, 290.4] SR:3 DR:6 LR:2.26 LO:16.34);ALT=G[chr9:125590750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	125659857	+	chr9	125667389	+	.	5	10	4434578_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4434578_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_125660501_125685501_407C;SPAN=7532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:10 DR:5 LR:-29.05 LO:29.82);ALT=T[chr9:125667389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	126554965	+	chr9	126692166	+	.	9	0	4438061_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4438061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:126554965(+)-9:126692166(-)__9_126689501_126714501D;SPAN=137201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=G[chr9:126692166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	126641300	+	chr9	126692167	+	.	5	4	4438062_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4438062_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_9_126689501_126714501_13C;SPAN=50867;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:40 GQ:8.9 PL:[8.9, 0.0, 88.1] SR:4 DR:5 LR:-8.969 LO:12.77);ALT=C[chr9:126692167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127020370	+	chr9	127074783	+	.	11	0	4439355_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4439355_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127020370(+)-9:127074783(-)__9_127057001_127082001D;SPAN=54413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:0 DR:11 LR:-21.68 LO:25.03);ALT=T[chr9:127074783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127020381	+	chr9	127064213	+	.	22	0	4439356_1	57.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4439356_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127020381(+)-9:127064213(-)__9_127057001_127082001D;SPAN=43832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:55 GQ:57.8 PL:[57.8, 0.0, 74.3] SR:0 DR:22 LR:-57.72 LO:57.86);ALT=T[chr9:127064213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127064333	+	chr9	127074785	+	.	2	23	4439373_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4439373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127057001_127082001_122C;SPAN=10452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:105 GQ:50.9 PL:[50.9, 0.0, 202.7] SR:23 DR:2 LR:-50.78 LO:55.98);ALT=G[chr9:127074785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127115990	+	chr9	127119042	+	.	5	60	4439594_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4439594_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127106001_127131001_300C;SPAN=3052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:122 GQ:99 PL:[178.4, 0.0, 115.7] SR:60 DR:5 LR:-178.9 LO:178.9);ALT=T[chr9:127119042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127119196	+	chr9	127167594	+	CCATGTCTGGCCTAAACTTATCTTCAAATACAGCCATTGCTGCCAAGGAGCCAGA	3	16	4439650_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=CCATGTCTGGCCTAAACTTATCTTCAAATACAGCCATTGCTGCCAAGGAGCCAGA;MAPQ=60;MATEID=4439650_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_127155001_127180001_246C;SPAN=48398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:46 GQ:47 PL:[47.0, 0.0, 63.5] SR:16 DR:3 LR:-46.96 LO:47.11);ALT=T[chr9:127167594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127167714	+	chr9	127174628	+	.	5	6	4439692_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCTG;MAPQ=60;MATEID=4439692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127155001_127180001_87C;SPAN=6914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:6 DR:5 LR:-1.533 LO:16.86);ALT=G[chr9:127174628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127174771	+	chr9	127176187	+	.	0	39	4439711_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4439711_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127155001_127180001_140C;SPAN=1416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:109 GQ:99 PL:[99.2, 0.0, 165.2] SR:39 DR:0 LR:-99.21 LO:100.1);ALT=A[chr9:127176187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127174819	+	chr9	127177650	+	.	20	0	4439712_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4439712_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127174819(+)-9:127177650(-)__9_127155001_127180001D;SPAN=2831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:103 GQ:38.3 PL:[38.3, 0.0, 209.9] SR:0 DR:20 LR:-38.12 LO:45.04);ALT=C[chr9:127177650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127176335	+	chr9	127177645	+	.	55	0	4439715_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4439715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127176335(+)-9:127177645(-)__9_127155001_127180001D;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:112 GQ:99 PL:[151.4, 0.0, 118.4] SR:0 DR:55 LR:-151.4 LO:151.4);ALT=A[chr9:127177645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127631719	+	chr9	127635971	+	.	0	36	4441266_1	83.0	.	EVDNC=ASSMB;HOMSEQ=A;MAPQ=60;MATEID=4441266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127620501_127645501_368C;SPAN=4252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:132 GQ:83.3 PL:[83.3, 0.0, 235.1] SR:36 DR:0 LR:-83.07 LO:87.2);ALT=A[chr9:127635971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127636044	+	chr9	127637252	+	.	0	14	4441277_1	16.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4441277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127620501_127645501_318C;SPAN=1208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:111 GQ:16.4 PL:[16.4, 0.0, 250.7] SR:14 DR:0 LR:-16.14 LO:28.65);ALT=G[chr9:127637252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127818331	+	chr9	127905694	+	.	8	0	4442432_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4442432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127818331(+)-9:127905694(-)__9_127890001_127915001D;SPAN=87363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=A[chr9:127905694[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127920662	+	chr9	127923119	+	.	0	11	4442583_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4442583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127914501_127939501_182C;SPAN=2457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:93 GQ:11.3 PL:[11.3, 0.0, 212.6] SR:11 DR:0 LR:-11.12 LO:22.18);ALT=C[chr9:127923119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127923187	+	chr9	127933364	+	.	0	21	4442599_1	40.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4442599_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127914501_127939501_301C;SPAN=10177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:106 GQ:40.7 PL:[40.7, 0.0, 215.6] SR:21 DR:0 LR:-40.6 LO:47.5);ALT=T[chr9:127933364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127923230	+	chr9	127951925	+	.	11	0	4442687_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4442687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127923230(+)-9:127951925(-)__9_127939001_127964001D;SPAN=28695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:60 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-20.06 LO:24.46);ALT=G[chr9:127951925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127933461	+	chr9	127951923	+	.	33	22	4442688_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4442688_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127939001_127964001_116C;SPAN=18462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:59 GQ:23.6 PL:[119.3, 0.0, 23.6] SR:22 DR:33 LR:-123.0 LO:123.0);ALT=T[chr9:127951923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127962904	+	chr9	127965284	+	.	11	0	4442786_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4442786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:127962904(+)-9:127965284(-)__9_127939001_127964001D;SPAN=2380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:0 DR:11 LR:-20.87 LO:24.74);ALT=C[chr9:127965284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127963186	+	chr9	127965285	+	.	6	11	4442788_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4442788_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127939001_127964001_176C;SPAN=2099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:11 DR:6 LR:-36.83 LO:38.71);ALT=G[chr9:127965285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	127965347	+	chr9	127969842	+	.	0	11	4442949_1	9.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=4442949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_127963501_127988501_212C;SPAN=4495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:11 DR:0 LR:-9.219 LO:21.81);ALT=T[chr9:127969842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	128024238	+	chr9	128061168	+	.	7	3	4443648_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4443648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_128012501_128037501_51C;SPAN=36930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:3 DR:7 LR:-15.84 LO:18.23);ALT=G[chr9:128061168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	128024239	+	chr9	128057736	+	.	4	2	4443649_1	6.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4443649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_128012501_128037501_387C;SPAN=33497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:38 GQ:6.2 PL:[6.2, 0.0, 85.4] SR:2 DR:4 LR:-6.21 LO:10.33);ALT=G[chr9:128057736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	129089291	+	chr9	129102786	+	.	9	0	4446619_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4446619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:129089291(+)-9:129102786(-)__9_129090501_129115501D;SPAN=13495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:47 GQ:17 PL:[17.0, 0.0, 96.2] SR:0 DR:9 LR:-16.98 LO:20.21);ALT=T[chr9:129102786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	129567408	+	chr9	129594762	+	.	13	0	4448627_1	25.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4448627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:129567408(+)-9:129594762(-)__9_129580501_129605501D;SPAN=27354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:64 GQ:25.7 PL:[25.7, 0.0, 128.0] SR:0 DR:13 LR:-25.57 LO:29.56);ALT=G[chr9:129594762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130565342	+	chr9	130566560	+	.	0	18	4452300_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CCAGG;MAPQ=60;MATEID=4452300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_130560501_130585501_19C;SPAN=1218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:129 GQ:24.5 PL:[24.5, 0.0, 288.5] SR:18 DR:0 LR:-24.47 LO:37.69);ALT=G[chr9:130566560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130677121	+	chr9	130678686	+	.	0	11	4452157_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4452157_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_130658501_130683501_109C;SPAN=1565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:88 GQ:12.5 PL:[12.5, 0.0, 200.6] SR:11 DR:0 LR:-12.47 LO:22.46);ALT=C[chr9:130678686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130677169	+	chr9	130679218	+	.	9	0	4452158_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4452158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:130677169(+)-9:130679218(-)__9_130658501_130683501D;SPAN=2049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:101 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:0 DR:9 LR:-2.346 LO:16.98);ALT=A[chr9:130679218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130698103	+	chr9	130699712	+	.	17	0	4452429_1	28.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4452429_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:130698103(+)-9:130699712(-)__9_130683001_130708001D;SPAN=1609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:104 GQ:28.1 PL:[28.1, 0.0, 222.8] SR:0 DR:17 LR:-27.94 LO:36.87);ALT=G[chr9:130699712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130698104	+	chr9	130700095	+	.	14	0	4452430_1	17.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4452430_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:130698104(+)-9:130700095(-)__9_130683001_130708001D;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:108 GQ:17 PL:[17.0, 0.0, 244.7] SR:0 DR:14 LR:-16.95 LO:28.83);ALT=G[chr9:130700095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130887725	+	chr9	130889718	+	.	0	7	4453167_1	0	.	EVDNC=ASSMB;HOMSEQ=CTGCG;MAPQ=60;MATEID=4453167_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_130879001_130904001_267C;SPAN=1993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:7 DR:0 LR:1.005 LO:12.81);ALT=G[chr9:130889718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	130922765	+	chr9	130925719	+	.	137	104	4453309_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4453309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_130903501_130928501_315C;SPAN=2954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:198 DP:184 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:104 DR:137 LR:-587.5 LO:587.5);ALT=G[chr9:130925719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131038678	+	chr9	131046788	+	.	16	0	4453857_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4453857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131038678(+)-9:131046788(-)__9_131026001_131051001D;SPAN=8110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:111 GQ:23 PL:[23.0, 0.0, 244.1] SR:0 DR:16 LR:-22.74 LO:33.74);ALT=G[chr9:131046788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131038682	+	chr9	131048218	+	ACTGAACCAAGACTTACCCGAAGTTGCCGCGGGGCCTTCCGATCCCCTAGGCCATTGCCCAAGTCTGGCCAGGCTGATGGGACCAGCGAGGAGTCTCTGCACCTTGACATTCAGAAACTGAAGGAGAAGAGGGACATGCTGGACAAGGAGATCTCCCAGTTCGTATCTGA	4	21	4453859_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ACTGAACCAAGACTTACCCGAAGTTGCCGCGGGGCCTTCCGATCCCCTAGGCCATTGCCCAAGTCTGGCCAGGCTGATGGGACCAGCGAGGAGTCTCTGCACCTTGACATTCAGAAACTGAAGGAGAAGAGGGACATGCTGGACAAGGAGATCTCCCAGTTCGTATCTGA;MAPQ=60;MATEID=4453859_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_9_131026001_131051001_24C;SPAN=9536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:113 GQ:38.9 PL:[38.9, 0.0, 233.6] SR:21 DR:4 LR:-38.71 LO:46.84);ALT=G[chr9:131048218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131079506	+	chr9	131083878	+	.	0	10	4453929_1	8.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4453929_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131075001_131100001_126C;SPAN=4372;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:92 GQ:8.3 PL:[8.3, 0.0, 212.9] SR:10 DR:0 LR:-8.085 LO:19.77);ALT=C[chr9:131083878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131085207	+	chr9	131088056	+	.	11	0	4453968_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4453968_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131085207(+)-9:131088056(-)__9_131075001_131100001D;SPAN=2849;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:117 GQ:4.7 PL:[4.7, 0.0, 278.6] SR:0 DR:11 LR:-4.613 LO:21.02);ALT=G[chr9:131088056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131085215	+	chr9	131087419	+	.	32	0	4453969_1	71.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4453969_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131085215(+)-9:131087419(-)__9_131075001_131100001D;SPAN=2204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:128 GQ:71 PL:[71.0, 0.0, 239.3] SR:0 DR:32 LR:-70.95 LO:76.08);ALT=G[chr9:131087419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131085426	+	chr9	131087421	+	.	0	35	4453972_1	80.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4453972_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_131075001_131100001_118C;SPAN=1995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:132 GQ:80 PL:[80.0, 0.0, 238.4] SR:35 DR:0 LR:-79.77 LO:84.27);ALT=G[chr9:131087421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131133734	+	chr9	131140313	+	.	13	0	4454409_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4454409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131133734(+)-9:131140313(-)__9_131124001_131149001D;SPAN=6579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:104 GQ:14.9 PL:[14.9, 0.0, 236.0] SR:0 DR:13 LR:-14.74 LO:26.55);ALT=G[chr9:131140313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131133737	+	chr9	131151539	+	.	24	0	4454411_1	63.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4454411_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131133737(+)-9:131151539(-)__9_131124001_131149001D;SPAN=17802;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:58 GQ:63.5 PL:[63.5, 0.0, 76.7] SR:0 DR:24 LR:-63.51 LO:63.59);ALT=G[chr9:131151539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131133738	+	chr9	131150094	+	.	27	0	4454412_1	73.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4454412_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131133738(+)-9:131150094(-)__9_131124001_131149001D;SPAN=16356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:58 GQ:66.8 PL:[73.4, 0.0, 66.8] SR:0 DR:27 LR:-73.43 LO:73.43);ALT=T[chr9:131150094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131140386	+	chr9	131150095	+	.	0	12	4454450_1	26.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4454450_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131124001_131149001_114C;SPAN=9709;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:48 GQ:26.6 PL:[26.6, 0.0, 89.3] SR:12 DR:0 LR:-26.61 LO:28.53);ALT=G[chr9:131150095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131183356	+	chr9	131185146	+	.	0	7	4454532_1	0	.	EVDNC=ASSMB;HOMSEQ=GGTG;MAPQ=60;MATEID=4454532_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131173001_131198001_406C;SPAN=1790;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:97 GQ:3 PL:[0.0, 3.0, 240.9] SR:7 DR:0 LR:3.173 LO:12.54);ALT=G[chr9:131185146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131218517	+	chr9	131222790	+	.	10	0	4455070_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4455070_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131218517(+)-9:131222790(-)__9_131222001_131247001D;SPAN=4273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:0 DR:10 LR:-17.3 LO:21.94);ALT=G[chr9:131222790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131218536	+	chr9	131221845	+	.	12	8	4455071_1	46.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4455071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131222001_131247001_264C;SPAN=3309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:0 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:8 DR:12 LR:-46.21 LO:46.21);ALT=T[chr9:131221845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131267184	+	chr9	131271153	+	.	0	7	4454934_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4454934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131271001_131296001_10C;SPAN=3969;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:48 GQ:10.1 PL:[10.1, 0.0, 105.8] SR:7 DR:0 LR:-10.1 LO:14.8);ALT=G[chr9:131271153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131403219	+	chr9	131418829	+	GTCTCCCC	32	6	4455770_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTCTCCCC;MAPQ=60;MATEID=4455770_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_131418001_131443001_242C;SPAN=15610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:39 GQ:7.2 PL:[108.9, 7.2, 0.0] SR:6 DR:32 LR:-110.1 LO:110.1);ALT=C[chr9:131418829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131412068	+	chr9	131413977	+	.	77	92	4455535_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AGGTCAGGAGTT;MAPQ=60;MATEID=4455535_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_131393501_131418501_219C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:147 DP:26 GQ:39.7 PL:[435.7, 39.7, 0.0] SR:92 DR:77 LR:-435.7 LO:435.7);ALT=T[chr9:131413977[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131425701	+	chr9	131446679	+	.	9	0	4455812_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4455812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:131425701(+)-9:131446679(-)__9_131418001_131443001D;SPAN=20978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=G[chr9:131446679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131484854	+	chr9	131486273	+	.	0	9	4455633_1	1.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4455633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131467001_131492001_169C;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:106 GQ:1.1 PL:[1.1, 0.0, 255.2] SR:9 DR:0 LR:-0.991 LO:16.78);ALT=C[chr9:131486273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131589471	+	chr9	131591013	+	.	0	8	4456470_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4456470_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131589501_131614501_113C;SPAN=1542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:8 DR:0 LR:-3.379 LO:15.29);ALT=C[chr9:131591013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	131873910	+	chr9	131882790	+	.	8	10	4457763_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4457763_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_131859001_131884001_50C;SPAN=8880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:114 GQ:22.1 PL:[22.1, 0.0, 253.1] SR:10 DR:8 LR:-21.93 LO:33.54);ALT=G[chr9:131882790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132026700	+	chr9	132028070	+	.	112	66	4458261_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCTGGGATTACAGGT;MAPQ=60;MATEID=4458261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132006001_132031001_79C;SPAN=1370;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:148 DP:42 GQ:40 PL:[439.0, 40.0, 0.0] SR:66 DR:112 LR:-439.0 LO:439.0);ALT=T[chr9:132028070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132388575	+	chr9	132396333	+	.	7	3	4459727_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4459727_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132373501_132398501_219C;SPAN=7758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:3 DR:7 LR:2.36 LO:12.64);ALT=G[chr9:132396333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132388575	+	chr9	132394929	+	.	12	4	4459726_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4459726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132373501_132398501_373C;SPAN=6354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:101 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:4 DR:12 LR:-18.85 LO:29.27);ALT=G[chr9:132394929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132585126	+	chr9	132586187	+	.	0	15	4460413_1	22.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4460413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132569501_132594501_53C;SPAN=1061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:101 GQ:22.4 PL:[22.4, 0.0, 220.4] SR:15 DR:0 LR:-22.15 LO:31.85);ALT=C[chr9:132586187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132591820	+	chr9	132593150	+	.	0	6	4460443_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4460443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132569501_132594501_385C;SPAN=1330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:102 GQ:7.5 PL:[0.0, 7.5, 260.7] SR:6 DR:0 LR:7.828 LO:10.2);ALT=A[chr9:132593150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132594252	+	chr9	132597418	+	TTATCTTTGCCCCTTTCCTTCAGTTTCTTCATATCCACCATACCACCTGTCTTCATCTGAAAGGGATCATCCACTAGAGTGGTCTCCTCTTGTACCTTCTCTCCCACCAGCAAGGCCACAGCACTCACCCCGTTGGGCCTCTTCCTCAAGTTCTGTACCTCTCTGGTCTCTTCCAGTTTTAAT	3	39	4460572_1	99.0	.	DISC_MAPQ=48;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TTATCTTTGCCCCTTTCCTTCAGTTTCTTCATATCCACCATACCACCTGTCTTCATCTGAAAGGGATCATCCACTAGAGTGGTCTCCTCTTGTACCTTCTCTCCCACCAGCAAGGCCACAGCACTCACCCCGTTGGGCCTCTTCCTCAAGTTCTGTACCTCTCTGGTCTCTTCCAGTTTTAAT;MAPQ=60;MATEID=4460572_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_9_132594001_132619001_389C;SPAN=3166;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:112 GQ:99 PL:[101.9, 0.0, 167.9] SR:39 DR:3 LR:-101.7 LO:102.6);ALT=C[chr9:132597418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132596040	+	chr9	132597461	+	.	16	0	4460590_1	26.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=4460590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:132596040(+)-9:132597461(-)__9_132594001_132619001D;SPAN=1421;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:97 GQ:26.6 PL:[26.6, 0.0, 208.1] SR:0 DR:16 LR:-26.54 LO:34.77);ALT=T[chr9:132597461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132658277	+	chr9	132662242	+	.	3	5	4460859_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4460859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132643001_132668001_212C;SPAN=3965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:114 GQ:7.5 PL:[0.0, 7.5, 290.4] SR:5 DR:3 LR:7.778 LO:12.03);ALT=T[chr9:132662242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132662828	+	chr9	132665147	+	.	2	4	4460876_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4460876_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_132643001_132668001_399C;SPAN=2319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:100 GQ:13.8 PL:[0.0, 13.8, 270.6] SR:4 DR:2 LR:13.89 LO:6.115);ALT=T[chr9:132665147[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132665282	+	chr9	132671169	+	.	3	2	4460903_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4460903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132667501_132692501_8C;SPAN=5887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:51 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:2 DR:3 LR:0.6132 LO:7.314);ALT=T[chr9:132671169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132740891	+	chr9	132757121	+	TTGTATTCTTCTTCCTCCTTCGAGTTCTTTTTAGGTTGGTACTTCTTTGAAAGATT	0	10	4461382_1	24.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTGA;INSERTION=TTGTATTCTTCTTCCTCCTTCGAGTTCTTTTTAGGTTGGTACTTCTTTGAAAGATT;MAPQ=60;MATEID=4461382_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_132741001_132766001_482C;SPAN=16230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:31 GQ:24.8 PL:[24.8, 0.0, 47.9] SR:10 DR:0 LR:-24.61 LO:25.11);ALT=C[chr9:132757121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	132757238	+	chr9	132805230	+	.	0	20	4461505_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4461505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_132790001_132815001_140C;SPAN=47992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:25 GQ:0 PL:[59.4, 0.0, 0.0] SR:20 DR:0 LR:-62.61 LO:62.61);ALT=C[chr9:132805230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	133383116	+	chr9	133387421	+	GTGATCC	41	51	4463328_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;INSERTION=GTGATCC;MAPQ=60;MATEID=4463328_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_9_133378001_133403001_411C;SPAN=4305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:71 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:51 DR:41 LR:-254.2 LO:254.2);ALT=C[chr9:133387421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	133570980	+	chr9	133573547	+	ATACATTGGTGAAGTAGGAGACATCGTAGTGGGACGAATCACAG	0	9	4463812_1	0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=ATACATTGGTGAAGTAGGAGACATCGTAGTGGGACGAATCACAG;MAPQ=60;MATEID=4463812_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_133549501_133574501_92C;SPAN=2567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:121 GQ:2.7 PL:[0.0, 2.7, 297.0] SR:9 DR:0 LR:3.073 LO:16.24);ALT=G[chr9:133573547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	134001137	+	chr9	134002909	+	.	10	3	4465529_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4465529_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_133990501_134015501_62C;SPAN=1772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:3 DR:10 LR:-8.627 LO:19.88);ALT=G[chr9:134002909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	134004864	+	chr9	134006152	+	.	0	4	4465538_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4465538_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_133990501_134015501_123C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:108 GQ:15.9 PL:[0.0, 15.9, 293.7] SR:4 DR:0 LR:16.06 LO:5.98);ALT=G[chr9:134006152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	134103720	+	chr9	134106016	+	.	0	15	4465988_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=4465988_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_134088501_134113501_91C;SPAN=2296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:15 DP:313 GQ:35 PL:[0.0, 35.0, 828.5] SR:15 DR:0 LR:35.28 LO:24.13);ALT=T[chr9:134106016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	134106157	+	chr9	134108841	+	GTTCAGCTTTGGGTCAAATAACTC	5	40	4465995_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTTCAGCTTTGGGTCAAATAACTC;MAPQ=60;MATEID=4465995_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_134088501_134113501_120C;SPAN=2684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:106 GQ:99 PL:[110.0, 0.0, 146.3] SR:40 DR:5 LR:-109.9 LO:110.2);ALT=G[chr9:134108841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	134269651	+	chr9	134305475	+	.	5	3	4467102_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4467102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_134284501_134309501_225C;SPAN=35824;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:45 GQ:11 PL:[11.0, 0.0, 96.8] SR:3 DR:5 LR:-10.92 LO:15.02);ALT=G[chr9:134305475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	135224876	+	chr9	135230303	+	.	9	0	4470258_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4470258_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:135224876(+)-9:135230303(-)__9_135215501_135240501D;SPAN=5427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:0 DR:9 LR:-1.533 LO:16.86);ALT=T[chr9:135230303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	135906551	+	chr9	135917473	+	.	0	11	4472658_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4472658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_135901501_135926501_214C;SPAN=10922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:135 GQ:0 PL:[0.0, 0.0, 326.7] SR:11 DR:0 LR:0.2638 LO:20.3);ALT=G[chr9:135917473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136037919	+	chr9	136039139	+	.	0	7	4473251_1	0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=4473251_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_136024001_136049001_135C;SPAN=1220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:105 GQ:5.1 PL:[0.0, 5.1, 264.0] SR:7 DR:0 LR:5.34 LO:12.29);ALT=C[chr9:136039139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136081121	-	chr9	138441408	+	CTTTCACCTACTCCCACGCCCTGCCAGGCCAAGTGAGAATCCTCGGC	6	38	4481010_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;INSERTION=CTTTCACCTACTCCCACGCCCTGCCAGGCCAAGTGAGAATCCTCGGC;MAPQ=39;MATEID=4481010_2;MATENM=1;NM=2;NUMPARTS=3;REPSEQ=TTT;SCTG=c_9_138425001_138450001_232C;SPAN=2360287;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:46 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:38 DR:6 LR:-135.3 LO:135.3);ALT=[chr9:138441408[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr9	136126534	+	chr9	136150576	+	.	15	0	4473685_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4473685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136126534(+)-9:136150576(-)__9_136146501_136171501D;SPAN=24042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:37 GQ:39.5 PL:[39.5, 0.0, 49.4] SR:0 DR:15 LR:-39.49 LO:39.56);ALT=G[chr9:136150576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136221872	+	chr9	136223144	+	.	53	0	4473912_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4473912_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136221872(+)-9:136223144(-)__9_136220001_136245001D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:81 GQ:41 PL:[153.2, 0.0, 41.0] SR:0 DR:53 LR:-156.4 LO:156.4);ALT=G[chr9:136223144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136234361	+	chr9	136242861	+	.	23	0	4473959_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4473959_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136234361(+)-9:136242861(-)__9_136220001_136245001D;SPAN=8500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:89 GQ:51.8 PL:[51.8, 0.0, 164.0] SR:0 DR:23 LR:-51.81 LO:55.07);ALT=C[chr9:136242861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136258365	+	chr16	22133566	+	.	20	58	4474595_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ATGGATGGATGGATGAGTGGATG;MAPQ=60;MATEID=4474595_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_136244501_136269501_153C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:57 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:58 DR:20 LR:-194.7 LO:194.7);ALT=G[chr16:22133566[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr9	136625194	+	chr9	136626268	+	TGGG	0	36	4475156_1	99.0	.	EVDNC=ASSMB;INSERTION=TGGG;MAPQ=60;MATEID=4475156_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_9_136612001_136637001_285C;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:66 GQ:58.1 PL:[101.0, 0.0, 58.1] SR:36 DR:0 LR:-101.5 LO:101.5);ALT=G[chr9:136626268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	136918729	+	chr9	136933066	+	.	14	0	4476342_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4476342_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:136918729(+)-9:136933066(-)__9_136930501_136955501D;SPAN=14337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:5 GQ:3.6 PL:[39.6, 3.6, 0.0] SR:0 DR:14 LR:-39.61 LO:39.61);ALT=A[chr9:136933066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	137001332	+	chr9	137004938	+	.	9	0	4476593_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4476593_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:137001332(+)-9:137004938(-)__9_136979501_137004501D;SPAN=3606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:18 GQ:18.2 PL:[24.8, 0.0, 18.2] SR:0 DR:9 LR:-24.88 LO:24.88);ALT=C[chr9:137004938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	137808310	+	chr9	137809615	+	.	27	10	4479041_1	70.0	.	DISC_MAPQ=49;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=4479041_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_9_137788001_137813001_195C;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:105 GQ:70.7 PL:[70.7, 0.0, 182.9] SR:10 DR:27 LR:-70.58 LO:73.39);ALT=G[chr9:137809615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	138392626	+	chr9	138393688	+	.	16	0	4480711_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4480711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:138392626(+)-9:138393688(-)__9_138376001_138401001D;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:66 GQ:35 PL:[35.0, 0.0, 124.1] SR:0 DR:16 LR:-34.94 LO:37.79);ALT=G[chr9:138393688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	138393821	+	chr9	138395385	+	.	2	6	4480714_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=4480714_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_138376001_138401001_187C;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:6 DR:2 LR:-2.567 LO:15.16);ALT=T[chr9:138395385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	138479103	+	chr9	138480200	+	.	78	48	4481204_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGC;MAPQ=60;MATEID=4481204_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_9_138474001_138499001_134C;SPAN=1097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:102 DP:26 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:48 DR:78 LR:-300.4 LO:300.4);ALT=C[chr9:138480200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139266593	+	chr9	139267985	+	.	13	0	4483794_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4483794_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139266593(+)-9:139267985(-)__9_139258001_139283001D;SPAN=1392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=C[chr9:139267985[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139560321	+	chr9	139563007	+	.	16	0	4484624_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4484624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139560321(+)-9:139563007(-)__9_139552001_139577001D;SPAN=2686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:55 GQ:38 PL:[38.0, 0.0, 94.1] SR:0 DR:16 LR:-37.92 LO:39.29);ALT=G[chr9:139563007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139562778	+	chr9	139564056	+	.	17	0	4484633_1	32.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4484633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139562778(+)-9:139564056(-)__9_139552001_139577001D;SPAN=1278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:89 GQ:32 PL:[32.0, 0.0, 183.8] SR:0 DR:17 LR:-32.01 LO:38.15);ALT=T[chr9:139564056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139572010	+	chr9	139581628	+	.	0	13	4484746_1	32.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4484746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_139576501_139601501_165C;SPAN=9618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:41 GQ:32 PL:[32.0, 0.0, 65.0] SR:13 DR:0 LR:-31.81 LO:32.52);ALT=T[chr9:139581628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139757500	+	chr9	139760662	+	.	18	0	4485709_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4485709_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139757500(+)-9:139760662(-)__9_139748001_139773001D;SPAN=3162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:137 GQ:22.4 PL:[22.4, 0.0, 309.5] SR:0 DR:18 LR:-22.3 LO:37.18);ALT=C[chr9:139760662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139757955	+	chr9	139760649	+	.	136	0	4485715_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4485715_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139757955(+)-9:139760649(-)__9_139748001_139773001D;SPAN=2694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:122 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:0 DR:136 LR:-402.7 LO:402.7);ALT=A[chr9:139760649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139758325	+	chr9	139760632	+	.	53	46	4485717_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=4485717_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_139748001_139773001_145C;SPAN=2307;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:122 GQ:99 PL:[155.3, 0.0, 138.8] SR:46 DR:53 LR:-155.1 LO:155.1);ALT=T[chr9:139760632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139872144	+	chr9	139873443	+	.	0	6	4485877_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4485877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_139870501_139895501_342C;SPAN=1299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:82 GQ:2.1 PL:[0.0, 2.1, 201.3] SR:6 DR:0 LR:2.41 LO:10.78);ALT=G[chr9:139873443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	139927735	+	chr9	139929103	+	.	12	0	4485815_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4485815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:139927735(+)-9:139929103(-)__9_139919501_139944501D;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:92 GQ:14.9 PL:[14.9, 0.0, 206.3] SR:0 DR:12 LR:-14.69 LO:24.74);ALT=C[chr9:139929103[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140135869	+	chr9	140136947	+	TTTTGGGAGGTGATCAGCGATGAGCACGGCATCGACCCCACGGGCACCTACCACGGGGACAGCGACCTGCAGCTGGAACGCATCAACGTGTACTACAATGAGGCCACCGGCGGCAAGTACGTGCCCCGCGCCGTGCTCGTGGATCTGGAGCCCGGCACCATGGACTCCGTGCGCTCGGGGCCCTTCGGGCAGATCTTCCGGCCGGACAACTTCGTTTTC	5	40	4486774_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=TTTTGGGAGGTGATCAGCGATGAGCACGGCATCGACCCCACGGGCACCTACCACGGGGACAGCGACCTGCAGCTGGAACGCATCAACGTGTACTACAATGAGGCCACCGGCGGCAAGTACGTGCCCCGCGCCGTGCTCGTGGATCTGGAGCCCGGCACCATGGACTCCGTGCGCTCGGGGCCCTTCGGGCAGATCTTCCGGCCGGACAACTTCGTTTTC;MAPQ=60;MATEID=4486774_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_9_140115501_140140501_400C;SPAN=1078;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:70 GQ:53.6 PL:[116.3, 0.0, 53.6] SR:40 DR:5 LR:-117.6 LO:117.6);ALT=G[chr9:140136947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140289860	+	chr9	140317566	+	.	3	4	4487169_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGC;MAPQ=60;MATEID=4487169_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140287001_140312001_310C;SPAN=27706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:32 GQ:8 PL:[8.0, 0.0, 67.4] SR:4 DR:3 LR:-7.835 LO:10.74);ALT=C[chr9:140317566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140346697	+	chr9	140344585	+	.	11	0	4487260_1	13.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=4487260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:140344585(-)-9:140346697(+)__9_140336001_140361001D;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:0 DR:11 LR:-13.55 LO:22.7);ALT=]chr9:140346697]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr9	140500224	+	chr9	140507863	+	.	10	0	4488056_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4488056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:140500224(+)-9:140507863(-)__9_140507501_140532501D;SPAN=7639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:0 DR:10 LR:-19.73 LO:22.76);ALT=A[chr9:140507863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140500287	+	chr9	140507346	+	.	57	33	4488057_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4488057_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140507501_140532501_419C;SPAN=7059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:0 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:33 DR:57 LR:-201.3 LO:201.3);ALT=G[chr9:140507346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140513548	+	chr9	140611075	+	.	14	0	4488760_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4488760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:140513548(+)-9:140611075(-)__9_140605501_140630501D;SPAN=97527;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:76 GQ:25.7 PL:[25.7, 0.0, 157.7] SR:0 DR:14 LR:-25.62 LO:31.17);ALT=G[chr9:140611075[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	140783384	+	chr9	140785281	+	.	66	31	4489230_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4489230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_140777001_140802001_444C;SPAN=1897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:173 GQ:99 PL:[240.5, 0.0, 177.8] SR:31 DR:66 LR:-240.8 LO:240.8);ALT=G[chr9:140785281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	2812387	+	chr10	3748412	+	.	11	0	4496763_1	29.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4496763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:2812387(+)-10:3748412(-)__10_3748501_3773501D;SPAN=936025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:2 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:11 LR:-29.71 LO:29.71);ALT=G[chr10:3748412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3109901	+	chr10	3124578	+	.	40	24	4495829_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4495829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3111501_3136501_3C;SPAN=14677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:44 GQ:12 PL:[132.0, 12.0, 0.0] SR:24 DR:40 LR:-132.0 LO:132.0);ALT=T[chr10:3124578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3109931	+	chr10	3141464	+	.	20	0	4495975_1	58.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4495975_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:3109931(+)-10:3141464(-)__10_3136001_3161001D;SPAN=31533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:29 GQ:11.9 PL:[58.1, 0.0, 11.9] SR:0 DR:20 LR:-59.85 LO:59.85);ALT=G[chr10:3141464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3141545	+	chr10	3143556	+	.	0	10	4495984_1	18.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4495984_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3136001_3161001_110C;SPAN=2011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:10 DR:0 LR:-18.65 LO:22.38);ALT=G[chr10:3143556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3357536	+	chr10	3356324	+	.	42	0	4496231_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=4496231_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:3356324(-)-10:3357536(+)__10_3356501_3381501D;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:20 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=]chr10:3357536]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	3822424	+	chr10	3823832	+	.	33	6	4497208_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4497208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3797501_3822501_18C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:6 DR:33 LR:-115.5 LO:115.5);ALT=G[chr10:3823832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	3824410	+	chr10	3827105	+	.	126	139	4496862_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTGT;MAPQ=60;MATEID=4496862_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_3822001_3847001_130C;SPAN=2695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:192 DP:254 GQ:50.2 PL:[565.1, 0.0, 50.2] SR:139 DR:126 LR:-590.1 LO:590.1);ALT=T[chr10:3827105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	4290063	+	chr10	4291683	+	.	74	51	4497691_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4497691_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_10_4287501_4312501_0C;SPAN=1620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:26 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:51 DR:74 LR:-293.8 LO:293.8);ALT=C[chr10:4291683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	4376586	+	chr10	4374452	+	.	39	0	4497876_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4497876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:4374452(-)-10:4376586(+)__10_4361001_4386001D;SPAN=2134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:39 LR:-125.4 LO:125.4);ALT=]chr10:4376586]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	4708518	+	chr10	4710523	+	ATAG	50	42	4498208_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATAG;MAPQ=60;MATEID=4498208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_4704001_4729001_49C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:22 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:42 DR:50 LR:-208.0 LO:208.0);ALT=T[chr10:4710523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5136722	+	chr10	5138608	+	TCCA	23	12	4498895_1	74.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCCA;MAPQ=60;MATEID=4498895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5120501_5145501_121C;SPAN=1886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:53 GQ:51.8 PL:[74.9, 0.0, 51.8] SR:12 DR:23 LR:-74.95 LO:74.95);ALT=T[chr10:5138608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5147869	+	chr10	5149651	+	.	0	11	4498916_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4498916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5145001_5170001_60C;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:11 DR:0 LR:-21.14 LO:24.83);ALT=G[chr10:5149651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5838825	+	chr10	5842561	+	.	0	25	4500010_1	64.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4500010_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5831001_5856001_68C;SPAN=3736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:67 GQ:64.4 PL:[64.4, 0.0, 97.4] SR:25 DR:0 LR:-64.37 LO:64.76);ALT=A[chr10:5842561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5838873	+	chr10	5855175	+	.	8	0	4500011_1	9.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4500011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:5838873(+)-10:5855175(-)__10_5831001_5856001D;SPAN=16302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:0 DR:8 LR:-9.34 LO:16.4);ALT=T[chr10:5855175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5842669	+	chr10	5855176	+	.	0	97	4500021_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4500021_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5831001_5856001_225C;SPAN=12507;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:102 GQ:27.3 PL:[300.3, 27.3, 0.0] SR:97 DR:0 LR:-300.4 LO:300.4);ALT=C[chr10:5855176[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5889586	+	chr10	5892818	+	.	41	34	4500385_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTCTGCCTCCCAGGTTCAAGCAATTCT;MAPQ=45;MATEID=4500385_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5880001_5905001_252C;SPAN=3232;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:21 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:34 DR:41 LR:-188.1 LO:188.1);ALT=T[chr10:5892818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	5969505	+	chr10	5978418	+	.	2	2	4500266_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4500266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_5953501_5978501_202C;SPAN=8913;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:46 GQ:0.8 PL:[0.8, 0.0, 109.7] SR:2 DR:2 LR:-0.7415 LO:7.501);ALT=G[chr10:5978418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	6131108	+	chr15	35591616	-	.	16	0	5924278_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5924278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:6131108(+)-15:35591616(+)__15_35574001_35599001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:30 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:0 DR:16 LR:-44.89 LO:44.89);ALT=C]chr15:35591616];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	6131119	+	chr10	6139007	+	.	39	0	4500777_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4500777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:6131119(+)-10:6139007(-)__10_6125001_6150001D;SPAN=7888;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:50 GQ:6.2 PL:[115.1, 0.0, 6.2] SR:0 DR:39 LR:-121.1 LO:121.1);ALT=C[chr10:6139007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	6156110	+	chr10	6157414	+	TTAATTGCTGATTCAACTCTCTCAAATTCTAAAAATATCCGTACTGCTTCATCATCAGGGGCACCAGGAAT	4	14	4500727_1	40.0	.	DISC_MAPQ=41;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTAATTGCTGATTCAACTCTCTCAAATTCTAAAAATATCCGTACTGCTTCATCATCAGGGGCACCAGGAAT;MAPQ=60;MATEID=4500727_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_6149501_6174501_0C;SPAN=1304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:59 GQ:40.1 PL:[40.1, 0.0, 102.8] SR:14 DR:4 LR:-40.13 LO:41.66);ALT=A[chr10:6157414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	6411580	+	chr10	6417630	+	.	40	24	4501537_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGCAAATCATTTTCCT;MAPQ=60;MATEID=4501537_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_6394501_6419501_193C;SPAN=6050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:139 GQ:99 PL:[147.2, 0.0, 190.1] SR:24 DR:40 LR:-147.2 LO:147.5);ALT=T[chr10:6417630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17396861	+	chr10	7059510	+	.	25	0	6752155_1	75.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6752155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:7059510(-)-19:17396861(+)__19_17395001_17420001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:26 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:0 DR:25 LR:-75.92 LO:75.92);ALT=]chr19:17396861]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	7077040	+	chr10	7078302	+	A	105	72	4502524_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4502524_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_7056001_7081001_305C;SPAN=1262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:37 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:72 DR:105 LR:-432.4 LO:432.4);ALT=T[chr10:7078302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7132876	+	chr19	17397640	+	.	31	28	6752156_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGAA;MAPQ=60;MATEID=6752156_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_17395001_17420001_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:31 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:28 DR:31 LR:-148.5 LO:148.5);ALT=A[chr19:17397640[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	7634373	-	chr18	9868617	+	.	9	18	6538428_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6538428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_9849001_9874001_132C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:40 GQ:28.7 PL:[68.3, 0.0, 28.7] SR:18 DR:9 LR:-69.27 LO:69.27);ALT=[chr18:9868617[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	7723778	+	chr17	746192	+	.	0	35	4503687_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GAAAGAAA;MAPQ=60;MATEID=4503687_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_7717501_7742501_245C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:11 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:35 DR:0 LR:-102.3 LO:102.3);ALT=A[chr17:746192[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	7825176	+	chr10	7829858	+	.	12	0	4503854_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4503854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:7825176(+)-10:7829858(-)__10_7815501_7840501D;SPAN=4682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:63 GQ:22.7 PL:[22.7, 0.0, 128.3] SR:0 DR:12 LR:-22.54 LO:26.91);ALT=T[chr10:7829858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7830227	+	chr10	7839010	+	ATTCAAGTTCGAAATATGGCAACTTTGAAAGATA	116	42	4503874_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GACTAAAGTCCATCAAAAACATCCAGAAAATTACCAAGTCTATGAAAATGGTAGCGGCAGCAAAATATGCCCGAGCTGAGAGAGAGCTGAAACCAGCTCGAATATATGGATTGGGATCTTTAG;INSERTION=ATTCAAGTTCGAAATATGGCAACTTTGAAAGATA;MAPQ=60;MATEID=4503874_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_7815501_7840501_181C;SECONDARY;SPAN=8783;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:97 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:42 DR:116 LR:-415.9 LO:415.9);ALT=G[chr10:7839010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7830256	+	chr10	7840947	+	.	36	0	4503875_1	99.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4503875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:7830256(+)-10:7840947(-)__10_7815501_7840501D;SPAN=10691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:36 LR:-115.5 LO:115.5);ALT=A[chr10:7840947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7839141	+	chr10	7840951	+	.	4	150	4504031_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4504031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_7840001_7865001_205C;SPAN=1810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:153 DP:63 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:150 DR:4 LR:-452.2 LO:452.2);ALT=G[chr10:7840951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	7842054	+	chr10	7844232	+	.	8	11	4504039_1	27.0	.	DISC_MAPQ=51;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=4504039_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_7840001_7865001_254C;SPAN=2178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:80 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:11 DR:8 LR:-27.84 LO:33.52);ALT=G[chr10:7844232[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	11207646	+	chr10	11252632	+	.	0	49	4511845_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4511845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_11196501_11221501_287C;SPAN=44986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:49 DR:0 LR:-155.1 LO:155.1);ALT=G[chr10:11252632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	11207647	+	chr10	11259386	+	.	0	31	4511846_1	88.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=4511846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_11196501_11221501_382C;SPAN=51739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:52 GQ:35.6 PL:[88.4, 0.0, 35.6] SR:31 DR:0 LR:-89.33 LO:89.33);ALT=T[chr10:11259386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12077479	+	chr10	12084753	+	.	42	0	4514265_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12077479(+)-10:12084753(-)__10_12054001_12079001D;SPAN=7274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:42 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=G[chr10:12084753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12209811	+	chr10	12215717	+	ATCAAGTCTCTGCAGCAGGTCATTCTTGGGTAAAGAAATGACTTCCACAAACTCTCCATCCCCTGGCTTTGGCTTCGGCCTTGCGTTTTCGGCATCATCTCCGTTAATGGTGACTGTCACGATGTGTATAGTACAGTTTGACAAGCCTGGGTCCATACAGACCG	0	48	4514812_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATCAAGTCTCTGCAGCAGGTCATTCTTGGGTAAAGAAATGACTTCCACAAACTCTCCATCCCCTGGCTTTGGCTTCGGCCTTGCGTTTTCGGCATCATCTCCGTTAATGGTGACTGTCACGATGTGTATAGTACAGTTTGACAAGCCTGGGTCCATACAGACCG;MAPQ=60;MATEID=4514812_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_10_12201001_12226001_127C;SPAN=5906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:88 GQ:78.5 PL:[134.6, 0.0, 78.5] SR:48 DR:0 LR:-135.4 LO:135.4);ALT=C[chr10:12215717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12215817	+	chr10	12226888	+	GGGAACTCTATGCAGTAGCCCCCCATTGGTGGTCGGAACTGTTTCACCAGAACGATACACTCATAGTGAAGTGTTCTCTGCAGCACGGGGATGACCGCGACACCATCCGCAGTCTGCTCTTTCCTGGTTGTACGTTTCACTGATTCCCAAGTT	0	49	4514830_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GGGAACTCTATGCAGTAGCCCCCCATTGGTGGTCGGAACTGTTTCACCAGAACGATACACTCATAGTGAAGTGTTCTCTGCAGCACGGGGATGACCGCGACACCATCCGCAGTCTGCTCTTTCCTGGTTGTACGTTTCACTGATTCCCAAGTT;MAPQ=60;MATEID=4514830_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_12201001_12226001_11C;SPAN=11071;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:33 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:49 DR:0 LR:-145.2 LO:145.2);ALT=A[chr10:12226888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12219900	+	chr10	12226888	+	ATCCGCAGTCTGCTCTTTCCTGGTTGTACGTTTCACTGATTCCCAAGTT	4	50	4514955_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=ATCCGCAGTCTGCTCTTTCCTGGTTGTACGTTTCACTGATTCCCAAGTT;MAPQ=60;MATEID=4514955_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_12225501_12250501_194C;SPAN=6988;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:45 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:50 DR:4 LR:-158.4 LO:158.4);ALT=C[chr10:12226888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12221181	+	chr10	12237767	+	.	13	0	4514958_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514958_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12221181(+)-10:12237767(-)__10_12225501_12250501D;SPAN=16586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:0 DR:13 LR:-30.18 LO:31.58);ALT=T[chr10:12237767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12226957	+	chr10	12228228	+	.	0	56	4514963_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4514963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_12225501_12250501_148C;SPAN=1271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:56 DP:92 GQ:61.1 PL:[160.1, 0.0, 61.1] SR:56 DR:0 LR:-162.2 LO:162.2);ALT=T[chr10:12228228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12226998	+	chr10	12237766	+	.	33	0	4514964_1	87.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=4514964_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12226998(+)-10:12237766(-)__10_12225501_12250501D;SPAN=10768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:80 GQ:87.2 PL:[87.2, 0.0, 107.0] SR:0 DR:33 LR:-87.26 LO:87.37);ALT=A[chr10:12237766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12228331	+	chr10	12237768	+	.	40	12	4514965_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4514965_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_12225501_12250501_423C;SPAN=9437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:89 GQ:94.7 PL:[121.1, 0.0, 94.7] SR:12 DR:40 LR:-121.3 LO:121.3);ALT=C[chr10:12237768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12238302	+	chr10	12257737	+	.	11	0	4514989_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514989_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12238302(+)-10:12257737(-)__10_12225501_12250501D;SPAN=19435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:0 DR:11 LR:-25.75 LO:26.84);ALT=G[chr10:12257737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12238316	+	chr10	12251963	+	.	31	0	4514990_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4514990_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:12238316(+)-10:12251963(-)__10_12225501_12250501D;SPAN=13647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=G[chr10:12251963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12238318	+	chr10	12240702	+	.	25	13	4514991_1	69.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4514991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_12225501_12250501_285C;SPAN=2384;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:72 GQ:69.8 PL:[69.8, 0.0, 102.8] SR:13 DR:25 LR:-69.62 LO:70.02);ALT=G[chr10:12240702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12240776	+	chr10	12257738	+	GATGATCCACCAACACATTCTCAGCCAGACAGTGATGATGAAGCAGAAGAAATACAGTGGTCTGATGATGAGAACACAGCCACGCTTAC	0	61	4514997_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GATGATCCACCAACACATTCTCAGCCAGACAGTGATGATGAAGCAGAAGAAATACAGTGGTCTGATGATGAGAACACAGCCACGCTTAC;MAPQ=60;MATEID=4514997_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_12225501_12250501_118C;SPAN=16962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:41 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:61 DR:0 LR:-178.2 LO:178.2);ALT=G[chr10:12257738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12391909	+	chr10	12595224	+	.	10	11	4516003_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4516003_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_12593001_12618001_174C;SPAN=203315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:39 GQ:45.5 PL:[48.8, 0.0, 45.5] SR:11 DR:10 LR:-48.86 LO:48.86);ALT=C[chr10:12595224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	12560473	+	chr10	12562974	+	.	79	58	4516315_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTTATTCATTCTT;MAPQ=60;MATEID=4516315_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_10_12544001_12569001_147C;SPAN=2501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:35 GQ:27 PL:[297.0, 27.0, 0.0] SR:58 DR:79 LR:-297.1 LO:297.1);ALT=T[chr10:12562974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	13337651	+	chr10	13342000	+	.	8	0	4518561_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4518561_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:13337651(+)-10:13342000(-)__10_13328001_13353001D;SPAN=4349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=A[chr10:13342000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	13629153	+	chr10	13639457	+	.	0	8	4519288_1	3.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4519288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_13622001_13647001_72C;SPAN=10304;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:8 DR:0 LR:-3.109 LO:15.25);ALT=G[chr10:13639457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	13652186	+	chr10	13653613	+	.	3	6	4519387_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4519387_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_13646501_13671501_170C;SPAN=1427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:6 DR:3 LR:3.764 LO:10.62);ALT=G[chr10:13653613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	14880459	+	chr10	14881902	+	.	11	7	4522544_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=4522544_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_10_14871501_14896501_333C;SPAN=1443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:73 GQ:29.9 PL:[29.9, 0.0, 145.4] SR:7 DR:11 LR:-29.74 LO:34.19);ALT=G[chr10:14881902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	8126012	+	chr10	15373880	+	.	2	11	4523962_1	33.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=ATATATATATATATAT;MAPQ=60;MATEID=4523962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_15361501_15386501_136C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:12 DP:10 GQ:3 PL:[33.0, 3.0, 0.0] SR:11 DR:2 LR:-33.01 LO:33.01);ALT=]chr18:8126012]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	22209894	+	chr10	22292141	+	CTGCCTTCGTTCATCATCCTTTAAAACTTCATAAATGGCCACCAATTGTCTAAACTGAGTTTCTGCATTTTCATCTTTATTCTTGTCTGGATGTAAAGTTAGTGAAAGCTTACGATATGCTTTTCTGATGTCTGCAGATGATGCAT	0	30	4540441_1	85.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=CTGCCTTCGTTCATCATCCTTTAAAACTTCATAAATGGCCACCAATTGTCTAAACTGAGTTTCTGCATTTTCATCTTTATTCTTGTCTGGATGTAAAGTTAGTGAAAGCTTACGATATGCTTTTCTGATGTCTGCAGATGATGCAT;MAPQ=60;MATEID=4540441_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_22197001_22222001_26C;SPAN=82247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:52 GQ:38.9 PL:[85.1, 0.0, 38.9] SR:30 DR:0 LR:-85.76 LO:85.76);ALT=T[chr10:22292141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	22218073	+	chr10	22292141	+	.	0	11	4540674_1	25.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=4540674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_22270501_22295501_77C;SPAN=74068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:11 DR:0 LR:-25.75 LO:26.84);ALT=G[chr10:22292141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	22605441	+	chr10	22607030	+	.	13	0	4541157_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4541157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:22605441(+)-10:22607030(-)__10_22589001_22614001D;SPAN=1589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:71 GQ:23.9 PL:[23.9, 0.0, 146.0] SR:0 DR:13 LR:-23.68 LO:28.9);ALT=C[chr10:22607030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	22605485	+	chr10	22606809	+	.	35	27	4541158_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTAG;MAPQ=60;MATEID=4541158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_22589001_22614001_239C;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:68 GQ:17.9 PL:[146.6, 0.0, 17.9] SR:27 DR:35 LR:-152.4 LO:152.4);ALT=G[chr10:22606809[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	23384656	+	chr10	23393070	+	.	0	10	4543119_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=4543119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_23373001_23398001_137C;SPAN=8414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:93 GQ:8 PL:[8.0, 0.0, 215.9] SR:10 DR:0 LR:-7.814 LO:19.72);ALT=G[chr10:23393070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	23393173	+	chr10	23399170	+	.	0	11	4543146_1	25.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4543146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_23373001_23398001_90C;SPAN=5997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:42 GQ:25.1 PL:[25.1, 0.0, 74.6] SR:11 DR:0 LR:-24.93 LO:26.41);ALT=G[chr10:23399170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	23408380	+	chr10	23409683	+	.	0	17	4543200_1	33.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=4543200_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_23397501_23422501_209C;SPAN=1303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:17 DR:0 LR:-33.63 LO:38.73);ALT=G[chr10:23409683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26727385	+	chr10	26781254	+	GGCCTTCCTTGCACCTCGGAGCAAAGCAGCTCGGATAGCGCCACACGTCTGCGCCCTGCGTGGGAAGGGCAGGGCTGACAGCACTTCCTCCCCGGGGCAGAGACCTGGAGCCCGGGTGCGGCAGTCTGCACCGCGCGTCGCTTTCCCGGCCGGAGCCTCGCCGCCTTCCCGCGCCCCGCAGCGCCCCGCAGAGCAGTCG	5	19	4551031_1	50.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GGCCTTCCTTGCACCTCGGAGCAAAGCAGCTCGGATAGCGCCACACGTCTGCGCCCTGCGTGGGAAGGGCAGGGCTGACAGCACTTCCTCCCCGGGGCAGAGACCTGGAGCCCGGGTGCGGCAGTCTGCACCGCGCGTCGCTTTCCCGGCCGGAGCCTCGCCGCCTTCCCGCGCCCCGCAGCGCCCCGCAGAGCAGTCG;MAPQ=60;MATEID=4551031_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_26778501_26803501_326C;SPAN=53869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:44 GQ:50.9 PL:[50.9, 0.0, 54.2] SR:19 DR:5 LR:-50.8 LO:50.81);ALT=G[chr10:26781254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26727782	+	chr10	26781254	+	.	11	10	4551032_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=4551032_2;MATENM=0;NM=3;NUMPARTS=3;SCTG=c_10_26778501_26803501_326C;SPAN=53472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:10 DR:11 LR:-44.2 LO:44.37);ALT=G[chr10:26781254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26727799	+	chr10	26785227	+	.	17	0	4551033_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4551033_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:26727799(+)-10:26785227(-)__10_26778501_26803501D;SPAN=57428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:39 GQ:45.5 PL:[45.5, 0.0, 48.8] SR:0 DR:17 LR:-45.55 LO:45.56);ALT=G[chr10:26785227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26781327	+	chr10	26785230	+	.	0	18	4551047_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=4551047_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_26778501_26803501_169C;SPAN=3903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:80 GQ:37.7 PL:[37.7, 0.0, 156.5] SR:18 DR:0 LR:-37.74 LO:41.84);ALT=G[chr10:26785230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26785320	+	chr10	26789747	+	.	3	11	4551058_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4551058_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_26778501_26803501_201C;SPAN=4427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:11 DR:3 LR:-23.73 LO:30.57);ALT=G[chr10:26789747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26790041	+	chr10	26800674	+	AAGAGGAAGAAGCCCAAGCCAAGGCTGATAAAATTAAGCTGGCGCTGGAAAAACTGAAGGAGGCCAAGGTTAAGA	0	15	4551074_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAGAGGAAGAAGCCCAAGCCAAGGCTGATAAAATTAAGCTGGCGCTGGAAAAACTGAAGGAGGCCAAGGTTAAGA;MAPQ=60;MATEID=4551074_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_26778501_26803501_86C;SPAN=10633;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:75 GQ:29.3 PL:[29.3, 0.0, 151.4] SR:15 DR:0 LR:-29.2 LO:34.0);ALT=G[chr10:26800674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26800835	+	chr10	26802467	+	.	0	12	4551099_1	22.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4551099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_26778501_26803501_192C;SPAN=1632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:65 GQ:22.1 PL:[22.1, 0.0, 134.3] SR:12 DR:0 LR:-22.0 LO:26.73);ALT=G[chr10:26802467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26849774	+	chr10	26851252	+	.	0	4	4551315_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=4551315_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_26827501_26852501_35C;SPAN=1478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:4 DR:0 LR:6.574 LO:6.671);ALT=G[chr10:26851252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	26999048	+	chr10	27002154	+	.	89	35	4551675_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=GAGGTTGCAGTGAGCCGAGATCACGCCATTGCA;MAPQ=0;MATEID=4551675_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_26999001_27024001_99C;SECONDARY;SPAN=3106;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:35 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:35 DR:89 LR:-320.2 LO:320.2);ALT=A[chr10:27002154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27112237	+	chr10	27149675	+	.	32	26	4552106_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4552106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_27146001_27171001_69C;SPAN=37438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:26 DR:32 LR:-128.7 LO:128.7);ALT=G[chr10:27149675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27192516	+	chr10	27601219	-	.	17	0	4553497_1	49.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=4553497_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:27192516(+)-10:27601219(+)__10_27587001_27612001D;SPAN=408703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:5 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:17 LR:-49.51 LO:49.51);ALT=A]chr10:27601219];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	27224203	+	chr10	27228086	+	.	107	79	4552299_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=4552299_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_10_27219501_27244501_51C;SPAN=3883;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:51 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:79 DR:107 LR:-445.6 LO:445.6);ALT=A[chr10:27228086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27229307	+	chr10	27224628	+	GATCCCGCCAAGGATGGCCGCCTCTCCACACCCGGGCTGGAATAAGAGTG	12	20	4552303_1	82.0	.	DISC_MAPQ=50;EVDNC=TSI_G;HOMSEQ=GCAGTGTCTGACATTCATAGAACCCCCTTTCCCCCATAATCTCTGAAACACTAACAAACTGGAAATAAG;INSERTION=GATCCCGCCAAGGATGGCCGCCTCTCCACACCCGGGCTGGAATAAGAGTG;MAPQ=60;MATEID=4552303_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_27219501_27244501_158C;SECONDARY;SPAN=4679;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:38 GQ:9.5 PL:[82.1, 0.0, 9.5] SR:20 DR:12 LR:-85.39 LO:85.39);ALT=]chr10:27229307]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	27403538	+	chr10	27404989	+	.	0	7	4552849_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=39;MATEID=4552849_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_27391001_27416001_63C;SPAN=1451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:7 DR:0 LR:-0.8912 LO:13.07);ALT=T[chr10:27404989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27437971	+	chr10	27443105	+	.	17	16	4552878_1	66.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4552878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_27440001_27465001_61C;SPAN=5134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:35 GQ:17 PL:[66.5, 0.0, 17.0] SR:16 DR:17 LR:-67.94 LO:67.94);ALT=T[chr10:27443105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	27775891	+	chr12	11191370	-	CGTATAAGTACTGGGACTTTTTTTTTT	8	27	5094303_1	92.0	.	DISC_MAPQ=37;EVDNC=ASDIS;INSERTION=CGTATAAGTACTGGGACTTTTTTTTTT;MAPQ=60;MATEID=5094303_2;MATENM=11;NM=3;NUMPARTS=2;SCTG=c_12_11172001_11197001_178C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:49 GQ:26.3 PL:[92.3, 0.0, 26.3] SR:27 DR:8 LR:-94.38 LO:94.38);ALT=A]chr12:11191370];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	27793366	+	chr10	27798801	+	.	8	2	4553786_1	10.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4553786_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_27783001_27808001_276C;SPAN=5435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:2 DR:8 LR:-10.52 LO:20.25);ALT=G[chr10:27798801[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	28527717	+	chr10	28591839	+	.	9	0	4555788_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4555788_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:28527717(+)-10:28591839(-)__10_28591501_28616501D;SPAN=64122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:0 DR:9 LR:-21.04 LO:21.94);ALT=A[chr10:28591839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	28663803	+	chr10	28665096	+	CCCAAGTAGCCTCCCAAGTAGCCTCCCAAG	27	27	4556263_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;INSERTION=CCCAAGTAGCCTCCCAAGTAGCCTCCCAAG;MAPQ=60;MATEID=4556263_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_28640501_28665501_280C;SPAN=1293;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:64 GQ:15.8 PL:[137.9, 0.0, 15.8] SR:27 DR:27 LR:-143.2 LO:143.2);ALT=T[chr10:28665096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	28677208	-	chr10	28678259	+	.	8	0	4556061_1	8.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4556061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:28677208(-)-10:28678259(-)__10_28665001_28690001D;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:0 DR:8 LR:-7.985 LO:16.11);ALT=[chr10:28678259[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	29975581	+	chr10	30024684	+	.	5	6	4560007_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4560007_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_30012501_30037501_208C;SPAN=49103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:23 GQ:23.6 PL:[23.6, 0.0, 30.2] SR:6 DR:5 LR:-23.48 LO:23.56);ALT=C[chr10:30024684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	30630571	+	chr10	30638047	+	.	5	11	4561707_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4561707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_30625001_30650001_384C;SPAN=7476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:80 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:11 DR:5 LR:-27.84 LO:33.52);ALT=T[chr10:30638047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	30723307	+	chr10	30727843	+	.	0	11	4562089_1	19.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4562089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_30698501_30723501_291C;SPAN=4536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:11 DR:0 LR:-19.51 LO:24.29);ALT=G[chr10:30727843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	30723677	+	chr10	30727844	+	.	38	3	4561932_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4561932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_30723001_30748001_156C;SPAN=4167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:98 GQ:99 PL:[108.8, 0.0, 128.6] SR:3 DR:38 LR:-108.8 LO:108.9);ALT=G[chr10:30727844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	30723705	+	chr10	30725849	+	.	11	0	4561933_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4561933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:30723705(+)-10:30725849(-)__10_30723001_30748001D;SPAN=2144;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:88 GQ:12.5 PL:[12.5, 0.0, 200.6] SR:0 DR:11 LR:-12.47 LO:22.46);ALT=C[chr10:30725849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	31443368	+	chr10	31444865	+	.	77	42	4564183_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=TTGGGAGGCTGAGGCAGG;MAPQ=60;MATEID=4564183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_31433501_31458501_235C;SPAN=1497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:51 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:42 DR:77 LR:-277.3 LO:277.3);ALT=G[chr10:31444865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	32324924	+	chr10	32326180	+	.	11	4	4566423_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4566423_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_32315501_32340501_242C;SPAN=1256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:4 DR:11 LR:-26.49 LO:33.08);ALT=T[chr10:32326180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	33221577	+	chr10	33247072	+	.	9	0	4568469_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4568469_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:33221577(+)-10:33247072(-)__10_33197501_33222501D;SPAN=25495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=G[chr10:33247072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	33386453	+	chr10	36119061	+	.	9	19	4573146_1	64.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=4573146_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_10_36113001_36138001_13C;SPAN=2732608;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:29 GQ:5.3 PL:[64.7, 0.0, 5.3] SR:19 DR:9 LR:-67.69 LO:67.69);ALT=T[chr10:36119061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	35248436	+	chr10	35255023	+	.	90	52	4571671_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4571671_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_10_35255501_35280501_292C;SPAN=6587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:0 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:52 DR:90 LR:-326.8 LO:326.8);ALT=G[chr10:35255023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	36148491	-	chr10	36302201	+	.	17	0	4573605_1	49.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=4573605_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:36148491(-)-10:36302201(-)__10_36284501_36309501D;SPAN=153710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:13 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:17 LR:-49.51 LO:49.51);ALT=[chr10:36302201[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	36420084	+	chr12	86504056	-	.	3	9	5274534_1	33.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=ATATATATAGACTATATATATA;MAPQ=60;MATEID=5274534_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_86485001_86510001_196C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:12 GQ:3 PL:[33.0, 3.0, 0.0] SR:9 DR:3 LR:-33.01 LO:33.01);ALT=T]chr12:86504056];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	37874848	+	chr10	36684296	+	.	16	0	4575971_1	49.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4575971_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:36684296(-)-10:37874848(+)__10_37852501_37877501D;SPAN=1190552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:17 GQ:4.5 PL:[49.5, 4.5, 0.0] SR:0 DR:16 LR:-49.51 LO:49.51);ALT=]chr10:37874848]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	37916288	-	chr10	37917420	+	.	12	0	4576107_1	27.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4576107_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:37916288(-)-10:37917420(-)__10_37901501_37926501D;SPAN=1132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:46 GQ:27.2 PL:[27.2, 0.0, 83.3] SR:0 DR:12 LR:-27.15 LO:28.79);ALT=[chr10:37917420[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	38310372	-	chr10	43123587	+	.	16	0	4581075_1	44.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4581075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38310372(-)-10:43123587(-)__10_43120001_43145001D;SPAN=4813215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:31 GQ:28.1 PL:[44.6, 0.0, 28.1] SR:0 DR:16 LR:-44.55 LO:44.55);ALT=[chr10:43123587[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	38645417	+	chr10	38647237	+	.	18	3	4577296_1	50.0	.	DISC_MAPQ=12;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=32;MATEID=4577296_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_38636501_38661501_125C;SPAN=1820;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:56 GQ:50.9 PL:[50.9, 0.0, 83.9] SR:3 DR:18 LR:-50.85 LO:51.32);ALT=G[chr10:38647237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	38778219	+	chr10	38776832	+	.	20	0	4577995_1	45.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=4577995_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38776832(-)-10:38778219(+)__10_38759001_38784001D;SPAN=1387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:76 GQ:45.5 PL:[45.5, 0.0, 137.9] SR:0 DR:20 LR:-45.43 LO:48.08);ALT=]chr10:38778219]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38783026	+	chr10	38781513	+	.	10	0	4578019_1	16.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4578019_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38781513(-)-10:38783026(+)__10_38759001_38784001D;SPAN=1513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.48 LO:21.7);ALT=]chr10:38783026]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38790808	+	chr10	38788969	+	.	9	0	4578527_1	11.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=4578527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38788969(-)-10:38790808(+)__10_38783501_38808501D;SPAN=1839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:0 DR:9 LR:-11.83 LO:18.75);ALT=]chr10:38790808]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38795208	+	chr10	38791686	+	.	8	0	4578543_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4578543_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38791686(-)-10:38795208(+)__10_38783501_38808501D;SPAN=3522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=]chr10:38795208]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38799034	+	chr10	38795559	+	.	10	0	4578564_1	10.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4578564_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38795559(-)-10:38799034(+)__10_38783501_38808501D;SPAN=3475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:0 DR:10 LR:-9.982 LO:20.14);ALT=]chr10:38799034]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38805168	+	chr10	38802842	+	.	13	0	4578626_1	25.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4578626_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38802842(-)-10:38805168(+)__10_38783501_38808501D;SPAN=2326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:65 GQ:25.4 PL:[25.4, 0.0, 131.0] SR:0 DR:13 LR:-25.3 LO:29.46);ALT=]chr10:38805168]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38805788	+	chr10	38802860	+	.	8	0	4578627_1	10.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4578627_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38802860(-)-10:38805788(+)__10_38783501_38808501D;SPAN=2928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=]chr10:38805788]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38871438	+	chr10	38869227	+	.	9	0	4578430_1	12.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=4578430_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38869227(-)-10:38871438(+)__10_38857001_38882001D;SPAN=2211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:0 DR:9 LR:-12.1 LO:18.81);ALT=]chr10:38871438]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	38876414	+	chr10	38875112	+	.	11	0	4578466_1	12.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4578466_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:38875112(-)-10:38876414(+)__10_38857001_38882001D;SPAN=1302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:0 DR:11 LR:-12.74 LO:22.52);ALT=]chr10:38876414]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39078602	+	chr10	39077454	+	.	11	0	4578908_1	23.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=4578908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39077454(-)-10:39078602(+)__10_39077501_39102501D;SPAN=1148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:0 DR:11 LR:-23.85 LO:25.91);ALT=]chr10:39078602]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39079801	+	chr10	39078784	+	.	12	0	4578918_1	19.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=4578918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39078784(-)-10:39079801(+)__10_39077501_39102501D;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:74 GQ:19.7 PL:[19.7, 0.0, 158.3] SR:0 DR:12 LR:-19.56 LO:25.98);ALT=]chr10:39079801]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39081733	+	chr10	39080263	+	.	12	0	4578927_1	16.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=4578927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39080263(-)-10:39081733(+)__10_39077501_39102501D;SPAN=1470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:85 GQ:16.7 PL:[16.7, 0.0, 188.3] SR:0 DR:12 LR:-16.58 LO:25.19);ALT=]chr10:39081733]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39090757	+	chr10	39087832	+	.	16	0	4578962_1	30.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4578962_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39087832(-)-10:39090757(+)__10_39077501_39102501D;SPAN=2925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:82 GQ:30.8 PL:[30.8, 0.0, 166.1] SR:0 DR:16 LR:-30.6 LO:36.07);ALT=]chr10:39090757]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39103265	+	chr10	39101962	+	.	9	0	4579075_1	8.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=4579075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39101962(-)-10:39103265(+)__10_39102001_39127001D;SPAN=1303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:0 DR:9 LR:-8.306 LO:17.99);ALT=]chr10:39103265]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39107791	+	chr10	39106533	+	.	9	0	4579097_1	5.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4579097_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39106533(-)-10:39107791(+)__10_39102001_39127001D;SPAN=1258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:0 DR:9 LR:-5.597 LO:17.5);ALT=]chr10:39107791]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39108429	+	chr10	39106602	+	.	12	0	4579098_1	19.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=4579098_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39106602(-)-10:39108429(+)__10_39102001_39127001D;SPAN=1827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:74 GQ:19.7 PL:[19.7, 0.0, 158.3] SR:0 DR:12 LR:-19.56 LO:25.98);ALT=]chr10:39108429]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39117164	+	chr10	39114067	+	.	10	0	4579143_1	16.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4579143_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39114067(-)-10:39117164(+)__10_39102001_39127001D;SPAN=3097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:0 DR:10 LR:-16.21 LO:21.62);ALT=]chr10:39117164]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39115169	+	chr10	39114108	+	.	8	0	4579149_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4579149_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39114108(-)-10:39115169(+)__10_39102001_39127001D;SPAN=1061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:153 GQ:14.8 PL:[0.0, 14.8, 399.3] SR:0 DR:8 LR:15.04 LO:13.18);ALT=]chr10:39115169]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39124571	+	chr10	39123134	+	.	21	0	4579188_1	44.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4579188_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39123134(-)-10:39124571(+)__10_39102001_39127001D;SPAN=1437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:92 GQ:44.6 PL:[44.6, 0.0, 176.6] SR:0 DR:21 LR:-44.4 LO:48.97);ALT=]chr10:39124571]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39130090	+	chr10	39128976	+	.	9	0	4579711_1	10.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4579711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39128976(-)-10:39130090(+)__10_39126501_39151501D;SPAN=1114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:0 DR:9 LR:-10.2 LO:18.38);ALT=]chr10:39130090]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39140646	+	chr10	39139249	+	.	11	0	4579786_1	18.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4579786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39139249(-)-10:39140646(+)__10_39126501_39151501D;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:0 DR:11 LR:-18.7 LO:24.04);ALT=]chr10:39140646]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39145368	+	chr10	39144044	+	.	10	0	4579823_1	13.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4579823_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39144044(-)-10:39145368(+)__10_39126501_39151501D;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:72 GQ:13.7 PL:[13.7, 0.0, 158.9] SR:0 DR:10 LR:-13.5 LO:20.92);ALT=]chr10:39145368]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39147532	+	chr10	39146496	+	.	18	0	4579831_1	41.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=4579831_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39146496(-)-10:39147532(+)__10_39126501_39151501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:65 GQ:41.9 PL:[41.9, 0.0, 114.5] SR:0 DR:18 LR:-41.81 LO:43.74);ALT=]chr10:39147532]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39150621	+	chr10	39149167	+	.	10	0	4579844_1	9.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4579844_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39149167(-)-10:39150621(+)__10_39126501_39151501D;SPAN=1454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:0 DR:10 LR:-9.711 LO:20.09);ALT=]chr10:39150621]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	39154178	+	chr10	39153114	+	.	10	0	4578694_1	15.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4578694_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:39153114(-)-10:39154178(+)__10_39151001_39176001D;SPAN=1064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:66 GQ:15.2 PL:[15.2, 0.0, 143.9] SR:0 DR:10 LR:-15.13 LO:21.33);ALT=]chr10:39154178]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42356560	+	chr10	42355518	+	.	9	0	4578821_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=4578821_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42355518(-)-10:42356560(+)__10_42336001_42361001D;SPAN=1042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:291 GQ:48.8 PL:[0.0, 48.8, 802.0] SR:0 DR:9 LR:49.13 LO:12.75);ALT=]chr10:42356560]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42665019	+	chr10	42661689	+	.	8	0	4579944_1	7.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4579944_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42661689(-)-10:42665019(+)__10_42654501_42679501D;SPAN=3330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.443 LO:16.0);ALT=]chr10:42665019]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42667527	+	chr10	42666389	+	.	9	0	4579969_1	2.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4579969_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42666389(-)-10:42667527(+)__10_42654501_42679501D;SPAN=1138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:102 GQ:2.3 PL:[2.3, 0.0, 243.2] SR:0 DR:9 LR:-2.075 LO:16.94);ALT=]chr10:42667527]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42792908	+	chr10	42791876	+	.	8	0	4580724_1	4.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=4580724_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42791876(-)-10:42792908(+)__10_42777001_42802001D;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:0 DR:8 LR:-4.192 LO:15.42);ALT=]chr10:42792908]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42809246	+	chr10	42805768	+	.	40	0	4580853_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=4580853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42805768(-)-10:42809246(+)__10_42801501_42826501D;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:70 GQ:56.9 PL:[113.0, 0.0, 56.9] SR:0 DR:40 LR:-114.1 LO:114.1);ALT=]chr10:42809246]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42814392	+	chr10	42812622	+	.	15	0	4580881_1	22.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4580881_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42812622(-)-10:42814392(+)__10_42801501_42826501D;SPAN=1770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:100 GQ:22.4 PL:[22.4, 0.0, 220.4] SR:0 DR:15 LR:-22.42 LO:31.92);ALT=]chr10:42814392]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42815604	+	chr10	42812662	+	.	15	0	4580882_1	33.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4580882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42812662(-)-10:42815604(+)__10_42801501_42826501D;SPAN=2942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:0 DR:15 LR:-33.8 LO:35.92);ALT=]chr10:42815604]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	42816250	+	chr10	42812760	+	.	10	0	4580883_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4580883_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:42812760(-)-10:42816250(+)__10_42801501_42826501D;SPAN=3490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:57 GQ:17.6 PL:[17.6, 0.0, 119.9] SR:0 DR:10 LR:-17.57 LO:22.03);ALT=]chr10:42816250]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	43022099	+	chr10	43290652	+	.	8	0	4581284_1	15.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=4581284_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43022099(+)-10:43290652(-)__10_43267001_43292001D;SPAN=268553;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=A[chr10:43290652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43634035	+	chr10	43650343	+	.	8	0	4582161_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4582161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43634035(+)-10:43650343(-)__10_43634501_43659501D;SPAN=16308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:20 GQ:20.9 PL:[20.9, 0.0, 27.5] SR:0 DR:8 LR:-20.99 LO:21.04);ALT=T[chr10:43650343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43799275	-	chr14	107156050	+	.	10	13	4582418_1	51.0	.	DISC_MAPQ=11;EVDNC=ASDIS;HOMSEQ=CCTGTGAGCTGGCGATCT;MAPQ=25;MATEID=4582418_2;MATENM=2;NM=4;NUMPARTS=2;SCTG=c_10_43781501_43806501_79C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:43 GQ:51.2 PL:[51.2, 0.0, 51.2] SR:13 DR:10 LR:-51.07 LO:51.07);ALT=[chr14:107156050[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	43883386	+	chr10	43890078	+	.	0	67	4582628_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4582628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_43879501_43904501_189C;SPAN=6692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:80 GQ:5.1 PL:[204.6, 5.1, 0.0] SR:67 DR:0 LR:-213.3 LO:213.3);ALT=T[chr10:43890078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43883433	+	chr10	43904574	+	.	28	0	4583002_1	81.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4583002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43883433(+)-10:43904574(-)__10_43904001_43929001D;SPAN=21141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:42 GQ:18.5 PL:[81.2, 0.0, 18.5] SR:0 DR:28 LR:-83.03 LO:83.03);ALT=C[chr10:43904574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43883433	+	chr10	43903162	+	.	17	0	4582629_1	41.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4582629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43883433(+)-10:43903162(-)__10_43879501_43904501D;SPAN=19729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:55 GQ:41.3 PL:[41.3, 0.0, 90.8] SR:0 DR:17 LR:-41.22 LO:42.29);ALT=C[chr10:43903162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43890137	+	chr10	43891903	+	.	2	79	4582645_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4582645_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_43879501_43904501_63C;SPAN=1766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:80 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:79 DR:2 LR:-237.7 LO:237.7);ALT=C[chr10:43891903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43890181	+	chr10	43904574	+	.	20	0	4583003_1	54.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4583003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43890181(+)-10:43904574(-)__10_43904001_43929001D;SPAN=14393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:42 GQ:44.9 PL:[54.8, 0.0, 44.9] SR:0 DR:20 LR:-54.67 LO:54.67);ALT=T[chr10:43904574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43890182	+	chr10	43903162	+	.	23	0	4582647_1	61.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4582647_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43890182(+)-10:43903162(-)__10_43879501_43904501D;SPAN=12980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:55 GQ:61.1 PL:[61.1, 0.0, 71.0] SR:0 DR:23 LR:-61.02 LO:61.08);ALT=A[chr10:43903162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43892036	+	chr10	43904535	+	.	24	0	4583004_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4583004_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43892036(+)-10:43904535(-)__10_43904001_43929001D;SPAN=12499;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:20 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:0 DR:24 LR:-69.32 LO:69.32);ALT=A[chr10:43904535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	43892044	+	chr10	43903163	+	.	31	0	4582649_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4582649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:43892044(+)-10:43903163(-)__10_43879501_43904501D;SPAN=11119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:48 GQ:26.6 PL:[89.3, 0.0, 26.6] SR:0 DR:31 LR:-91.16 LO:91.16);ALT=A[chr10:43903163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	44140249	+	chr10	44141512	+	.	0	11	4583263_1	17.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4583263_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_44124501_44149501_63C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:11 DR:0 LR:-17.89 LO:23.8);ALT=T[chr10:44141512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	44140298	+	chr10	44144245	+	.	9	0	4583264_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4583264_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:44140298(+)-10:44144245(-)__10_44124501_44149501D;SPAN=3947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=T[chr10:44144245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	44141699	+	chr10	44144174	+	.	12	0	4583265_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4583265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:44141699(+)-10:44144174(-)__10_44124501_44149501D;SPAN=2475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=G[chr10:44144174[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	54316902	+	chr10	54320766	+	.	0	32	4599072_1	89.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4599072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_54316501_54341501_171C;SPAN=3864;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:58 GQ:50.3 PL:[89.9, 0.0, 50.3] SR:32 DR:0 LR:-90.5 LO:90.5);ALT=C[chr10:54320766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	54316954	+	chr10	54515099	+	.	9	0	4599313_1	21.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4599313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:54316954(+)-10:54515099(-)__10_54512501_54537501D;SPAN=198145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:30 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.58 LO:22.25);ALT=A[chr10:54515099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	54320878	+	chr10	54515064	+	.	24	7	4599314_1	75.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=4599314_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_54512501_54537501_131C;SPAN=194186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:21 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:7 DR:24 LR:-75.92 LO:75.92);ALT=G[chr10:54515064[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	54483781	+	chr10	54515065	+	.	14	2	4599316_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4599316_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_54512501_54537501_219C;SPAN=31284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:21 GQ:7.7 PL:[40.7, 0.0, 7.7] SR:2 DR:14 LR:-41.52 LO:41.52);ALT=G[chr10:54515065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	60029064	+	chr10	60036875	+	.	7	10	4606374_1	37.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4606374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_60025001_60050001_153C;SPAN=7811;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:56 GQ:37.7 PL:[37.7, 0.0, 97.1] SR:10 DR:7 LR:-37.64 LO:39.14);ALT=G[chr10:60036875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	60477422	+	chr12	72667074	-	G	34	69	5244021_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=5244021_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_72642501_72667501_147C;SPAN=-1;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:57 GQ:25.5 PL:[280.5, 25.5, 0.0] SR:69 DR:34 LR:-280.6 LO:280.6);ALT=G]chr12:72667074];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	61361964	+	chr10	61365009	+	.	47	29	4608151_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AATCA;MAPQ=60;MATEID=4608151_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_61348001_61373001_127C;SPAN=3045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:16 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:29 DR:47 LR:-184.8 LO:184.8);ALT=A[chr10:61365009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	64510899	+	chr19	38299507	+	.	0	37	4612519_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTC;MAPQ=60;MATEID=4612519_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_64508501_64533501_225C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:27 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:37 DR:0 LR:-108.9 LO:108.9);ALT=C[chr19:38299507[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	65024524	+	chr10	65028423	+	.	0	9	4613527_1	18.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4613527_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_65023001_65048001_128C;SPAN=3899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:9 DR:0 LR:-18.33 LO:20.7);ALT=T[chr10:65028423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	65140244	+	chr10	65281495	+	.	15	6	4613928_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=4613928_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_65268001_65293001_25C;SPAN=141251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:15 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:6 DR:15 LR:-52.81 LO:52.81);ALT=T[chr10:65281495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	69833006	+	chr10	69834897	+	.	17	0	4620251_1	42.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4620251_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:69833006(+)-10:69834897(-)__10_69825001_69850001D;SPAN=1891;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:0 DR:17 LR:-42.84 LO:43.35);ALT=A[chr10:69834897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70091992	+	chr10	70096955	+	.	55	14	4620900_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4620900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70070001_70095001_81C;SPAN=4963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:29 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:14 DR:55 LR:-184.8 LO:184.8);ALT=G[chr10:70096955[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70097091	+	chr10	70098258	+	GTTGGAAATCGTGCCAAATGGGATAACATTGACGATGGACTACCAGGGGAGAAGCACAGGGGAGGCCTTCGTGCAGTTTGCTTCAAAGGAGATAGCAGAAAATGCTCTGGGGAAACACAAGGAAAGAATAGGGCAC	3	28	4620800_1	85.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=GTTGGAAATCGTGCCAAATGGGATAACATTGACGATGGACTACCAGGGGAGAAGCACAGGGGAGGCCTTCGTGCAGTTTGCTTCAAAGGAGATAGCAGAAAATGCTCTGGGGAAACACAAGGAAAGAATAGGGCAC;MAPQ=60;MATEID=4620800_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_70094501_70119501_110C;SPAN=1167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:62 GQ:62.6 PL:[85.7, 0.0, 62.6] SR:28 DR:3 LR:-85.68 LO:85.68);ALT=G[chr10:70098258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70097092	+	chr10	70098895	+	.	2	5	4620801_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4620801_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70094501_70119501_6C;SPAN=1803;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:67 GQ:5 PL:[5.0, 0.0, 156.8] SR:5 DR:2 LR:-4.955 LO:13.71);ALT=T[chr10:70098895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70097802	+	chr10	70098895	+	.	10	0	4620806_1	14.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4620806_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:70097802(+)-10:70098895(-)__10_70094501_70119501D;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:0 DR:10 LR:-14.59 LO:21.18);ALT=T[chr10:70098895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70099312	+	chr10	70100931	+	.	4	10	4620809_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4620809_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70094501_70119501_290C;SPAN=1619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:60 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:10 DR:4 LR:-29.96 LO:32.8);ALT=T[chr10:70100931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70099353	+	chr10	70101341	+	.	12	0	4620810_1	24.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4620810_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:70099353(+)-10:70101341(-)__10_70094501_70119501D;SPAN=1988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:56 GQ:24.5 PL:[24.5, 0.0, 110.3] SR:0 DR:12 LR:-24.44 LO:27.6);ALT=C[chr10:70101341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70481082	+	chr10	70482214	+	.	8	0	4621850_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4621850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:70481082(+)-10:70482214(-)__10_70462001_70487001D;SPAN=1132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.59 LO:17.19);ALT=C[chr10:70482214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70481082	+	chr10	70496630	+	.	14	0	4621851_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4621851_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:70481082(+)-10:70496630(-)__10_70462001_70487001D;SPAN=15548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:26 GQ:22.7 PL:[39.2, 0.0, 22.7] SR:0 DR:14 LR:-39.37 LO:39.37);ALT=C[chr10:70496630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70482334	+	chr10	70496631	+	.	0	11	4621854_1	30.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4621854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70462001_70487001_291C;SPAN=14297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:22 GQ:20.6 PL:[30.5, 0.0, 20.6] SR:11 DR:0 LR:-30.4 LO:30.4);ALT=G[chr10:70496631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70525838	+	chr10	70530961	+	.	3	11	4621898_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4621898_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70511001_70536001_104C;SPAN=5123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:57 GQ:27.5 PL:[27.5, 0.0, 110.0] SR:11 DR:3 LR:-27.47 LO:30.31);ALT=T[chr10:70530961[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70661227	+	chr10	70666465	+	.	0	8	4622233_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4622233_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70658001_70683001_182C;SPAN=5238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:77 GQ:5.6 PL:[5.6, 0.0, 180.5] SR:8 DR:0 LR:-5.547 LO:15.65);ALT=G[chr10:70666465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70716068	+	chr10	70719560	+	.	56	32	4622304_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4622304_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70707001_70732001_245C;SPAN=3492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:73 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:32 DR:56 LR:-214.6 LO:214.6);ALT=G[chr10:70719560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70847992	+	chr10	70852819	+	.	9	32	4622673_1	78.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4622673_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70829501_70854501_37C;SPAN=4827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:185 GQ:78.7 PL:[78.7, 0.0, 369.2] SR:32 DR:9 LR:-78.62 LO:89.4);ALT=G[chr10:70852819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70847994	+	chr10	70856838	+	.	128	42	4622876_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4622876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70854001_70879001_121C;SPAN=8844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:142 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:42 DR:128 LR:-419.2 LO:419.2);ALT=T[chr10:70856838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70856987	+	chr10	70863627	+	.	18	54	4622894_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=4622894_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_70854001_70879001_63C;SPAN=6640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:74 DP:275 GQ:99 PL:[169.9, 0.0, 496.7] SR:54 DR:18 LR:-169.8 LO:178.7);ALT=C[chr10:70863627[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70884036	+	chr10	70892653	+	.	14	2	4622712_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4622712_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70878501_70903501_197C;SPAN=8617;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:50 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:2 DR:14 LR:-35.97 LO:37.08);ALT=G[chr10:70892653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	70892808	+	chr10	70915566	+	.	0	9	4622736_1	23.0	.	EVDNC=ASSMB;HOMSEQ=AGGTAAA;MAPQ=60;MATEID=4622736_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_70878501_70903501_243C;SPAN=22758;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:23 GQ:23.6 PL:[23.6, 0.0, 30.2] SR:9 DR:0 LR:-23.48 LO:23.56);ALT=A[chr10:70915566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	71078766	+	chr10	71103581	+	.	0	13	4623270_1	34.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4623270_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_71099001_71124001_77C;SPAN=24815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:33 GQ:34.1 PL:[34.1, 0.0, 44.0] SR:13 DR:0 LR:-33.97 LO:34.07);ALT=G[chr10:71103581[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	71812756	+	chr10	71835354	+	.	16	6	4624493_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4624493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_71834001_71859001_80C;SPAN=22598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:28 GQ:15.5 PL:[51.8, 0.0, 15.5] SR:6 DR:16 LR:-52.87 LO:52.87);ALT=G[chr10:71835354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	71977704	+	chr10	71993084	+	.	16	0	4624932_1	52.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=4624932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:71977704(+)-10:71993084(-)__10_71956501_71981501D;SPAN=15380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:18 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:16 LR:-52.35 LO:52.35);ALT=T[chr10:71993084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72448740	+	chr10	72451335	+	.	7	46	4625763_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TGGCT;MAPQ=60;MATEID=4625763_2;MATENM=1;NM=1;NUMPARTS=4;SCTG=c_10_72446501_72471501_11C;SPAN=2595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:23 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:46 DR:7 LR:-145.2 LO:145.2);ALT=A[chr10:72451335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72642244	+	chr10	72644907	+	.	0	7	4625951_1	12.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4625951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_72642501_72667501_134C;SPAN=2663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:7 DR:0 LR:-12.54 LO:15.5);ALT=T[chr10:72644907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72643807	+	chr10	72644907	+	.	0	39	4625954_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4625954_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_72642501_72667501_202C;SPAN=1100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:75 GQ:72.2 PL:[108.5, 0.0, 72.2] SR:39 DR:0 LR:-108.8 LO:108.8);ALT=T[chr10:72644907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72643852	+	chr10	72648286	+	.	16	0	4625956_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4625956_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:72643852(+)-10:72648286(-)__10_72642501_72667501D;SPAN=4434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:67 GQ:34.7 PL:[34.7, 0.0, 127.1] SR:0 DR:16 LR:-34.66 LO:37.67);ALT=C[chr10:72648286[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72645038	+	chr10	72648286	+	.	43	0	4625960_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4625960_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:72645038(+)-10:72648286(-)__10_72642501_72667501D;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:73 GQ:53 PL:[122.3, 0.0, 53.0] SR:0 DR:43 LR:-123.5 LO:123.5);ALT=T[chr10:72648286[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	72645687	+	chr10	72648287	+	.	55	8	4625962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4625962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_72642501_72667501_263C;SPAN=2600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:83 GQ:23.9 PL:[175.7, 0.0, 23.9] SR:8 DR:55 LR:-182.0 LO:182.0);ALT=C[chr10:72648287[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73511621	+	chr10	73515113	+	TCCATCCGCACCAGCTCCTGGG	3	4	4627447_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCCATCCGCACCAGCTCCTGGG;MAPQ=60;MATEID=4627447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73500001_73525001_152C;SPAN=3492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:53 GQ:5.6 PL:[5.6, 0.0, 121.1] SR:4 DR:3 LR:-5.447 LO:11.98);ALT=G[chr10:73515113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73521785	+	chr10	73533113	+	.	137	78	4627482_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4627482_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73500001_73525001_60C;SPAN=11328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:173 DP:45 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:78 DR:137 LR:-511.6 LO:511.6);ALT=T[chr10:73533113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73577233	+	chr10	73578373	+	.	3	11	4627542_1	31.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4627542_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_10_73573501_73598501_223C;SPAN=1140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:56 GQ:31.1 PL:[31.1, 0.0, 103.7] SR:11 DR:3 LR:-31.04 LO:33.29);ALT=C[chr10:73578373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73577233	+	chr10	73578788	+	ATTGCACTGGGCTGCTGTCTCTGTGTTCTGGCACCAGTAGCTTGGGCCCCATATACACTTCTCAGTTCCCAACAAGGGCTTATGGGCCGAGGGGCAGGCTCCAATTTT	6	17	4627543_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATTGCACTGGGCTGCTGTCTCTGTGTTCTGGCACCAGTAGCTTGGGCCCCATATACACTTCTCAGTTCCCAACAAGGGCTTATGGGCCGAGGGGCAGGCTCCAATTTT;MAPQ=60;MATEID=4627543_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_73573501_73598501_223C;SPAN=1555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:55 GQ:44.6 PL:[44.6, 0.0, 87.5] SR:17 DR:6 LR:-44.52 LO:45.33);ALT=C[chr10:73578788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73579659	+	chr10	73581633	+	CAGTCTTGTTGTTGTCAATCAGCTTGGTCACCTCCTTCACCAGGAATTCACACACCTCACAGTAAACATCAGACTTTGCTGGGACCTCGTGCTT	4	16	4627551_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CAGTCTTGTTGTTGTCAATCAGCTTGGTCACCTCCTTCACCAGGAATTCACACACCTCACAGTAAACATCAGACTTTGCTGGGACCTCGTGCTT;MAPQ=60;MATEID=4627551_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_73573501_73598501_11C;SPAN=1974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:68 GQ:44.3 PL:[44.3, 0.0, 120.2] SR:16 DR:4 LR:-44.3 LO:46.26);ALT=T[chr10:73581633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73581765	+	chr10	73585594	+	.	4	8	4627557_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4627557_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_10_73573501_73598501_240C;SPAN=3829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:78 GQ:15.2 PL:[15.2, 0.0, 173.6] SR:8 DR:4 LR:-15.18 LO:23.09);ALT=C[chr10:73585594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73581765	+	chr10	73587771	+	ATGTGCATCATCATCTGGATAGCAATTTCAGAATACTGGCTGATATAGTTCTTGCA	8	19	4627558_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATGTGCATCATCATCTGGATAGCAATTTCAGAATACTGGCTGATATAGTTCTTGCA;MAPQ=60;MATEID=4627558_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_73573501_73598501_240C;SPAN=6006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:74 GQ:52.7 PL:[52.7, 0.0, 125.3] SR:19 DR:8 LR:-52.57 LO:54.28);ALT=C[chr10:73587771[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73588835	+	chr10	73590883	+	.	2	4	4627578_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4627578_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_10_73573501_73598501_213C;SPAN=2048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:51 GQ:6.2 PL:[6.2, 0.0, 115.1] SR:4 DR:2 LR:-5.989 LO:12.08);ALT=C[chr10:73590883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73588835	+	chr10	73591602	+	ATTTCTCCTTTAATGATGTCCAGGATGACAGGGAGGTAGGAGTCCACTATCTCCTTGCATGAAGCAGACATGTTCGGTTTCGGAAGCCAGTCACAGGTCTTCTCCAAGTAAACAAGGATCTCCT	2	34	4627579_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=ATTTCTCCTTTAATGATGTCCAGGATGACAGGGAGGTAGGAGTCCACTATCTCCTTGCATGAAGCAGACATGTTCGGTTTCGGAAGCCAGTCACAGGTCTTCTCCAAGTAAACAAGGATCTCCT;MAPQ=60;MATEID=4627579_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_73573501_73598501_213C;SPAN=2767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:66 GQ:58.1 PL:[101.0, 0.0, 58.1] SR:34 DR:2 LR:-101.5 LO:101.5);ALT=C[chr10:73591602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73591058	+	chr10	73610945	+	.	14	0	4627815_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4627815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73591058(+)-10:73610945(-)__10_73598001_73623001D;SPAN=19887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:44 GQ:34.4 PL:[34.4, 0.0, 70.7] SR:0 DR:14 LR:-34.29 LO:35.04);ALT=A[chr10:73610945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73591678	+	chr10	73610939	+	ACTGTTGGCTTGTTCCAAACGGTCTGCAGGCAGTGCTTCACTGCCCCGCAGTCGGACGCCGTCTTCACATTCTGGCACCACACTGCCGAGCCCCTGGTGCATTCTTTCAGTCCAAGGACCGGGCCGGCTAGAG	29	65	4627817_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ACTGTTGGCTTGTTCCAAACGGTCTGCAGGCAGTGCTTCACTGCCCCGCAGTCGGACGCCGTCTTCACATTCTGGCACCACACTGCCGAGCCCCTGGTGCATTCTTTCAGTCCAAGGACCGGGCCGGCTAGAG;MAPQ=60;MATEID=4627817_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_10_73598001_73623001_31C;SPAN=19261;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:30 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:65 DR:29 LR:-217.9 LO:217.9);ALT=C[chr10:73610939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73594317	+	chr10	73610945	+	.	60	0	4627819_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4627819_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73594317(+)-10:73610945(-)__10_73598001_73623001D;SPAN=16628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:44 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=C[chr10:73610945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73970591	+	chr10	73972944	+	.	0	8	4628437_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4628437_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_138C;SPAN=2353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:8 DR:0 LR:-10.69 LO:16.71);ALT=T[chr10:73972944[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73973102	+	chr10	73975973	+	.	13	0	4628442_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4628442_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73973102(+)-10:73975973(-)__10_73965501_73990501D;SPAN=2871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:56 GQ:27.8 PL:[27.8, 0.0, 107.0] SR:0 DR:13 LR:-27.74 LO:30.42);ALT=A[chr10:73975973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975896	+	chr10	73990122	+	.	25	3	4628451_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4628451_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_105C;SPAN=14226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:78 GQ:61.4 PL:[61.4, 0.0, 127.4] SR:3 DR:25 LR:-61.39 LO:62.68);ALT=G[chr10:73990122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975898	+	chr10	73979810	+	.	17	6	4628452_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4628452_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_209C;SPAN=3912;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:58 GQ:50.3 PL:[50.3, 0.0, 89.9] SR:6 DR:17 LR:-50.31 LO:50.93);ALT=T[chr10:73979810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975946	+	chr10	73983639	+	.	71	0	4628454_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4628454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73975946(+)-10:73983639(-)__10_73965501_73990501D;SPAN=7693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:58 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=T[chr10:73983639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73975992	+	chr10	73992757	+	.	33	0	4628455_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4628455_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:73975992(+)-10:73992757(-)__10_73965501_73990501D;SPAN=16765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:39 GQ:3.9 PL:[102.3, 3.9, 0.0] SR:0 DR:33 LR:-105.5 LO:105.5);ALT=T[chr10:73992757[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73980137	+	chr10	73983645	+	.	3	5	4628458_1	7.0	.	DISC_MAPQ=20;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4628458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_193C;SPAN=3508;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:57 GQ:7.7 PL:[7.7, 0.0, 129.8] SR:5 DR:3 LR:-7.664 LO:14.24);ALT=G[chr10:73983645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73983814	+	chr10	73990122	+	.	0	79	4628475_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4628475_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_207C;SPAN=6308;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:91 GQ:17.7 PL:[254.1, 17.7, 0.0] SR:79 DR:0 LR:-255.3 LO:255.3);ALT=G[chr10:73990122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	73990198	+	chr10	73992758	+	.	2	65	4628490_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4628490_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_73965501_73990501_241C;SPAN=2560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:35 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:65 DR:2 LR:-194.7 LO:194.7);ALT=G[chr10:73992758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	74322823	+	chr10	74326390	+	.	0	10	4629011_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4629011_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_74308501_74333501_72C;SPAN=3567;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:10 DR:0 LR:-16.75 LO:21.78);ALT=T[chr10:74326390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	74326552	+	chr10	74385767	+	.	14	2	4629082_1	43.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4629082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_74382001_74407001_100C;SPAN=59215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:35 GQ:40.1 PL:[43.4, 0.0, 40.1] SR:2 DR:14 LR:-43.34 LO:43.34);ALT=C[chr10:74385767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	74382031	+	chr10	74385767	+	.	8	0	4629156_1	19.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=4629156_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:74382031(+)-10:74385767(-)__10_74357501_74382501D;SPAN=3736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:26 GQ:19.4 PL:[19.4, 0.0, 42.5] SR:0 DR:8 LR:-19.36 LO:19.88);ALT=G[chr10:74385767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	32673414	+	chr10	74767593	+	AAACATAACACCTAGATACATCC	42	83	6372196_1	99.0	.	DISC_MAPQ=48;EVDNC=ASDIS;INSERTION=AAACATAACACCTAGATACATCC;MAPQ=60;MATEID=6372196_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_17_32658501_32683501_14C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:25 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:83 DR:42 LR:-340.0 LO:340.0);ALT=]chr17:32673414]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	74767593	-	chr17	32673409	+	ATACATCC	44	67	6372195_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;INSERTION=ATACATCC;MAPQ=57;MATEID=6372195_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_32658501_32683501_57C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:23 GQ:27 PL:[297.0, 27.0, 0.0] SR:67 DR:44 LR:-297.1 LO:297.1);ALT=[chr17:32673409[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	74833597	+	chr10	74856520	+	.	9	0	4630067_1	23.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4630067_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:74833597(+)-10:74856520(-)__10_74847501_74872501D;SPAN=22923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=A[chr10:74856520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	74834663	+	chr10	74856520	+	.	10	0	4630068_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4630068_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:74834663(+)-10:74856520(-)__10_74847501_74872501D;SPAN=21857;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:22 GQ:23.9 PL:[27.2, 0.0, 23.9] SR:0 DR:10 LR:-27.05 LO:27.05);ALT=G[chr10:74856520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75148176	+	chr10	75156277	+	.	0	8	4630552_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CTGA;MAPQ=60;MATEID=4630552_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_75141501_75166501_167C;SPAN=8101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:8 DR:0 LR:-13.4 LO:17.42);ALT=A[chr10:75156277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75157034	+	chr10	75160561	+	CCGGGATAGGATGGAGCTCCCCCTGGCTGTGGGGCACCAGGATAGCCTCCAGGGGCTGGATAACCTCCAGGCGCAGGGTAGCCTCCAGCTCCTGGGTAGCCACTACTTGGCACTTGTGGGTAGGCACCTCCTCCCATTGGAGGAAAGCCACTAGGATAAGGATACTGACCAGAAGGGGGAAAAGATGACTCCTGACCTGCAGG	5	31	4630563_1	90.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCGGGATAGGATGGAGCTCCCCCTGGCTGTGGGGCACCAGGATAGCCTCCAGGGGCTGGATAACCTCCAGGCGCAGGGTAGCCTCCAGCTCCTGGGTAGCCACTACTTGGCACTTGTGGGTAGGCACCTCCTCCCATTGGAGGAAAGCCACTAGGATAAGGATACTGACCAGAAGGGGGAAAAGATGACTCCTGACCTGCAGG;MAPQ=60;MATEID=4630563_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_75141501_75166501_289C;SPAN=3527;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:56 GQ:44.3 PL:[90.5, 0.0, 44.3] SR:31 DR:5 LR:-91.26 LO:91.26);ALT=T[chr10:75160561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75158143	+	chr10	75160561	+	.	12	6	4630566_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4630566_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_10_75141501_75166501_289C;SPAN=2418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:59 GQ:43.4 PL:[43.4, 0.0, 99.5] SR:6 DR:12 LR:-43.43 LO:44.65);ALT=G[chr10:75160561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75158173	+	chr10	75173768	+	.	76	0	4630725_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4630725_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:75158173(+)-10:75173768(-)__10_75166001_75191001D;SPAN=15595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:55 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:0 DR:76 LR:-224.5 LO:224.5);ALT=T[chr10:75173768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75632841	+	chr10	75634154	+	.	14	11	4631573_1	47.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4631573_2;MATENM=0;NM=1;NUMPARTS=4;REPSEQ=CCC;SCTG=c_10_75631501_75656501_217C;SPAN=1313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:44 GQ:47.6 PL:[47.6, 0.0, 57.5] SR:11 DR:14 LR:-47.5 LO:47.57);ALT=C[chr10:75634154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75898188	+	chr10	75910516	+	.	8	0	4632150_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4632150_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:75898188(+)-10:75910516(-)__10_75901001_75926001D;SPAN=12328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=T[chr10:75910516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75936635	+	chr10	75984295	+	.	10	0	4632299_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4632299_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:75936635(+)-10:75984295(-)__10_75974501_75999501D;SPAN=47660;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=C[chr10:75984295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75936644	+	chr10	75960520	+	.	28	18	4632105_1	95.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4632105_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_75950001_75975001_201C;SPAN=23876;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:28 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:18 DR:28 LR:-95.72 LO:95.72);ALT=G[chr10:75960520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	75936657	+	chr10	76074424	+	.	17	0	4632390_1	48.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4632390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:75936657(+)-10:76074424(-)__10_76072501_76097501D;SPAN=137767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:29 GQ:21.8 PL:[48.2, 0.0, 21.8] SR:0 DR:17 LR:-48.79 LO:48.79);ALT=C[chr10:76074424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	76430029	+	chr10	76468077	+	.	10	9	4632980_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4632980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_76464501_76489501_74C;SPAN=38048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:27 GQ:15.8 PL:[48.8, 0.0, 15.8] SR:9 DR:10 LR:-49.67 LO:49.67);ALT=T[chr10:76468077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	76598512	+	chr10	76602357	+	.	0	9	4633236_1	16.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=4633236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_76587001_76612001_129C;SPAN=3845;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:9 DR:0 LR:-16.16 LO:19.94);ALT=T[chr10:76602357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	76871515	+	chr10	76910269	+	.	13	0	4633752_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4633752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:76871515(+)-10:76910269(-)__10_76905501_76930501D;SPAN=38754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:39 GQ:32.3 PL:[32.3, 0.0, 62.0] SR:0 DR:13 LR:-32.35 LO:32.87);ALT=T[chr10:76910269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	77191514	+	chr10	77198152	+	.	0	24	4634296_1	63.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=4634296_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_77175001_77200001_103C;SPAN=6638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:57 GQ:63.8 PL:[63.8, 0.0, 73.7] SR:24 DR:0 LR:-63.78 LO:63.83);ALT=T[chr10:77198152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	77191566	+	chr10	77795763	+	.	30	0	4635012_1	88.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4635012_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:77191566(+)-10:77795763(-)__10_77787501_77812501D;SPAN=604197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:39 GQ:5.9 PL:[88.4, 0.0, 5.9] SR:0 DR:30 LR:-92.71 LO:92.71);ALT=A[chr10:77795763[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	77198254	+	chr10	77806922	+	CACTGGAAGGACTGAGCGCATTCAGGAGCCTGGAGGAACTCATCTTGGACAACAATCAGCTGGGGGACGACCTTGTGTTGCCAGGGTTACCCAGACTGCATACCTTAACCCTCAACAAGAACCGA	0	41	4634308_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AT;INSERTION=CACTGGAAGGACTGAGCGCATTCAGGAGCCTGGAGGAACTCATCTTGGACAACAATCAGCTGGGGGACGACCTTGTGTTGCCAGGGTTACCCAGACTGCATACCTTAACCCTCAACAAGAACCGA;MAPQ=60;MATEID=4634308_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_77175001_77200001_53C;SPAN=608668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:33 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:41 DR:0 LR:-118.8 LO:118.8);ALT=T[chr10:77806922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78255578	+	chr10	78261020	+	.	42	36	4635628_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCAGT;MAPQ=60;MATEID=4635628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_78253001_78278001_187C;SPAN=5442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:18 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:36 DR:42 LR:-178.2 LO:178.2);ALT=T[chr10:78261020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78346604	+	chr10	78351578	+	.	53	25	4636083_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAATACTTAATTT;MAPQ=60;MATEID=4636083_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_78351001_78376001_169C;SPAN=4974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:10 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:25 DR:53 LR:-184.8 LO:184.8);ALT=T[chr10:78351578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	78516976	+	chr14	51644864	+	.	4	9	4635937_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TATATATATGTGTGTATATATA;MAPQ=60;MATEID=4635937_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_10_78498001_78523001_203C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:17 GQ:8.6 PL:[31.7, 0.0, 8.6] SR:9 DR:4 LR:-32.36 LO:32.36);ALT=A[chr14:51644864[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	79184909	+	chr22	44376043	-	.	31	33	7319557_1	99.0	.	DISC_MAPQ=10;EVDNC=ASDIS;HOMSEQ=ATGGATGGATGGATGGATGGATGGATG;MAPQ=25;MATEID=7319557_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_44369501_44394501_144C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:86 GQ:52.7 PL:[155.0, 0.0, 52.7] SR:33 DR:31 LR:-157.6 LO:157.6);ALT=G]chr22:44376043];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr10	79793707	+	chr10	79795266	+	.	113	0	4638092_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4638092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:79793707(+)-10:79795266(-)__10_79772001_79797001D;SPAN=1559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:113 DP:146 GQ:20 PL:[333.5, 0.0, 20.0] SR:0 DR:113 LR:-349.9 LO:349.9);ALT=C[chr10:79795266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81107368	+	chr10	81109419	+	.	9	0	4640186_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4640186_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:81107368(+)-10:81109419(-)__10_81095001_81120001D;SPAN=2051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:0 DR:9 LR:-17.25 LO:20.3);ALT=C[chr10:81109419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81803484	+	chr10	81787670	+	.	15	10	4641564_1	65.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTGAGACAGAGTCTTGCTGTGTTGCCCAGGC;MAPQ=60;MATEID=4641564_2;MATENM=1;NM=5;NUMPARTS=2;SCTG=c_10_81781001_81806001_184C;SPAN=15814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:37 GQ:23 PL:[65.9, 0.0, 23.0] SR:10 DR:15 LR:-66.98 LO:66.98);ALT=]chr10:81803484]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	81915669	+	chr10	81917396	+	.	0	26	4641955_1	68.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4641955_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_81903501_81928501_290C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:66 GQ:68 PL:[68.0, 0.0, 91.1] SR:26 DR:0 LR:-67.95 LO:68.15);ALT=C[chr10:81917396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81929115	+	chr10	81930555	+	.	2	7	4641981_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4641981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_81928001_81953001_151C;SPAN=1440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:7 DR:2 LR:-9.932 LO:18.32);ALT=C[chr10:81930555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81930674	+	chr10	81965096	+	GTGCAGCTGGTGGGTAGCCACCTGGGGGCGGGGGATAGCCAGGGTAGCTCATGGTTAGATCTTTGACTCAGCAACTCCACTTCTGTAAGTCTCTTCCCCAGACACA	16	64	4642027_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CACCTG;INSERTION=GTGCAGCTGGTGGGTAGCCACCTGGGGGCGGGGGATAGCCAGGGTAGCTCATGGTTAGATCTTTGACTCAGCAACTCCACTTCTGTAAGTCTCTTCCCCAGACACA;MAPQ=60;MATEID=4642027_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_81952501_81977501_188C;SPAN=34422;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:29 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:64 DR:16 LR:-234.4 LO:234.4);ALT=G[chr10:81965096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81932629	+	chr10	81965099	+	.	0	15	4642029_1	40.0	.	EVDNC=ASSMB;HOMSEQ=CTGG;MAPQ=60;MATEID=4642029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_81952501_81977501_7C;SPAN=32470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:34 GQ:40.4 PL:[40.4, 0.0, 40.4] SR:15 DR:0 LR:-40.3 LO:40.31);ALT=G[chr10:81965099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	81935962	+	chr10	81965183	+	.	28	0	4642032_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4642032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:81935962(+)-10:81965183(-)__10_81952501_81977501D;SPAN=29221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:33 GQ:5.4 PL:[89.1, 5.4, 0.0] SR:0 DR:28 LR:-89.59 LO:89.59);ALT=C[chr10:81965183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	82295395	+	chr16	75503315	+	.	15	0	6252462_1	42.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=6252462_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:82295395(+)-16:75503315(-)__16_75484501_75509501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:10 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=G[chr16:75503315[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr10	83641806	+	chr10	83827666	+	ATTAT	5	6	4644547_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATTAT;MAPQ=60;MATEID=4644547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_83814501_83839501_13C;SPAN=185860;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:24 GQ:26.6 PL:[29.9, 0.0, 26.6] SR:6 DR:5 LR:-29.81 LO:29.81);ALT=T[chr10:83827666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	84127819	+	chr10	84130365	+	.	32	33	4645094_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TTTTC;MAPQ=60;MATEID=4645094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_84108501_84133501_213C;SPAN=2546;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:17 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:33 DR:32 LR:-161.7 LO:161.7);ALT=C[chr10:84130365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	92631814	+	chr10	92635778	+	.	8	0	4658040_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4658040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:92631814(+)-10:92635778(-)__10_92634501_92659501D;SPAN=3964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=C[chr10:92635778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	92631821	+	chr10	92635312	+	.	11	0	4658041_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4658041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:92631821(+)-10:92635312(-)__10_92634501_92659501D;SPAN=3491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=T[chr10:92635312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	92980593	+	chr10	92982445	+	.	19	6	4658638_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4658638_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_92977501_93002501_108C;SPAN=1852;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:63 GQ:55.7 PL:[55.7, 0.0, 95.3] SR:6 DR:19 LR:-55.55 LO:56.18);ALT=G[chr10:92982445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	93683848	+	chr10	93695411	+	.	2	2	4659497_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4659497_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_93663501_93688501_213C;SPAN=11563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:22 GQ:7.4 PL:[7.4, 0.0, 43.7] SR:2 DR:2 LR:-7.244 LO:8.88);ALT=G[chr10:93695411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	94134599	+	chr10	94137654	+	GTTGACTTATCTTTT	0	25	4660739_1	58.0	.	EVDNC=ASSMB;INSERTION=GTTGACTTATCTTTT;MAPQ=60;MATEID=4660739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_94129001_94154001_34C;SPAN=3055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:88 GQ:58.7 PL:[58.7, 0.0, 154.4] SR:25 DR:0 LR:-58.68 LO:61.08);ALT=A[chr10:94137654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	94608393	+	chr10	94653105	+	.	17	5	4661355_1	56.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4661355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_94594501_94619501_82C;SPAN=44712;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:15 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:5 DR:17 LR:-56.11 LO:56.11);ALT=T[chr10:94653105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	95545477	+	chr10	95546496	+	CCACCACATGGCACACAAAAGGGTG	0	53	4662977_1	99.0	.	EVDNC=ASSMB;INSERTION=CCACCACATGGCACACAAAAGGGTG;MAPQ=60;MATEID=4662977_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_10_95525501_95550501_86C;SPAN=1019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:18 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:53 DR:0 LR:-155.1 LO:155.1);ALT=A[chr10:95546496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	101492115	+	chr10	101499464	+	.	10	0	4672637_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4672637_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:101492115(+)-10:101499464(-)__10_101479001_101504001D;SPAN=7349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=C[chr10:101499464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	101492167	+	chr10	101496002	+	.	17	13	4672638_1	55.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4672638_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_101479001_101504001_92C;SPAN=3835;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:65 GQ:55.1 PL:[55.1, 0.0, 101.3] SR:13 DR:17 LR:-55.01 LO:55.8);ALT=G[chr10:101496002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	101496076	+	chr10	101502909	+	GCTGATCGGATTGAATTATGTTCTGGTTTATCAGAGGGGGGAACTACACCCAGCATG	0	23	4672646_1	60.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=GCTGATCGGATTGAATTATGTTCTGGTTTATCAGAGGGGGGAACTACACCCAGCATG;MAPQ=60;MATEID=4672646_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_101479001_101504001_4C;SPAN=6833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:57 GQ:60.5 PL:[60.5, 0.0, 77.0] SR:23 DR:0 LR:-60.48 LO:60.6);ALT=T[chr10:101502909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102040811	+	chr10	102045854	+	.	0	21	4673881_1	61.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4673881_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_102018001_102043001_34C;SPAN=5043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:28 GQ:5.6 PL:[61.7, 0.0, 5.6] SR:21 DR:0 LR:-64.39 LO:64.39);ALT=C[chr10:102045854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102040860	+	chr10	102046361	+	.	22	0	4673882_1	66.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4673882_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:102040860(+)-10:102046361(-)__10_102018001_102043001D;SPAN=5501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:23 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:22 LR:-66.02 LO:66.02);ALT=A[chr10:102046361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102286312	+	chr10	102289135	+	GGTTCACCCCAGTTCAACCTCAGGCCCGGCTGGTCCCAGCTATACCATGGATCTCTCTCATGCTGTGAGCGGTCAGGGAGCTTCGGGTAGTCGCCAT	5	71	4674318_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=GGTTCACCCCAGTTCAACCTCAGGCCCGGCTGGTCCCAGCTATACCATGGATCTCTCTCATGCTGTGAGCGGTCAGGGAGCTTCGGGTAGTCGCCAT;MAPQ=60;MATEID=4674318_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_102263001_102288001_65C;SPAN=2823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:34 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:71 DR:5 LR:-221.2 LO:221.2);ALT=C[chr10:102289135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102286832	+	chr10	102289135	+	.	3	32	4674319_1	99.0	.	DISC_MAPQ=38;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=4674319_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_10_102263001_102288001_65C;SPAN=2303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:46 GQ:10.7 PL:[99.8, 0.0, 10.7] SR:32 DR:3 LR:-103.8 LO:103.8);ALT=C[chr10:102289135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102741300	+	chr10	102743512	+	.	0	24	4675104_1	62.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4675104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_102728501_102753501_62C;SPAN=2212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:64 GQ:62 PL:[62.0, 0.0, 91.7] SR:24 DR:0 LR:-61.89 LO:62.24);ALT=T[chr10:102743512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102792239	+	chr10	102794449	+	.	9	2	4675207_1	18.0	.	DISC_MAPQ=55;EVDNC=ASDIS;MAPQ=60;MATEID=4675207_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_102777501_102802501_262C;SPAN=2210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:2 DR:9 LR:-18.65 LO:22.38);ALT=C[chr10:102794449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	102792288	+	chr10	102795250	+	.	8	0	4675208_1	13.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4675208_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:102792288(+)-10:102795250(-)__10_102777501_102802501D;SPAN=2962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=A[chr10:102795250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	103912287	+	chr10	103916946	+	ACACAGCAGGATGCCAATGCCTCTTCCCTCTTAGACATCTATAGCTTCTGGCTCAA	10	15	4677264_1	46.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=ACACAGCAGGATGCCAATGCCTCTTCCCTCTTAGACATCTATAGCTTCTGGCTCAA;MAPQ=60;MATEID=4677264_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_103904501_103929501_225C;SPAN=4659;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:62 GQ:46.1 PL:[46.1, 0.0, 102.2] SR:15 DR:10 LR:-45.92 LO:47.18);ALT=T[chr10:103916946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21903372	+	chr10	104027094	+	.	5	22	6562716_1	69.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=TCTACTAAAAATACAAAAATTAGC;MAPQ=39;MATEID=6562716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21903001_21928001_274C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:8 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:22 DR:5 LR:-69.32 LO:69.32);ALT=]chr18:21903372]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	104184552	+	chr10	104192283	+	AGGTCGGCCTCCGGGAGGTGTGTCTGGACAAAGGCAAGGAGGGCTGCACTGACGATCCTCTCCAGCTCCATGCTCTCTCTT	66	32	4677795_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=AGGTCGGCCTCCGGGAGGTGTGTCTGGACAAAGGCAAGGAGGGCTGCACTGACGATCCTCTCCAGCTCCATGCTCTCTCTT;MAPQ=60;MATEID=4677795_2;MATENM=0;NM=88;NUMPARTS=3;SCTG=c_10_104174001_104199001_158C;SPAN=7731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:71 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:32 DR:66 LR:-227.8 LO:227.8);ALT=G[chr10:104192283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104184958	+	chr10	104192283	+	.	9	7	4677796_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=4677796_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_104174001_104199001_158C;SPAN=7325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:66 GQ:25.1 PL:[25.1, 0.0, 134.0] SR:7 DR:9 LR:-25.03 LO:29.37);ALT=G[chr10:104192283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104248895	+	chr10	104262356	+	TAGTTTGGAAAGCAGTATTTGGGGATCTGATCACCAGCAAAACCAGCTTTAATCACACCGGATC	13	15	4678203_1	59.0	.	DISC_MAPQ=50;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TAGTTTGGAAAGCAGTATTTGGGGATCTGATCACCAGCAAAACCAGCTTTAATCACACCGGATC;MAPQ=60;MATEID=4678203_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_104247501_104272501_110C;SPAN=13461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:63 GQ:59 PL:[59.0, 0.0, 92.0] SR:15 DR:13 LR:-58.86 LO:59.3);ALT=A[chr10:104262356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104250370	+	chr10	104262356	+	.	7	6	4678207_1	12.0	.	DISC_MAPQ=12;EVDNC=TSI_L;HOMSEQ=C;MAPQ=56;MATEID=4678207_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_10_104247501_104272501_110C;SPAN=11986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:52 GQ:12.5 PL:[12.5, 0.0, 111.5] SR:6 DR:7 LR:-12.32 LO:17.12);ALT=C[chr10:104262356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104459249	+	chr10	104465102	+	.	4	4	4678693_1	3.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4678693_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_104443501_104468501_146C;SPAN=5853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:60 GQ:3.5 PL:[3.5, 0.0, 142.1] SR:4 DR:4 LR:-3.551 LO:11.63);ALT=G[chr10:104465102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104614120	+	chr10	104620085	+	.	26	0	4678778_1	82.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4678778_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:104614120(+)-10:104620085(-)__10_104615001_104640001D;SPAN=5965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:0 DR:26 LR:-82.52 LO:82.52);ALT=C[chr10:104620085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104614184	+	chr10	104622630	+	CTGCTAGGTCAGGCAGCTCGAAACATGGTACTCCAGGAAGATGCCATCTTGCACTCAGAAGATAGTTTAAGGAAGATGGCAATAATAACAACACATCTTCAATACCAGCAAGAAGCTATTCAGAAGAA	0	29	4678780_1	85.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTGCTAGGTCAGGCAGCTCGAAACATGGTACTCCAGGAAGATGCCATCTTGCACTCAGAAGATAGTTTAAGGAAGATGGCAATAATAACAACACATCTTCAATACCAGCAAGAAGCTATTCAGAAGAA;MAPQ=60;MATEID=4678780_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_104615001_104640001_136C;SPAN=8446;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:25 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:29 DR:0 LR:-85.82 LO:85.82);ALT=G[chr10:104622630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104899237	+	chr10	104934614	+	.	4	4	4679511_1	16.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4679511_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_104933501_104958501_110C;SPAN=35377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:26 GQ:16.1 PL:[16.1, 0.0, 45.8] SR:4 DR:4 LR:-16.06 LO:16.91);ALT=C[chr10:104934614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	104934740	+	chr10	104940942	+	.	0	9	4679515_1	11.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4679515_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_104933501_104958501_63C;SPAN=6202;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:9 DR:0 LR:-11.56 LO:18.68);ALT=C[chr10:104940942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105148933	+	chr10	105156165	+	.	16	0	4679883_1	29.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=4679883_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:105148933(+)-10:105156165(-)__10_105154001_105179001D;SPAN=7232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:85 GQ:29.9 PL:[29.9, 0.0, 175.1] SR:0 DR:16 LR:-29.79 LO:35.79);ALT=A[chr10:105156165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105152063	+	chr10	105156165	+	.	55	0	4679884_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=4679884_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:105152063(+)-10:105156165(-)__10_105154001_105179001D;SPAN=4102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:85 GQ:46.4 PL:[158.6, 0.0, 46.4] SR:0 DR:55 LR:-161.8 LO:161.8);ALT=A[chr10:105156165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105156166	-	chrX	73393696	+	.	119	6	7450102_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GGAATTTGCGGCTTTGGCAG;MAPQ=60;MATEID=7450102_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_23_73377501_73402501_55C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:41 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:6 DR:119 LR:-359.8 LO:359.8);ALT=[chrX:73393696[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr10	105642599	+	chr10	105648830	+	.	3	14	4681005_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4681005_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_105619501_105644501_84C;SPAN=6231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:33 GQ:30.8 PL:[47.3, 0.0, 30.8] SR:14 DR:3 LR:-47.31 LO:47.31);ALT=T[chr10:105648830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105664916	+	chr10	105670285	+	.	0	13	4680918_1	34.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4680918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_105644001_105669001_15C;SPAN=5369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:32 GQ:34.4 PL:[34.4, 0.0, 41.0] SR:13 DR:0 LR:-34.24 LO:34.3);ALT=T[chr10:105670285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105670382	+	chr10	105677218	+	.	0	22	4680932_1	56.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4680932_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_105668501_105693501_230C;SPAN=6836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:60 GQ:56.3 PL:[56.3, 0.0, 89.3] SR:22 DR:0 LR:-56.37 LO:56.77);ALT=T[chr10:105677218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	105670429	+	chr10	105677857	+	.	10	0	4680933_1	16.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4680933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:105670429(+)-10:105677857(-)__10_105668501_105693501D;SPAN=7428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:0 DR:10 LR:-16.21 LO:21.62);ALT=T[chr10:105677857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	106014721	+	chr10	106019330	+	AAGCGCGCCCCCGGGGCCGGTCCCGGAGGGCTCGATCCGCATCTACAGCATGAGGTTCTGCCCGTTTGCTGAGAGGACGCGTCTAGTCCTGAAGGCCAAGGGAA	18	70	4681479_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TCAGG;INSERTION=AAGCGCGCCCCCGGGGCCGGTCCCGGAGGGCTCGATCCGCATCTACAGCATGAGGTTCTGCCCGTTTGCTGAGAGGACGCGTCTAGTCCTGAAGGCCAAGGGAA;MAPQ=60;MATEID=4681479_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_106011501_106036501_111C;SPAN=4609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:87 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:70 DR:18 LR:-257.5 LO:257.5);ALT=G[chr10:106019330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	106015030	+	chr10	106019330	+	.	83	58	4681482_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=TCAGG;MAPQ=60;MATEID=4681482_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_10_106011501_106036501_111C;SPAN=4300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:82 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:58 DR:83 LR:-356.5 LO:356.5);ALT=G[chr10:106019330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	106019558	+	chr10	106025840	+	GCCATCCTTGGTAGGAAGCTTTATTAGAAGCCAAAATAAAGAAGACTATGATGGCCTAAAAGAAGAATTTCGTAAAGAATTTACCAAGCTAGAGG	9	35	4681497_1	99.0	.	DISC_MAPQ=22;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=GCCATCCTTGGTAGGAAGCTTTATTAGAAGCCAAAATAAAGAAGACTATGATGGCCTAAAAGAAGAATTTCGTAAAGAATTTACCAAGCTAGAGG;MAPQ=51;MATEID=4681497_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_106011501_106036501_112C;SPAN=6282;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:56 GQ:21.2 PL:[113.6, 0.0, 21.2] SR:35 DR:9 LR:-117.0 LO:117.0);ALT=T[chr10:106025840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	106019558	+	chr10	106022735	+	.	11	10	4681496_1	36.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4681496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_106011501_106036501_267C;SPAN=3177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:59 GQ:36.8 PL:[36.8, 0.0, 106.1] SR:10 DR:11 LR:-36.83 LO:38.71);ALT=T[chr10:106022735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	106022833	+	chr10	106025840	+	.	0	21	4681501_1	53.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4681501_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_106011501_106036501_47C;SPAN=3007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:60 GQ:53 PL:[53.0, 0.0, 92.6] SR:21 DR:0 LR:-53.07 LO:53.65);ALT=G[chr10:106025840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46237807	+	chr10	126145906	+	.	5	19	4712002_1	59.0	.	DISC_MAPQ=21;EVDNC=ASDIS;HOMSEQ=CTCTCTCTCTCTCTCTCTCTCTTTCTTTCTTT;MAPQ=16;MATEID=4712002_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_10_126126001_126151001_199C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:6 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:19 DR:5 LR:-59.41 LO:59.41);ALT=]chr13:46237807]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr10	126150556	+	chr10	126172705	+	.	31	11	4712009_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4712009_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_126126001_126151001_159C;SPAN=22149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:34 DP:21 GQ:9 PL:[99.0, 9.0, 0.0] SR:11 DR:31 LR:-99.02 LO:99.02);ALT=G[chr10:126172705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	126477727	+	chr10	126480293	+	AGATTTCACCTGTATCTCCATATTCTCGGAAAGTTTGCAGTTCTCTCTCATAGACAGCATCCCAA	11	22	4712487_1	64.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGATTTCACCTGTATCTCCATATTCTCGGAAAGTTTGCAGTTCTCTCTCATAGACAGCATCCCAA;MAPQ=60;MATEID=4712487_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_126469001_126494001_163C;SPAN=2566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:66 GQ:64.7 PL:[64.7, 0.0, 94.4] SR:22 DR:11 LR:-64.64 LO:64.97);ALT=C[chr10:126480293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	126478943	+	chr10	126480356	+	.	15	0	4712494_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4712494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:126478943(+)-10:126480356(-)__10_126469001_126494001D;SPAN=1413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:52 GQ:35.6 PL:[35.6, 0.0, 88.4] SR:0 DR:15 LR:-35.43 LO:36.77);ALT=A[chr10:126480356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127190418	-	chr10	127201102	+	.	7	54	4713844_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=4713844_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ACAC;SCTG=c_10_127179501_127204501_72C;SPAN=10684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:84 GQ:26.9 PL:[175.4, 0.0, 26.9] SR:54 DR:7 LR:-181.3 LO:181.3);ALT=[chr10:127201102[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	127201222	+	chr10	127190797	+	.	24	32	4713846_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CCACCAT;MAPQ=60;MATEID=4713846_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_10_127179501_127204501_72C;SPAN=10425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:69 GQ:7.7 PL:[159.5, 0.0, 7.7] SR:32 DR:24 LR:-167.8 LO:167.8);ALT=]chr10:127201222]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	127191657	+	chr10	127197235	+	.	81	55	4713856_1	99.0	.	DISC_MAPQ=32;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=4713856_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127179501_127204501_169C;SPAN=5578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:47 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:55 DR:81 LR:-323.5 LO:323.5);ALT=C[chr10:127197235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127408485	+	chr10	127409771	+	.	3	4	4714236_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4714236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127400001_127425001_221C;SPAN=1286;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:60 GQ:3.5 PL:[3.5, 0.0, 142.1] SR:4 DR:3 LR:-3.551 LO:11.63);ALT=G[chr10:127409771[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127477576	+	chr10	127483449	+	.	2	2	4714189_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4714189_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127473501_127498501_4C;SPAN=5873;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:65 GQ:4.2 PL:[0.0, 4.2, 165.0] SR:2 DR:2 LR:4.406 LO:6.878);ALT=T[chr10:127483449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127503701	+	chr10	127504746	+	.	0	6	4714264_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4714264_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127498001_127523001_136C;SPAN=1045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:60 GQ:3.5 PL:[3.5, 0.0, 142.1] SR:6 DR:0 LR:-3.551 LO:11.63);ALT=T[chr10:127504746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127505096	+	chr10	127511598	+	.	0	42	4714267_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4714267_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_127498001_127523001_268C;SPAN=6502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:70 GQ:50.3 PL:[119.6, 0.0, 50.3] SR:42 DR:0 LR:-121.2 LO:121.2);ALT=T[chr10:127511598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127512292	+	chr10	127516125	+	AAGTGAATATTGAATTTGAAGCTTATTCCCTATCAGATAATGATTATGACGGAATTAAGAAATTACTGCAGC	10	31	4714283_1	95.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAGTGAATATTGAATTTGAAGCTTATTCCCTATCAGATAATGATTATGACGGAATTAAGAAATTACTGCAGC;MAPQ=60;MATEID=4714283_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_127498001_127523001_161C;SPAN=3833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:64 GQ:58.7 PL:[95.0, 0.0, 58.7] SR:31 DR:10 LR:-95.3 LO:95.3);ALT=G[chr10:127516125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	127512292	+	chr10	127515158	+	.	20	18	4714282_1	74.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=4714282_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_10_127498001_127523001_161C;SPAN=2866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:68 GQ:74 PL:[74.0, 0.0, 90.5] SR:18 DR:20 LR:-74.01 LO:74.1);ALT=G[chr10:127515158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	129060203	+	chr10	129058857	+	.	34	0	4716743_1	93.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=4716743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:129058857(-)-10:129060203(+)__10_129041501_129066501D;SPAN=1346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:69 GQ:73.7 PL:[93.5, 0.0, 73.7] SR:0 DR:34 LR:-93.66 LO:93.66);ALT=]chr10:129060203]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	129846101	+	chr10	129847792	+	.	0	9	4717903_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4717903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_129825501_129850501_25C;SPAN=1691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:9 DR:0 LR:-9.661 LO:18.26);ALT=G[chr10:129847792[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131265562	+	chr10	131334504	+	.	63	9	4720138_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=4720138_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_131320001_131345001_266C;SPAN=68942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:31 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:9 DR:63 LR:-201.3 LO:201.3);ALT=T[chr10:131334504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131265562	+	chr10	131557464	+	ACTTGGAAAAATGGACAAGGATTGTGAAATGAAACGCACCACACTGGACAGCCCTTTGGGGAAGCTGGAGCTGTCTGGTTGTGAGCAGGGTCTGCACGAAATAAAGCTCCTGGGCAAGGGGACGTCTGCAGCTGATGCCGTGGAGGTCCCAGCCCCCGCTGCGGTTCTCGGAGGTCCGGAGCCCCTGATGCAGTGCACAGCCTGGCTGAATGCCTATTTCCACCAGCCCGAGGCTATCGAAGAGTTCCCCGTGCCGGCTCTTCACCATCCCGTTTTCCAGCA	2	19	4719938_1	59.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACTTGGAAAAATGGACAAGGATTGTGAAATGAAACGCACCACACTGGACAGCCCTTTGGGGAAGCTGGAGCTGTCTGGTTGTGAGCAGGGTCTGCACGAAATAAAGCTCCTGGGCAAGGGGACGTCTGCAGCTGATGCCGTGGAGGTCCCAGCCCCCGCTGCGGTTCTCGGAGGTCCGGAGCCCCTGATGCAGTGCACAGCCTGGCTGAATGCCTATTTCCACCAGCCCGAGGCTATCGAAGAGTTCCCCGTGCCGGCTCTTCACCATCCCGTTTTCCAGCA;MAPQ=60;MATEID=4719938_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_131246501_131271501_225C;SPAN=291902;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:36 GQ:26.6 PL:[59.6, 0.0, 26.6] SR:19 DR:2 LR:-60.19 LO:60.19);ALT=T[chr10:131557464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131265613	+	chr10	131506157	+	.	60	0	4719939_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4719939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:131265613(+)-10:131506157(-)__10_131246501_131271501D;SPAN=240544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:25 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:60 LR:-178.2 LO:178.2);ALT=A[chr10:131506157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131334641	+	chr10	131506159	+	.	4	77	4720298_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=4720298_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_10_131491501_131516501_52C;SPAN=171518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:53 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:77 DR:4 LR:-237.7 LO:237.7);ALT=A[chr10:131506159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131557607	+	chr10	131565052	+	.	4	19	4720443_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=4720443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_131540501_131565501_166C;SPAN=7445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:60 GQ:53 PL:[53.0, 0.0, 92.6] SR:19 DR:4 LR:-53.07 LO:53.65);ALT=T[chr10:131565052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	131934756	+	chr10	131943474	+	.	10	0	4721041_1	22.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4721041_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:131934756(+)-10:131943474(-)__10_131932501_131957501D;SPAN=8718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:40 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-22.17 LO:23.78);ALT=G[chr10:131943474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	132840299	+	chr10	132841347	+	.	16	3	4722507_1	56.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GGGGTAAGATAGGGTATGGGGGGTGGGGTAAGATAGGGTATCGGG;MAPQ=60;MATEID=4722507_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GGG;SCTG=c_10_132839001_132864001_202C;SECONDARY;SPAN=1048;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:10 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:3 DR:16 LR:-56.11 LO:56.11);ALT=G[chr10:132841347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	132909062	+	chr10	132912780	+	.	48	33	4722583_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTCA;MAPQ=60;MATEID=4722583_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_132912501_132937501_31C;SPAN=3718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:11 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:33 DR:48 LR:-204.7 LO:204.7);ALT=A[chr10:132912780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	13023198	+	chr18	53590863	-	.	40	48	4764331_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CATTAGATTCTCATAAGGAGCATGCAGCCTAG;MAPQ=60;MATEID=4764331_2;MATENM=2;NM=1;NUMPARTS=2;SCTG=c_11_13009501_13034501_28C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:24 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:48 DR:40 LR:-241.0 LO:241.0);ALT=G]chr18:53590863];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	13565922	+	chr20	37970249	+	.	8	46	4765729_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCTGCCTCAGCCTCCCAAGTAGATGG;MAPQ=60;MATEID=4765729_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_13548501_13573501_234C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:11 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:46 DR:8 LR:-141.9 LO:141.9);ALT=G[chr20:37970249[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr20	37970324	+	chr11	13566291	+	.	7	17	7006922_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GCCACCATGCCTGGCTAATTTTTGTATTTTTAGTAG;MAPQ=60;MATEID=7006922_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCACCA;SCTG=c_20_37950501_37975501_188C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:55 GQ:47.7 PL:[47.7, 0.0, 50.3] SR:17 DR:7 LR:-47.55 LO:47.56);ALT=]chr20:37970324]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	14501261	+	chr11	14502305	+	.	2	4	4768172_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4768172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14479501_14504501_95C;SPAN=1044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:75 GQ:0.3 PL:[0.0, 0.3, 181.5] SR:4 DR:2 LR:0.5133 LO:11.02);ALT=C[chr11:14502305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14526796	+	chr11	14529202	+	.	3	12	4768312_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4768312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14504001_14529001_224C;SPAN=2406;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:46 GQ:37.1 PL:[37.1, 0.0, 73.4] SR:12 DR:3 LR:-37.05 LO:37.75);ALT=T[chr11:14529202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14529314	+	chr11	14532418	+	.	2	10	4768399_1	18.0	.	DISC_MAPQ=14;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4768399_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14528501_14553501_192C;SPAN=3104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:78 GQ:18.5 PL:[18.5, 0.0, 170.3] SR:10 DR:2 LR:-18.48 LO:25.68);ALT=T[chr11:14532418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14532497	+	chr11	14535112	+	.	2	4	4768411_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TTAC;MAPQ=60;MATEID=4768411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14528501_14553501_196C;SPAN=2615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:75 GQ:0.3 PL:[0.0, 0.3, 181.5] SR:4 DR:2 LR:0.5133 LO:11.02);ALT=C[chr11:14535112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14535462	+	chr11	14539187	+	.	8	0	4768423_1	4.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4768423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:14535462(+)-11:14539187(-)__11_14528501_14553501D;SPAN=3725;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=C[chr11:14539187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14536038	+	chr11	14539188	+	.	3	43	4768424_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4768424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14528501_14553501_333C;SPAN=3150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:92 GQ:94.1 PL:[127.1, 0.0, 94.1] SR:43 DR:3 LR:-127.1 LO:127.1);ALT=C[chr11:14539188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14536082	+	chr11	14541842	+	.	16	0	4768425_1	18.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4768425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:14536082(+)-11:14541842(-)__11_14528501_14553501D;SPAN=5760;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:127 GQ:18.5 PL:[18.5, 0.0, 289.1] SR:0 DR:16 LR:-18.41 LO:32.73);ALT=A[chr11:14541842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14539330	+	chr11	14541841	+	.	82	0	4768435_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4768435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:14539330(+)-11:14541841(-)__11_14528501_14553501D;SPAN=2511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:116 GQ:41.3 PL:[239.3, 0.0, 41.3] SR:0 DR:82 LR:-247.1 LO:247.1);ALT=A[chr11:14541841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14540641	+	chr11	14541840	+	.	17	0	4768444_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4768444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:14540641(+)-11:14541840(-)__11_14528501_14553501D;SPAN=1199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:123 GQ:23 PL:[23.0, 0.0, 273.8] SR:0 DR:17 LR:-22.79 LO:35.52);ALT=C[chr11:14541840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	14632698	+	chr11	14664998	+	.	0	7	4768743_1	14.0	.	EVDNC=ASSMB;HOMSEQ=TACC;MAPQ=60;MATEID=4768743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_14651001_14676001_35C;SPAN=32300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:34 GQ:14 PL:[14.0, 0.0, 66.8] SR:7 DR:0 LR:-13.9 LO:15.96);ALT=C[chr11:14664998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	22844680	+	chr11	22851240	+	CTAAGTCCACCTTCTGGTGGGGGCCCGGATGTAGCAATTTGTTTTTCTATTTTTTCCTTTTTCTTTCTCTTTTCTTGCACAGATTGAACATCTAAAATTCCCCGAGATGCAGCCTCTTTTTGTCTTCTCTCTGCAGCCTCTGCAAGCTTTGCTCTTTTCTCTT	0	34	4790228_1	85.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CTAAGTCCACCTTCTGGTGGGGGCCCGGATGTAGCAATTTGTTTTTCTATTTTTTCCTTTTTCTTTCTCTTTTCTTGCACAGATTGAACATCTAAAATTCCCCGAGATGCAGCCTCTTTTTGTCTTCTCTCTGCAGCCTCTGCAAGCTTTGCTCTTTTCTCTT;MAPQ=60;MATEID=4790228_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_22834001_22859001_165C;SPAN=6560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:100 GQ:85.1 PL:[85.1, 0.0, 157.7] SR:34 DR:0 LR:-85.14 LO:86.33);ALT=C[chr11:22851240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	22844680	+	chr11	22848753	+	.	3	17	4790227_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4790227_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_22834001_22859001_165C;SPAN=4073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:81 GQ:44.3 PL:[44.3, 0.0, 149.9] SR:17 DR:3 LR:-44.08 LO:47.43);ALT=C[chr11:22848753[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	22848934	+	chr11	22851256	+	.	31	0	4790244_1	74.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4790244_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:22848934(+)-11:22851256(-)__11_22834001_22859001D;SPAN=2322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:102 GQ:74.9 PL:[74.9, 0.0, 170.6] SR:0 DR:31 LR:-74.7 LO:76.84);ALT=T[chr11:22851256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	22849421	+	chr11	22851240	+	.	13	15	4790247_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=4790247_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_11_22834001_22859001_165C;SPAN=1819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:106 GQ:37.4 PL:[37.4, 0.0, 218.9] SR:15 DR:13 LR:-37.3 LO:44.76);ALT=C[chr11:22851240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	23205525	+	chr11	23211205	+	.	8	0	4791011_1	12.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=4791011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:23205525(+)-11:23211205(-)__11_23201501_23226501D;SPAN=5680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=G[chr11:23211205[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32605476	+	chr11	32608555	+	.	70	18	4813771_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4813771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_32585001_32610001_63C;SPAN=3079;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:95 GQ:0.8 PL:[228.5, 0.0, 0.8] SR:18 DR:70 LR:-242.1 LO:242.1);ALT=G[chr11:32608555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32605482	+	chr11	32610136	+	.	52	0	4813773_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4813773_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:32605482(+)-11:32610136(-)__11_32585001_32610001D;SPAN=4654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:47 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=T[chr11:32610136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32608690	+	chr11	32610138	+	.	0	104	4813782_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4813782_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_32585001_32610001_160C;SPAN=1448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:65 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:104 DR:0 LR:-307.0 LO:307.0);ALT=G[chr11:32610138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32611187	+	chr11	32615410	+	.	2	17	4813585_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=4813585_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_11_32609501_32634501_346C;SPAN=4223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:74 GQ:36.2 PL:[36.2, 0.0, 141.8] SR:17 DR:2 LR:-36.07 LO:39.69);ALT=G[chr11:32615410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32611187	+	chr11	32616458	+	TGATGCTGCTTCAAAAGTCATGGTGGAATTGCTCGGAAGTTACACAGAGGACAATGCTTCCCAGGCTCGAGTTGATGCCCAC	7	30	4813586_1	88.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=TGATGCTGCTTCAAAAGTCATGGTGGAATTGCTCGGAAGTTACACAGAGGACAATGCTTCCCAGGCTCGAGTTGATGCCCAC;MAPQ=60;MATEID=4813586_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_32609501_32634501_346C;SPAN=5271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:76 GQ:88.4 PL:[88.4, 0.0, 95.0] SR:30 DR:7 LR:-88.34 LO:88.36);ALT=G[chr11:32616458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32617594	+	chr11	32623823	+	CCTGTTACATGAACAGAATATGGCAAAAATGAGACTACTTACTTTTATGGGAATGGCAGTAGAAAATAAGGAAATTTCTTTTGACACAATGCAGCAAGAACTTCAGATTGGAGCTGATGATGTTGAAGCATTTGTTATTGACGCCGTAAGAACTAAAATGGTCTACTGCAAAATTGATCAGACCCAGAGAAAAGTAGTTGTC	0	142	4813602_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCTGTTACATGAACAGAATATGGCAAAAATGAGACTACTTACTTTTATGGGAATGGCAGTAGAAAATAAGGAAATTTCTTTTGACACAATGCAGCAAGAACTTCAGATTGGAGCTGATGATGTTGAAGCATTTGTTATTGACGCCGTAAGAACTAAAATGGTCTACTGCAAAATTGATCAGACCCAGAGAAAAGTAGTTGTC;MAPQ=60;MATEID=4813602_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_32609501_32634501_330C;SPAN=6229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:142 DP:126 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:142 DR:0 LR:-419.2 LO:419.2);ALT=G[chr11:32623823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	32617594	+	chr11	32622234	+	.	9	11	4813601_1	41.0	.	DISC_MAPQ=51;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4813601_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_11_32609501_32634501_330C;SPAN=4640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:90 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:11 DR:9 LR:-41.64 LO:46.37);ALT=G[chr11:32622234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	33163535	+	chr11	33182844	+	.	27	12	4815475_1	96.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4815475_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_33148501_33173501_67C;SPAN=19309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:47 GQ:17 PL:[96.2, 0.0, 17.0] SR:12 DR:27 LR:-99.25 LO:99.25);ALT=G[chr11:33182844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	33731890	+	chr11	33738915	+	.	0	15	4817285_1	32.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=4817285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_33736501_33761501_127C;SPAN=7025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:15 DR:0 LR:-32.72 LO:35.42);ALT=C[chr11:33738915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	33731925	+	chr11	33757925	+	.	8	0	4817286_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4817286_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:33731925(+)-11:33757925(-)__11_33736501_33761501D;SPAN=26000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:0 DR:8 LR:-10.97 LO:16.77);ALT=T[chr11:33757925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	33739019	+	chr11	33743923	+	.	0	8	4817300_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4817300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_33736501_33761501_2C;SPAN=4904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:8 DR:0 LR:2.039 LO:14.52);ALT=T[chr11:33743923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	33739065	+	chr11	33757925	+	.	16	0	4817301_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4817301_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:33739065(+)-11:33757925(-)__11_33736501_33761501D;SPAN=18860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:112 GQ:22.7 PL:[22.7, 0.0, 247.1] SR:0 DR:16 LR:-22.47 LO:33.68);ALT=T[chr11:33757925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34127339	+	chr11	34129756	+	.	2	2	4818771_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4818771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34104001_34129001_307C;SPAN=2417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:60 GQ:3 PL:[0.0, 3.0, 151.8] SR:2 DR:2 LR:3.051 LO:7.022);ALT=G[chr11:34129756[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34460626	+	chr11	34470737	+	.	111	48	4819533_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4819533_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_34447001_34472001_46C;SPAN=10111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:124 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:48 DR:111 LR:-399.4 LO:399.4);ALT=G[chr11:34470737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34460627	+	chr11	34472533	+	.	20	4	4819534_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4819534_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34447001_34472001_359C;SPAN=11906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:50 GQ:59 PL:[62.3, 0.0, 59.0] SR:4 DR:20 LR:-62.38 LO:62.38);ALT=G[chr11:34472533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34470911	+	chr11	34472533	+	.	7	23	4819738_1	76.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4819738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_162C;SPAN=1622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:59 GQ:66.5 PL:[76.4, 0.0, 66.5] SR:23 DR:7 LR:-76.48 LO:76.48);ALT=G[chr11:34472533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34473805	+	chr11	34475344	+	.	9	0	4819743_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4819743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:34473805(+)-11:34475344(-)__11_34471501_34496501D;SPAN=1539;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-7.764 LO:17.89);ALT=A[chr11:34475344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34475473	+	chr11	34477556	+	.	18	10	4819752_1	50.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4819752_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_24C;SPAN=2083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:83 GQ:50.3 PL:[50.3, 0.0, 149.3] SR:10 DR:18 LR:-50.14 LO:52.96);ALT=G[chr11:34477556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34478365	+	chr11	34482795	+	.	13	22	4819762_1	67.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4819762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_335C;SPAN=4430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:116 GQ:67.7 PL:[67.7, 0.0, 212.9] SR:22 DR:13 LR:-67.6 LO:71.85);ALT=G[chr11:34482795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34478415	+	chr11	34485650	+	.	12	0	4819763_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4819763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:34478415(+)-11:34485650(-)__11_34471501_34496501D;SPAN=7235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:105 GQ:11.3 PL:[11.3, 0.0, 242.3] SR:0 DR:12 LR:-11.17 LO:24.01);ALT=C[chr11:34485650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34482938	+	chr11	34485651	+	.	25	14	4819780_1	77.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4819780_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_250C;SPAN=2713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:115 GQ:77.9 PL:[77.9, 0.0, 200.0] SR:14 DR:25 LR:-77.78 LO:80.8);ALT=T[chr11:34485651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34485784	+	chr11	34489832	+	.	9	29	4819791_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=4819791_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_240C;SPAN=4048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:123 GQ:89 PL:[89.0, 0.0, 207.8] SR:29 DR:9 LR:-88.81 LO:91.51);ALT=T[chr11:34489832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34489944	+	chr11	34492504	+	.	6	18	4819802_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=4819802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_34471501_34496501_141C;SPAN=2560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:92 GQ:47.9 PL:[47.9, 0.0, 173.3] SR:18 DR:6 LR:-47.7 LO:51.81);ALT=T[chr11:34492504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	34489984	+	chr11	34492911	+	.	26	0	4819803_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4819803_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:34489984(+)-11:34492911(-)__11_34471501_34496501D;SPAN=2927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:102 GQ:58.4 PL:[58.4, 0.0, 187.1] SR:0 DR:26 LR:-58.19 LO:62.08);ALT=G[chr11:34492911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35160917	+	chr11	35198121	+	.	59	53	4821704_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4821704_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35157501_35182501_184C;SPAN=37204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:112 DP:201 GQ:99 PL:[315.5, 0.0, 170.3] SR:53 DR:59 LR:-317.5 LO:317.5);ALT=G[chr11:35198121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35201954	+	chr11	35208377	+	.	2	6	4822001_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4822001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35206501_35231501_150C;SPAN=6423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:38 GQ:12.8 PL:[12.8, 0.0, 78.8] SR:6 DR:2 LR:-12.81 LO:15.58);ALT=G[chr11:35208377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35208447	+	chr11	35211382	+	.	4	26	4822008_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4822008_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35206501_35231501_149C;SPAN=2935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:108 GQ:59.9 PL:[59.9, 0.0, 201.8] SR:26 DR:4 LR:-59.87 LO:64.2);ALT=A[chr11:35211382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35240934	+	chr11	35243197	+	.	0	14	4821646_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=4821646_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35231001_35256001_71C;SPAN=2263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:86 GQ:23 PL:[23.0, 0.0, 184.7] SR:14 DR:0 LR:-22.91 LO:30.33);ALT=G[chr11:35243197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35243281	+	chr11	35250674	+	.	0	7	4821656_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=4821656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_35231001_35256001_311C;SPAN=7393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:88 GQ:0.6 PL:[0.0, 0.6, 214.5] SR:7 DR:0 LR:0.7344 LO:12.84);ALT=T[chr11:35250674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	35720740	+	chr11	35729094	-	.	13	0	4823159_1	37.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4823159_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:35720740(+)-11:35729094(+)__11_35721001_35746001D;SPAN=8354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:21 GQ:11 PL:[37.4, 0.0, 11.0] SR:0 DR:13 LR:-37.82 LO:37.82);ALT=G]chr11:35729094];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	36300213	+	chr11	36310910	+	.	33	0	4824914_1	95.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4824914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:36300213(+)-11:36310910(-)__11_36309001_36334001D;SPAN=10697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:52 GQ:29 PL:[95.0, 0.0, 29.0] SR:0 DR:33 LR:-96.6 LO:96.6);ALT=C[chr11:36310910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	36302389	+	chr11	36310911	+	.	19	4	4824916_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4824916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_36309001_36334001_243C;SPAN=8522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:54 GQ:48.2 PL:[48.2, 0.0, 81.2] SR:4 DR:19 LR:-48.09 LO:48.6);ALT=T[chr11:36310911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	36616142	+	chr11	36631629	+	.	16	2	4825591_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4825591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_36627501_36652501_41C;SPAN=15487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:43 GQ:41.3 PL:[41.3, 0.0, 61.1] SR:2 DR:16 LR:-41.17 LO:41.42);ALT=G[chr11:36631629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	9239910	+	chr11	37130845	+	.	5	9	6102834_1	23.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGAGAGAGAGAGAGAGAGAGAGAGAGA;MAPQ=60;MATEID=6102834_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_9236501_9261501_171C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:60 GQ:23.3 PL:[23.3, 0.0, 122.3] SR:9 DR:5 LR:-23.36 LO:27.2);ALT=]chr16:9239910]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	43380609	+	chr11	43400778	+	.	12	0	4841357_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4841357_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:43380609(+)-11:43400778(-)__11_43365001_43390001D;SPAN=20169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:0 DR:12 LR:-24.71 LO:27.71);ALT=G[chr11:43400778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	43380665	+	chr11	43411200	+	GGATTCACCAATGAACTTGAAGCATCCTCATGACCTAGTCATATTAATGAGACAAGAAGCAACAGTTAACTACCTCAAAGAATTAG	0	21	4841359_1	58.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GGATTCACCAATGAACTTGAAGCATCCTCATGACCTAGTCATATTAATGAGACAAGAAGCAACAGTTAACTACCTCAAAGAATTAG;MAPQ=60;MATEID=4841359_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_43365001_43390001_105C;SPAN=30535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:41 GQ:38.6 PL:[58.4, 0.0, 38.6] SR:21 DR:0 LR:-58.37 LO:58.37);ALT=T[chr11:43411200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	43702537	+	chr11	43775594	+	TTGTCACAGGTAGTACTGATGGAATTGGAAAATCATATGCAGAAG	0	13	4842186_1	32.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTGTCACAGGTAGTACTGATGGAATTGGAAAATCATATGCAGAAG;MAPQ=60;MATEID=4842186_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_43757001_43782001_109C;SPAN=73057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:39 GQ:32.3 PL:[32.3, 0.0, 62.0] SR:13 DR:0 LR:-32.35 LO:32.87);ALT=G[chr11:43775594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	43902729	+	chr11	43904131	+	.	5	4	4842830_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4842830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_43879501_43904501_310C;SPAN=1402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:4 DR:5 LR:-2.788 LO:13.35);ALT=G[chr11:43904131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587286	+	chr11	44609022	+	.	35	11	4844335_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4844335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_44590001_44615001_66C;SPAN=21736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:11 DR:35 LR:-120.9 LO:120.9);ALT=G[chr11:44609022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587310	+	chr11	44616190	+	.	59	0	4844390_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4844390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:44587310(+)-11:44616190(-)__11_44614501_44639501D;SPAN=28880;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:55 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=G[chr11:44616190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587324	+	chr11	44621707	+	.	36	0	4844391_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4844391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:44587324(+)-11:44621707(-)__11_44614501_44639501D;SPAN=34383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:65 GQ:55.1 PL:[101.3, 0.0, 55.1] SR:0 DR:36 LR:-101.9 LO:101.9);ALT=A[chr11:44621707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44587334	+	chr11	44626607	+	.	8	0	4844392_1	13.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4844392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:44587334(+)-11:44626607(-)__11_44614501_44639501D;SPAN=39273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=G[chr11:44626607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44616275	+	chr11	44626608	+	ATCCTGGGCGCAGTGATCCTGGGCTTCGGGGTGTGGATCCTGGCCGACAAGAGCAGTTTCATCTCTGTCCTGC	0	75	4844398_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=ATCCTGGGCGCAGTGATCCTGGGCTTCGGGGTGTGGATCCTGGCCGACAAGAGCAGTTTCATCTCTGTCCTGC;MAPQ=60;MATEID=4844398_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_44614501_44639501_335C;SPAN=10333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:106 GQ:37.4 PL:[218.9, 0.0, 37.4] SR:75 DR:0 LR:-226.1 LO:226.1);ALT=T[chr11:44626608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	44636927	+	chr11	44639709	+	.	3	4	4844672_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGTGA;MAPQ=60;MATEID=4844672_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_44639001_44664001_325C;SPAN=2782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:37 GQ:9.8 PL:[9.8, 0.0, 79.1] SR:4 DR:3 LR:-9.782 LO:12.99);ALT=A[chr11:44639709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45429849	+	chr11	45431614	+	.	73	40	4846777_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCC;MAPQ=60;MATEID=4846777_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_45423001_45448001_5C;SPAN=1765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:23 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:40 DR:73 LR:-290.5 LO:290.5);ALT=C[chr11:45431614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45932513	+	chr11	45935369	+	.	0	13	4847869_1	23.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4847869_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_45913001_45938001_60C;SPAN=2856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:72 GQ:23.6 PL:[23.6, 0.0, 149.0] SR:13 DR:0 LR:-23.41 LO:28.82);ALT=C[chr11:45935369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45937388	+	chr11	45939249	+	ACAGGCAACTTTTTCCGAAGCTCCTTCCGTAGGATCCCGTCATTGAGCAGCACAAGCAGGTTAGAGGCAGAGTACACCAGCTCTGACAGCTCGTGCGAATCGGCGAATCG	0	32	4847891_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=ACAGGCAACTTTTTCCGAAGCTCCTTCCGTAGGATCCCGTCATTGAGCAGCACAAGCAGGTTAGAGGCAGAGTACACCAGCTCTGACAGCTCGTGCGAATCGGCGAATCG;MAPQ=60;MATEID=4847891_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_11_45913001_45938001_351C;SPAN=1861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:32 DR:0 LR:-99.02 LO:99.02);ALT=C[chr11:45939249[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45937909	+	chr11	45939319	+	.	30	0	4847893_1	88.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4847893_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:45937909(+)-11:45939319(-)__11_45913001_45938001D;SPAN=1410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:41 GQ:8.9 PL:[88.1, 0.0, 8.9] SR:0 DR:30 LR:-91.3 LO:91.3);ALT=A[chr11:45939319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	45987161	+	chr11	45991364	+	.	4	4	4847903_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4847903_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_45986501_46011501_269C;SPAN=4203;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:4 DR:4 LR:-0.8912 LO:13.07);ALT=T[chr11:45991364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	46958414	+	chr11	47073938	+	.	10	0	4851207_1	21.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4851207_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:46958414(+)-11:47073938(-)__11_47064501_47089501D;SPAN=115524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:44 GQ:21.2 PL:[21.2, 0.0, 83.9] SR:0 DR:10 LR:-21.09 LO:23.3);ALT=C[chr11:47073938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47236816	+	chr11	47237886	+	.	0	11	4851921_1	11.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=4851921_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47236001_47261001_377C;SPAN=1070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:11 DR:0 LR:-11.39 LO:22.24);ALT=T[chr11:47237886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47279681	+	chr11	47280730	+	.	0	4	4851714_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=4851714_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47260501_47285501_258C;SPAN=1049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:4 DR:0 LR:13.62 LO:6.133);ALT=G[chr11:47280730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47381592	+	chr11	47397184	+	.	2	78	4852586_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4852586_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47383001_47408001_357C;SPAN=15592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:70 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:78 DR:2 LR:-237.7 LO:237.7);ALT=C[chr11:47397184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47381644	+	chr11	47399859	+	.	51	0	4852587_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4852587_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:47381644(+)-11:47399859(-)__11_47383001_47408001D;SPAN=18215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:77 GQ:38.6 PL:[147.5, 0.0, 38.6] SR:0 DR:51 LR:-151.0 LO:151.0);ALT=G[chr11:47399859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47397283	+	chr11	47399860	+	.	0	94	4852643_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4852643_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47383001_47408001_285C;SPAN=2577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:162 GQ:99 PL:[266.6, 0.0, 124.7] SR:94 DR:0 LR:-269.1 LO:269.1);ALT=G[chr11:47399860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47405385	+	chr11	47417041	+	.	12	5	4852668_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4852668_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47383001_47408001_11C;SPAN=11656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:39 GQ:29 PL:[29.0, 0.0, 65.3] SR:5 DR:12 LR:-29.05 LO:29.82);ALT=T[chr11:47417041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47440751	+	chr11	47441815	+	.	0	30	4852820_1	77.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4852820_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47432001_47457001_420C;SPAN=1064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:82 GQ:77 PL:[77.0, 0.0, 119.9] SR:30 DR:0 LR:-76.81 LO:77.38);ALT=G[chr11:47441815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47446310	+	chr11	47447755	+	.	15	0	4852850_1	21.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=4852850_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:47446310(+)-11:47447755(-)__11_47432001_47457001D;SPAN=1445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:105 GQ:21.2 PL:[21.2, 0.0, 232.4] SR:0 DR:15 LR:-21.07 LO:31.57);ALT=G[chr11:47447755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47587407	+	chr11	47591248	+	.	27	0	4853497_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4853497_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:47587407(+)-11:47591248(-)__11_47579001_47604001D;SPAN=3841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:73 GQ:69.5 PL:[69.5, 0.0, 105.8] SR:0 DR:27 LR:-69.35 LO:69.81);ALT=G[chr11:47591248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47587539	+	chr11	47593018	+	AGTGGAAGAGACTAGGAGTCGAGCAGCTGCGGCTCAGCACAGTAGACATGACTGGGATCCCCACCTTGGACAACCTCCAGAAGGGAGTCCAATTTGCTCTCAAGTACCAGTCGCTGGGCCAGTGTGTTTACGTGCATTGTAAGGCTGGGCGCTCCAGGAGTGCCACTATGGTGGCAGCATACCTGA	0	52	4853499_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TTCAGGT;INSERTION=AGTGGAAGAGACTAGGAGTCGAGCAGCTGCGGCTCAGCACAGTAGACATGACTGGGATCCCCACCTTGGACAACCTCCAGAAGGGAGTCCAATTTGCTCTCAAGTACCAGTCGCTGGGCCAGTGTGTTTACGTGCATTGTAAGGCTGGGCGCTCCAGGAGTGCCACTATGGTGGCAGCATACCTGA;MAPQ=60;MATEID=4853499_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_47579001_47604001_148C;SPAN=5479;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:80 GQ:44.3 PL:[149.9, 0.0, 44.3] SR:52 DR:0 LR:-153.2 LO:153.2);ALT=G[chr11:47593018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47600711	+	chr11	47602077	+	GACTGGGCGACCCTCCGTTCTGTTGCTGCCGGTGAGGCGGGAGAGCGCCGGGGCCGACACGCGCC	60	55	4853543_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GACTGGGCGACCCTCCGTTCTGTTGCTGCCGGTGAGGCGGGAGAGCGCCGGGGCCGACACGCGCC;MAPQ=60;MATEID=4853543_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_47579001_47604001_182C;SPAN=1366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:127 DP:106 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:55 DR:60 LR:-376.3 LO:376.3);ALT=G[chr11:47602077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47604020	+	chr11	47605864	+	.	0	39	4852902_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4852902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47603501_47628501_82C;SPAN=1844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:84 GQ:96.2 PL:[106.1, 0.0, 96.2] SR:39 DR:0 LR:-106.0 LO:106.0);ALT=G[chr11:47605864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47612371	+	chr11	47615699	+	.	6	11	4852924_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTGG;MAPQ=60;MATEID=4852924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47603501_47628501_175C;SPAN=3328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:71 GQ:27.2 PL:[27.2, 0.0, 142.7] SR:11 DR:6 LR:-26.98 LO:31.63);ALT=G[chr11:47615699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47660605	+	chr11	47663929	+	.	35	30	4853303_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4853303_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47652501_47677501_379C;SPAN=3324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:91 GQ:84.5 PL:[134.0, 0.0, 84.5] SR:30 DR:35 LR:-134.3 LO:134.3);ALT=T[chr11:47663929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47776218	+	chr11	47786821	+	.	2	5	4853726_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4853726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47775001_47800001_399C;SPAN=10603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:79 GQ:1.5 PL:[0.0, 1.5, 194.7] SR:5 DR:2 LR:1.597 LO:10.88);ALT=T[chr11:47786821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47786916	+	chr11	47788621	+	.	0	20	4853770_1	43.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4853770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_47775001_47800001_39C;SPAN=1705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:84 GQ:43.4 PL:[43.4, 0.0, 158.9] SR:20 DR:0 LR:-43.26 LO:47.06);ALT=T[chr11:47788621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	47924170	+	chr19	57838857	-	.	4	26	6877244_1	85.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=AGTAGCTGGGATTACAGGC;MAPQ=31;MATEID=6877244_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_57820001_57845001_390C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:28 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:26 DR:4 LR:-85.82 LO:85.82);ALT=T]chr19:57838857];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	48600858	+	chr11	48604283	+	.	92	72	4856306_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=TC;MAPQ=60;MATEID=4856306_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_48583501_48608501_6C;SPAN=3425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:32 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:72 DR:92 LR:-373.0 LO:373.0);ALT=C[chr11:48604283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	48734780	+	chr11	48736949	+	.	58	11	4856572_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=TTCTCAGAAAGCTTCTTTCTAGTTTTTATTTGAAGATATTTCCTTTTT;MAPQ=60;MATEID=4856572_2;MATENM=1;NM=4;NUMPARTS=2;SCTG=c_11_48730501_48755501_161C;SPAN=2169;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:15 GQ:18.3 PL:[201.3, 18.3, 0.0] SR:11 DR:58 LR:-201.3 LO:201.3);ALT=T[chr11:48736949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57094365	+	chr11	57095768	+	CTTAGAAGACTCGCCTCGGCCCCCTTCATATTCTTTCATGGCTTTTTCATAGTCCCTCCTGGCATCCTCAGCCTTGCGATCCCACTCCTCTTTCTTCTCTTTGGACATTCCCTTCCAGATCTCGCCTGCCTTCTTGGAAAGATCCGTGATGCTGATGCCAGGATGGTCTGACTTGATCTTCTCTCGGCTGGCATTGAGCCACAGCATGTATGCAGACATGGGCCTCTTGGGGGCATTGGGGTCTTTGCCCTTCTT	0	15	4868706_1	22.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CACCT;INSERTION=CTTAGAAGACTCGCCTCGGCCCCCTTCATATTCTTTCATGGCTTTTTCATAGTCCCTCCTGGCATCCTCAGCCTTGCGATCCCACTCCTCTTTCTTCTCTTTGGACATTCCCTTCCAGATCTCGCCTGCCTTCTTGGAAAGATCCGTGATGCTGATGCCAGGATGGTCTGACTTGATCTTCTCTCGGCTGGCATTGAGCCACAGCATGTATGCAGACATGGGCCTCTTGGGGGCATTGGGGTCTTTGCCCTTCTT;MAPQ=60;MATEID=4868706_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_57085001_57110001_44C;SPAN=1403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:102 GQ:22.1 PL:[22.1, 0.0, 223.4] SR:15 DR:0 LR:-21.88 LO:31.78);ALT=T[chr11:57095768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57296394	+	chr11	57297592	+	.	0	39	4869171_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=4869171_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_57281001_57306001_104C;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:100 GQ:99 PL:[101.6, 0.0, 141.2] SR:39 DR:0 LR:-101.6 LO:102.0);ALT=G[chr11:57297592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57296438	+	chr11	57298129	+	.	32	0	4869172_1	83.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4869172_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57296438(+)-11:57298129(-)__11_57281001_57306001D;SPAN=1691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:80 GQ:83.9 PL:[83.9, 0.0, 110.3] SR:0 DR:32 LR:-83.96 LO:84.15);ALT=T[chr11:57298129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57322144	+	chr11	57335056	+	.	88	0	4869296_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4869296_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57322144(+)-11:57335056(-)__11_57330001_57355001D;SPAN=12912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:55 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:0 DR:88 LR:-260.8 LO:260.8);ALT=T[chr11:57335056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57327907	+	chr11	57335057	+	.	25	3	4869297_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=4869297_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACCAC;SCTG=c_11_57330001_57355001_13C;SPAN=7150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:55 GQ:45.1 PL:[52.9, 0.0, 45.1] SR:3 DR:25 LR:-52.78 LO:52.78);ALT=T[chr11:57335057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	71492565	+	chr11	57343970	+	.	8	0	7447647_1	0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=7447647_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57343970(-)-23:71492565(+)__23_71491001_71516001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:628 GQ:99 PL:[0.0, 143.5, 1812.0] SR:0 DR:8 LR:143.7 LO:8.283);ALT=]chrX:71492565]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	57425356	+	chr11	57426924	+	.	8	0	4869616_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4869616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:57425356(+)-11:57426924(-)__11_57403501_57428501D;SPAN=1568;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=C[chr11:57426924[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	57472703	+	chr11	57479433	+	.	3	6	4869907_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4869907_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_57477001_57502001_263C;SPAN=6730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:6 DR:3 LR:-19.14 LO:21.04);ALT=T[chr11:57479433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	58166999	+	chr11	58168150	+	.	0	49	4871618_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGTACTAAAGATTTTAT;MAPQ=60;MATEID=4871618_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_11_58163001_58188001_271C;SPAN=1151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:28 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:49 DR:0 LR:-145.2 LO:145.2);ALT=T[chr11:58168150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	58322415	+	chr11	58338028	+	GTAGACATTGAGCTCCTGGATATTGGTAGTATACACGAGCTGCG	0	18	4872001_1	48.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GTAGACATTGAGCTCCTGGATATTGGTAGTATACACGAGCTGCG;MAPQ=60;MATEID=4872001_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_58334501_58359501_176C;SPAN=15613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:41 GQ:48.5 PL:[48.5, 0.0, 48.5] SR:18 DR:0 LR:-48.31 LO:48.32);ALT=T[chr11:58338028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	58338238	+	chr11	58343254	+	.	30	0	4872011_1	82.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4872011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:58338238(+)-11:58343254(-)__11_58334501_58359501D;SPAN=5016;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:63 GQ:68.9 PL:[82.1, 0.0, 68.9] SR:0 DR:30 LR:-82.0 LO:82.0);ALT=A[chr11:58343254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	58594188	+	chr11	58596020	+	.	90	62	4872674_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4872674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_58579501_58604501_80C;SPAN=1832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:30 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:62 DR:90 LR:-369.7 LO:369.7);ALT=T[chr11:58596020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59575324	+	chr11	59577328	+	.	0	19	4874773_1	41.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4874773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59559501_59584501_72C;SPAN=2004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:81 GQ:41 PL:[41.0, 0.0, 153.2] SR:19 DR:0 LR:-40.77 LO:44.56);ALT=T[chr11:59577328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59575370	+	chr11	59578076	+	.	15	0	4874774_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4874774_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:59575370(+)-11:59578076(-)__11_59559501_59584501D;SPAN=2706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:111 GQ:19.7 PL:[19.7, 0.0, 247.4] SR:0 DR:15 LR:-19.44 LO:31.18);ALT=A[chr11:59578076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59940602	+	chr11	59942874	+	.	6	7	4875754_1	21.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4875754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59927001_59952001_261C;SPAN=2272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:81 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:7 DR:6 LR:-20.97 LO:28.08);ALT=C[chr11:59942874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59943085	+	chr11	59947304	+	AAAAGCTTGGTCAACCTTTTCTCTGTGGCGATTGATAGAGAGCCAGAGATGATAAA	4	15	4875760_1	35.0	.	DISC_MAPQ=48;EVDNC=TSI_G;HOMSEQ=CACC;INSERTION=AAAAGCTTGGTCAACCTTTTCTCTGTGGCGATTGATAGAGAGCCAGAGATGATAAA;MAPQ=60;MATEID=4875760_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_59927001_59952001_282C;SPAN=4219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:15 DR:4 LR:-35.58 LO:40.99);ALT=C[chr11:59947304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59945790	+	chr11	59949054	+	.	2	7	4875771_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4875771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59927001_59952001_204C;SPAN=3264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:7 DR:2 LR:-3.158 LO:17.1);ALT=C[chr11:59949054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59947439	+	chr11	59949054	+	.	7	48	4875780_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4875780_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59927001_59952001_276C;SPAN=1615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:101 GQ:98.3 PL:[144.5, 0.0, 98.3] SR:48 DR:7 LR:-144.7 LO:144.7);ALT=C[chr11:59949054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59947487	+	chr11	59950450	+	.	26	0	4875781_1	61.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4875781_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:59947487(+)-11:59950450(-)__11_59927001_59952001D;SPAN=2963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:91 GQ:61.4 PL:[61.4, 0.0, 157.1] SR:0 DR:26 LR:-61.17 LO:63.6);ALT=G[chr11:59950450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59949216	+	chr11	59950451	+	.	111	16	4875786_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4875786_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_59927001_59952001_152C;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:114 DP:100 GQ:30.6 PL:[336.6, 30.6, 0.0] SR:16 DR:111 LR:-336.7 LO:336.7);ALT=T[chr11:59950451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	59997546	+	chr11	60010431	+	.	23	8	4875885_1	75.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4875885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_60000501_60025501_289C;SPAN=12885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:26 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:8 DR:23 LR:-75.92 LO:75.92);ALT=T[chr11:60010431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60146137	+	chr11	60150599	+	.	12	1	4876250_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=4876250_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_60147501_60172501_277C;SPAN=4462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:1 DR:12 LR:-28.83 LO:30.91);ALT=G[chr11:60150599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60150761	+	chr11	60156863	+	TTTGGCATTACTGGATCCCTCTCAATTATCTCTGGAAAACAATCAACTAAGCCCTTT	4	9	4876257_1	13.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTGGCATTACTGGATCCCTCTCAATTATCTCTGGAAAACAATCAACTAAGCCCTTT;MAPQ=60;MATEID=4876257_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_60147501_60172501_157C;SPAN=6102;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:9 DR:4 LR:-12.96 LO:20.79);ALT=G[chr11:60156863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60671333	+	chr11	60673836	+	.	20	16	4877243_1	79.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=4877243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_60662001_60687001_201C;SPAN=2503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:74 GQ:79.1 PL:[79.1, 0.0, 98.9] SR:16 DR:20 LR:-78.98 LO:79.13);ALT=A[chr11:60673836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60681765	+	chr11	60687155	+	.	40	0	4877513_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4877513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:60681765(+)-11:60687155(-)__11_60686501_60711501D;SPAN=5390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:40 LR:-130.9 LO:130.9);ALT=G[chr11:60687155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	60857830	-	chr11	60859316	+	CGCACCCCCCAT	7	15	4877985_1	24.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=TGGTGGGGGGTG;INSERTION=CGCACCCCCCAT;MAPQ=60;MATEID=4877985_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_60833501_60858501_295C;SPAN=1486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:153 GQ:24.8 PL:[24.8, 0.0, 344.9] SR:15 DR:7 LR:-24.57 LO:41.26);ALT=[chr11:60859316[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	60859356	+	chr11	60857833	+	A	7	26	4877986_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CACCCCCCACCA;INSERTION=A;MAPQ=60;MATEID=4877986_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGGGGG;SCTG=c_11_60833501_60858501_71C;SPAN=1523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:189 GQ:27 PL:[27.0, 0.0, 313.1] SR:26 DR:7 LR:-26.86 LO:43.77);ALT=]chr11:60859356]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	60857882	+	chr11	60859356	-	CGCACCCCCCAT	6	19	4877988_1	30.0	.	DISC_MAPQ=52;EVDNC=TSI_L;INSERTION=CGCACCCCCCAT;MAPQ=60;MATEID=4877988_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_11_60833501_60858501_295C;SPAN=1474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:182 GQ:30.1 PL:[30.1, 0.0, 409.7] SR:19 DR:6 LR:-29.92 LO:49.61);ALT=C]chr11:60859356];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	60868963	+	chr11	60866748	+	.	8	0	4878209_1	0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=4878209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:60866748(-)-11:60868963(+)__11_60858001_60883001D;SPAN=2215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=]chr11:60868963]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	61081966	+	chr11	61083760	+	.	3	2	4878568_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GATAA;MAPQ=60;MATEID=4878568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61078501_61103501_256C;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:95 GQ:9 PL:[0.0, 9.0, 247.5] SR:2 DR:3 LR:9.233 LO:8.25);ALT=A[chr11:61083760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61100795	+	chr11	61102089	+	.	10	0	4878621_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4878621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61100795(+)-11:61102089(-)__11_61078501_61103501D;SPAN=1294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:0 DR:10 LR:-12.96 LO:20.79);ALT=G[chr11:61102089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61100812	+	chr11	61105411	+	.	10	0	4878711_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4878711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61100812(+)-11:61105411(-)__11_61103001_61128001D;SPAN=4599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:40 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-22.17 LO:23.78);ALT=G[chr11:61105411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61102203	+	chr11	61105412	+	.	0	14	4878712_1	35.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4878712_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61103001_61128001_191C;SPAN=3209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:39 GQ:35.6 PL:[35.6, 0.0, 58.7] SR:14 DR:0 LR:-35.65 LO:35.96);ALT=G[chr11:61105412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61129944	+	chr11	61131774	+	.	8	0	4879353_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4879353_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61129944(+)-11:61131774(-)__11_61127501_61152501D;SPAN=1830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=G[chr11:61131774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61197689	+	chr11	61213409	+	.	19	0	4878933_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4878933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61197689(+)-11:61213409(-)__11_61201001_61226001D;SPAN=15720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:42 GQ:48.2 PL:[51.5, 0.0, 48.2] SR:0 DR:19 LR:-51.34 LO:51.34);ALT=G[chr11:61213409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61197689	+	chr11	61204381	+	.	27	0	4878932_1	78.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4878932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61197689(+)-11:61204381(-)__11_61201001_61226001D;SPAN=6692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:39 GQ:15.8 PL:[78.5, 0.0, 15.8] SR:0 DR:27 LR:-80.89 LO:80.89);ALT=G[chr11:61204381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61432089	-	chr11	61433848	+	.	9	0	4879851_1	8.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4879851_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61432089(-)-11:61433848(-)__11_61421501_61446501D;SPAN=1759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:77 GQ:8.9 PL:[8.9, 0.0, 177.2] SR:0 DR:9 LR:-8.848 LO:18.1);ALT=[chr11:61433848[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	61556754	+	chr11	61560026	+	.	17	0	4880058_1	12.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=4880058_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61556754(+)-11:61560026(-)__11_61544001_61569001D;SPAN=3272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:162 GQ:12.4 PL:[12.4, 0.0, 378.8] SR:0 DR:17 LR:-12.23 LO:33.34);ALT=C[chr11:61560026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61557426	+	chr11	61560024	+	.	87	0	4880064_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=4880064_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61557426(+)-11:61560024(-)__11_61544001_61569001D;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:158 GQ:99 PL:[244.4, 0.0, 138.8] SR:0 DR:87 LR:-245.9 LO:245.9);ALT=T[chr11:61560024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61558075	+	chr11	61560027	+	.	36	50	4880068_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4880068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_61544001_61569001_50C;SPAN=1952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:191 GQ:99 PL:[209.3, 0.0, 252.2] SR:50 DR:36 LR:-209.0 LO:209.3);ALT=C[chr11:61560027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61560499	+	chr11	61562812	+	.	16	0	4880074_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4880074_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:61560499(+)-11:61562812(-)__11_61544001_61569001D;SPAN=2313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:78 GQ:31.7 PL:[31.7, 0.0, 157.1] SR:0 DR:16 LR:-31.68 LO:36.46);ALT=A[chr11:61562812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	61841813	+	chr14	81786774	+	C	43	42	5819167_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=5819167_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_81781001_81806001_356C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:32 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:42 DR:43 LR:-221.2 LO:221.2);ALT=G[chr14:81786774[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	62105641	+	chr11	62123795	+	.	3	10	4881869_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=4881869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62107501_62132501_74C;SPAN=18154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:37 GQ:29.6 PL:[29.6, 0.0, 59.3] SR:10 DR:3 LR:-29.59 LO:30.16);ALT=T[chr11:62123795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62301547	+	chr11	62303416	+	AGAACCACTTCAGAGCTGCAGGAGCTGAAGACTTCACGGGTCCAGGTCTGGCCAGGCTCGGGAGAGCGGTCCCCCTTGCGGTGCAGCTTCAGGCCCACCGTGTGGTGCCCCATGGTGTTCAGCAGCTGGGTCACCTCACCCGACTGCAGGTTGTCAAAGTAGATGGTGGCACCCACAATCTGGTCC	2	10	4882564_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AGAACCACTTCAGAGCTGCAGGAGCTGAAGACTTCACGGGTCCAGGTCTGGCCAGGCTCGGGAGAGCGGTCCCCCTTGCGGTGCAGCTTCAGGCCCACCGTGTGGTGCCCCATGGTGTTCAGCAGCTGGGTCACCTCACCCGACTGCAGGTTGTCAAAGTAGATGGTGGCACCCACAATCTGGTCC;MAPQ=60;MATEID=4882564_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_62303501_62328501_231C;SPAN=1869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:4 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:10 DR:2 LR:-29.71 LO:29.71);ALT=C[chr11:62303416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62303619	+	chr11	62314128	+	.	22	0	4882568_1	50.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4882568_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62303619(+)-11:62314128(-)__11_62303501_62328501D;SPAN=10509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:81 GQ:50.9 PL:[50.9, 0.0, 143.3] SR:0 DR:22 LR:-50.68 LO:53.24);ALT=C[chr11:62314128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62304041	+	chr11	62314130	+	.	0	28	4882571_1	73.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4882571_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62303501_62328501_188C;SPAN=10089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:71 GQ:73.4 PL:[73.4, 0.0, 96.5] SR:28 DR:0 LR:-73.19 LO:73.41);ALT=T[chr11:62314130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62430805	+	chr11	62432319	+	.	0	22	4883104_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=4883104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62426001_62451001_143C;SPAN=1514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:81 GQ:50.9 PL:[50.9, 0.0, 143.3] SR:22 DR:0 LR:-50.68 LO:53.24);ALT=C[chr11:62432319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62430848	+	chr11	62432600	+	.	31	0	4883105_1	80.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4883105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62430848(+)-11:62432600(-)__11_62426001_62451001D;SPAN=1752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:83 GQ:80 PL:[80.0, 0.0, 119.6] SR:0 DR:31 LR:-79.84 LO:80.32);ALT=C[chr11:62432600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62491899	+	chr11	62494090	+	.	5	4	4882949_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=4882949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62475001_62500001_311C;SPAN=2191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:81 GQ:1.8 PL:[0.0, 1.8, 198.0] SR:4 DR:5 LR:2.139 LO:10.82);ALT=C[chr11:62494090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62529157	+	chr11	62530336	+	.	69	0	4883505_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4883505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62529157(+)-11:62530336(-)__11_62524001_62549001D;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:69 DP:112 GQ:72.2 PL:[197.6, 0.0, 72.2] SR:0 DR:69 LR:-200.5 LO:200.5);ALT=A[chr11:62530336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62529378	+	chr11	62533123	+	ATGGCTTTGTAATTGCTGTCACCACCATTGACAATATTGGTGCTGGTGTGATCCAGCCAGGCCGAGGCTTTGTCCTTTATCCAGTTAAGTACAAGGCCATTGTTTTCCGGCCATTTAAAGGGGAGGTCGTGGATGCTGTTGTCACTCAGGTCAACAAGGTTGGACTCTTCACAGAAATTGGGCCCATGTCTTGCTTCATCTCTCGACATTCCATCCCTTCAGAGATGGAGTTTGATCCTAACTCCAACCCACCATGTTACAAGACAATGGATG	0	96	4883509_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGGCTTTGTAATTGCTGTCACCACCATTGACAATATTGGTGCTGGTGTGATCCAGCCAGGCCGAGGCTTTGTCCTTTATCCAGTTAAGTACAAGGCCATTGTTTTCCGGCCATTTAAAGGGGAGGTCGTGGATGCTGTTGTCACTCAGGTCAACAAGGTTGGACTCTTCACAGAAATTGGGCCCATGTCTTGCTTCATCTCTCGACATTCCATCCCTTCAGAGATGGAGTTTGATCCTAACTCCAACCCACCATGTTACAAGACAATGGATG;MAPQ=60;MATEID=4883509_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_11_62524001_62549001_217C;SPAN=3745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:116 GQ:4.8 PL:[290.4, 4.8, 0.0] SR:96 DR:0 LR:-304.2 LO:304.2);ALT=T[chr11:62533123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62555000	+	chr11	62556492	+	.	104	25	4883323_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4883323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_62548501_62573501_83C;SPAN=1492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:94 GQ:30 PL:[330.0, 30.0, 0.0] SR:25 DR:104 LR:-330.1 LO:330.1);ALT=G[chr11:62556492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	62621802	+	chr11	62622855	+	.	30	0	4883728_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4883728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:62621802(+)-11:62622855(-)__11_62597501_62622501D;SPAN=1053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:49 GQ:32.9 PL:[85.7, 0.0, 32.9] SR:0 DR:30 LR:-87.03 LO:87.03);ALT=G[chr11:62622855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63088186	-	chr11	63089363	+	.	8	0	4884986_1	8.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4884986_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63088186(-)-11:63089363(-)__11_63087501_63112501D;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=[chr11:63089363[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	63304400	+	chr11	63306994	+	.	11	0	4885569_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4885569_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63304400(+)-11:63306994(-)__11_63283501_63308501D;SPAN=2594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:0 DR:11 LR:-15.72 LO:23.22);ALT=C[chr11:63306994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63304400	+	chr11	63312092	+	.	41	0	4885570_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4885570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63304400(+)-11:63312092(-)__11_63283501_63308501D;SPAN=7692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:35 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=C[chr11:63312092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63307098	+	chr11	63312093	+	.	3	25	4885575_1	81.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=4885575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63283501_63308501_346C;SPAN=4995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:41 GQ:15.5 PL:[81.5, 0.0, 15.5] SR:25 DR:3 LR:-83.57 LO:83.57);ALT=T[chr11:63312093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63312363	+	chr11	63313618	+	.	0	7	4885365_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=4885365_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_63308001_63333001_265C;SPAN=1255;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:80 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:7 DR:0 LR:-1.433 LO:13.15);ALT=T[chr11:63313618[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63426726	+	chr11	63438762	+	.	6	5	4886030_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4886030_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63430501_63455501_9C;SPAN=12036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:36 GQ:16.7 PL:[16.7, 0.0, 69.5] SR:5 DR:6 LR:-16.65 LO:18.55);ALT=T[chr11:63438762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63449188	+	chr11	63517460	+	.	23	0	4886202_1	67.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=4886202_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63449188(+)-11:63517460(-)__11_63504001_63529001D;SPAN=68272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:33 GQ:11 PL:[67.1, 0.0, 11.0] SR:0 DR:23 LR:-69.03 LO:69.03);ALT=G[chr11:63517460[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63742267	+	chr11	63743696	+	.	138	160	4886969_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4886969_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63724501_63749501_182C;SPAN=1429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:260 DP:248 GQ:70.3 PL:[772.3, 70.3, 0.0] SR:160 DR:138 LR:-772.4 LO:772.4);ALT=G[chr11:63743696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63754008	+	chr11	63755818	+	.	44	0	4887026_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4887026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63754008(+)-11:63755818(-)__11_63749001_63774001D;SPAN=1810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:73 GQ:49.7 PL:[125.6, 0.0, 49.7] SR:0 DR:44 LR:-127.1 LO:127.1);ALT=T[chr11:63755818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63754037	+	chr11	63763998	+	.	35	0	4887027_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4887027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63754037(+)-11:63763998(-)__11_63749001_63774001D;SPAN=9961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:89 GQ:91.4 PL:[91.4, 0.0, 124.4] SR:0 DR:35 LR:-91.42 LO:91.7);ALT=G[chr11:63763998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63755870	+	chr11	63764000	+	ATTGCTGTGCAGAACCCTCTGGTGTCAGAGCGGCTGGAGCTCTCGGTCCTATACAAGGAGTATGCTGAAGATGACAACATCTATCAACAGAAGATCA	0	70	4887032_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTGCTGTGCAGAACCCTCTGGTGTCAGAGCGGCTGGAGCTCTCGGTCCTATACAAGGAGTATGCTGAAGATGACAACATCTATCAACAGAAGATCA;MAPQ=60;MATEID=4887032_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_63749001_63774001_145C;SPAN=8130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:112 GQ:68.9 PL:[200.9, 0.0, 68.9] SR:70 DR:0 LR:-204.1 LO:204.1);ALT=G[chr11:63764000[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63923406	-	chr11	63924524	+	.	13	0	4887621_1	20.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=4887621_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63923406(-)-11:63924524(-)__11_63920501_63945501D;SPAN=1118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:83 GQ:20.6 PL:[20.6, 0.0, 179.0] SR:0 DR:13 LR:-20.43 LO:27.93);ALT=[chr11:63924524[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	63953771	+	chr11	63960545	+	.	28	0	4887856_1	68.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4887856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63953771(+)-11:63960545(-)__11_63945001_63970001D;SPAN=6774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:90 GQ:68 PL:[68.0, 0.0, 150.5] SR:0 DR:28 LR:-68.05 LO:69.75);ALT=C[chr11:63960545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63962093	+	chr11	63963117	+	.	2	8	4887891_1	5.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4887891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63945001_63970001_233C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:8 DR:2 LR:-5.276 LO:15.61);ALT=G[chr11:63963117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63974315	+	chr11	63978082	+	.	14	0	4887541_1	24.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4887541_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63974315(+)-11:63978082(-)__11_63969501_63994501D;SPAN=3767;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:82 GQ:24.2 PL:[24.2, 0.0, 172.7] SR:0 DR:14 LR:-24.0 LO:30.65);ALT=G[chr11:63978082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63974996	+	chr11	63978083	+	.	0	41	4887542_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4887542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63969501_63994501_315C;SPAN=3087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:93 GQ:99 PL:[110.3, 0.0, 113.6] SR:41 DR:0 LR:-110.1 LO:110.2);ALT=A[chr11:63978083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63992482	+	chr11	63993549	+	.	8	0	4887597_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4887597_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63992482(+)-11:63993549(-)__11_63969501_63994501D;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:0 DR:8 LR:-6.089 LO:15.75);ALT=G[chr11:63993549[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	63995142	+	chr11	63996717	+	.	0	7	4887927_1	2.0	.	EVDNC=ASSMB;HOMSEQ=AGGTGA;MAPQ=60;MATEID=4887927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63994001_64019001_145C;SPAN=1575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:7 DR:0 LR:-2.788 LO:13.35);ALT=A[chr11:63996717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64000338	+	chr11	64001363	+	.	0	16	4887946_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=4887946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63994001_64019001_287C;SPAN=1025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:84 GQ:30.2 PL:[30.2, 0.0, 172.1] SR:16 DR:0 LR:-30.06 LO:35.88);ALT=G[chr11:64001363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64008604	+	chr11	64009854	+	.	0	7	4887965_1	2.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4887965_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_63994001_64019001_25C;SPAN=1250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:76 GQ:2.6 PL:[2.6, 0.0, 180.8] SR:7 DR:0 LR:-2.517 LO:13.31);ALT=G[chr11:64009854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64039277	+	chr11	64051653	+	.	0	16	4887757_1	43.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=4887757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64043001_64068001_321C;SPAN=12376;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:34 GQ:37.1 PL:[43.7, 0.0, 37.1] SR:16 DR:0 LR:-43.62 LO:43.62);ALT=T[chr11:64051653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64085858	+	chr11	64088131	+	.	29	9	4888483_1	81.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4888483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64067501_64092501_442C;SPAN=2273;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:149 GQ:81.8 PL:[81.8, 0.0, 279.8] SR:9 DR:29 LR:-81.77 LO:87.85);ALT=G[chr11:64088131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64085861	+	chr11	64087204	+	.	104	121	4888484_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGGTG;MAPQ=60;MATEID=4888484_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=GAGA;SCTG=c_11_64067501_64092501_370C;SPAN=1343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:180 DP:176 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:121 DR:104 LR:-534.7 LO:534.7);ALT=G[chr11:64087204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64494604	+	chr11	64496335	+	ATCTATTACAAGTGGATGTCAAACACCCCATCCTCCACCGTCTGTACCTCCTCCTCACGGATCT	3	20	4889284_1	43.0	.	DISC_MAPQ=42;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATCTATTACAAGTGGATGTCAAACACCCCATCCTCCACCGTCTGTACCTCCTCCTCACGGATCT;MAPQ=60;MATEID=4889284_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_11_64484001_64509001_79C;SPAN=1731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:96 GQ:43.4 PL:[43.4, 0.0, 188.6] SR:20 DR:3 LR:-43.31 LO:48.52);ALT=C[chr11:64496335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64496516	+	chr11	64497525	+	CGGCATTTGAGGCCCTGCTTGTAGATGCCCAGGAT	5	5	4889294_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CGGCATTTGAGGCCCTGCTTGTAGATGCCCAGGAT;MAPQ=60;MATEID=4889294_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_64484001_64509001_61C;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:5 DR:5 LR:-6.139 LO:17.59);ALT=T[chr11:64497525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64508973	+	chr11	64510266	+	ATGTGGAGCAGCTTGGCCGCCAG	3	25	4889360_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATGTGGAGCAGCTTGGCCGCCAG;MAPQ=60;MATEID=4889360_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64508501_64533501_255C;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:87 GQ:65.6 PL:[65.6, 0.0, 144.8] SR:25 DR:3 LR:-65.56 LO:67.23);ALT=G[chr11:64510266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64510370	+	chr11	64512212	+	.	10	0	4889367_1	16.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4889367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:64510370(+)-11:64512212(-)__11_64508501_64533501D;SPAN=1842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.75 LO:21.78);ALT=C[chr11:64512212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64532990	+	chr11	64534371	+	.	5	5	4889513_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4889513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64533001_64558001_59C;SPAN=1381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:5 DR:5 LR:-10.2 LO:18.38);ALT=C[chr11:64534371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64537884	+	chr11	64543970	+	CCTCAGGGTTAGGGGGGATGCCCAGGTCTCCTGTGCGCAGTTTACGAGTCAGGTCTTCTATCTGCAGTTGCA	6	12	4889527_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCTCAGGGTTAGGGGGGATGCCCAGGTCTCCTGTGCGCAGTTTACGAGTCAGGTCTTCTATCTGCAGTTGCA;MAPQ=60;MATEID=4889527_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_64533001_64558001_11C;SPAN=6086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:106 GQ:27.5 PL:[27.5, 0.0, 228.8] SR:12 DR:6 LR:-27.4 LO:36.71);ALT=T[chr11:64543970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64544099	+	chr11	64545834	+	.	111	93	4889559_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4889559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64533001_64558001_3C;SPAN=1735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:160 DP:106 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:93 DR:111 LR:-475.3 LO:475.3);ALT=C[chr11:64545834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64781744	+	chr11	64787889	+	TGGCCTGGACAATGCTGGAAAGACAACCATCCTGAAGAAGTTCAATGGGGAGGACATCGACACCATCTCCCCAACGCTGGGCTTCAACATCAAGACCCTGGAGCACCGAGGATTCAAGCTGAACATCTGGGATGTGGGTGGCCAGAAGTCCCTGCGGTCCTACTGGCGGAACTACTTTGAGAGCACCGATGGCCTCATCTGGGTAGTGGACAGCGCAGACCGCCAGCGCATGCAGGACTGCCAGCGGGAGCTCCAGAGCCTGCTGGTGGAGG	2	34	4890442_1	91.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGGCCTGGACAATGCTGGAAAGACAACCATCCTGAAGAAGTTCAATGGGGAGGACATCGACACCATCTCCCCAACGCTGGGCTTCAACATCAAGACCCTGGAGCACCGAGGATTCAAGCTGAACATCTGGGATGTGGGTGGCCAGAAGTCCCTGCGGTCCTACTGGCGGAACTACTTTGAGAGCACCGATGGCCTCATCTGGGTAGTGGACAGCGCAGACCGCCAGCGCATGCAGGACTGCCAGCGGGAGCTCCAGAGCCTGCTGGTGGAGG;MAPQ=60;MATEID=4890442_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_64778001_64803001_34C;SPAN=6145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:76 GQ:91.7 PL:[91.7, 0.0, 91.7] SR:34 DR:2 LR:-91.64 LO:91.65);ALT=T[chr11:64787889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64781744	+	chr11	64785836	+	.	114	21	4890441_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=4890441_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_11_64778001_64803001_34C;SPAN=4092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:88 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:21 DR:114 LR:-356.5 LO:356.5);ALT=T[chr11:64785836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64787972	+	chr11	64789195	+	C	4	2	4890458_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=4890458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64778001_64803001_108C;SPAN=1223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:101 GQ:7.2 PL:[0.0, 7.2, 257.4] SR:2 DR:4 LR:7.557 LO:10.22);ALT=G[chr11:64789195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64795057	+	chr11	64799900	+	.	11	0	4890474_1	8.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4890474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:64795057(+)-11:64799900(-)__11_64778001_64803001D;SPAN=4843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:104 GQ:8.3 PL:[8.3, 0.0, 242.6] SR:0 DR:11 LR:-8.135 LO:21.61);ALT=G[chr11:64799900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64814004	+	chr11	64815119	+	.	11	2	4890114_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGGGG;MAPQ=60;MATEID=4890114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64802501_64827501_235C;SPAN=1115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:84 GQ:17 PL:[17.0, 0.0, 185.3] SR:2 DR:11 LR:-16.85 LO:25.26);ALT=G[chr11:64815119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	64889896	+	chr11	64891973	+	.	9	3	4890621_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4890621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_64876001_64901001_53C;SPAN=2077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:3 DR:9 LR:-4.784 LO:17.36);ALT=G[chr11:64891973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65101429	+	chr11	65108433	+	.	9	0	4891311_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4891311_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65101429(+)-11:65108433(-)__11_65096501_65121501D;SPAN=7004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=T[chr11:65108433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65405690	+	chr11	65408333	+	.	10	0	4892275_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4892275_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65405690(+)-11:65408333(-)__11_65390501_65415501D;SPAN=2643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:0 DR:10 LR:-18.11 LO:22.2);ALT=C[chr11:65408333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65623202	+	chr11	65625567	+	AGAAGATAAACACCAGATCCTCCTTCTTGCTCTCCTTGGTCTCATAGGTTGCATCATAGAGGGCATAGCGGCAGTCCTTATCTGGCAGCATCTTGACAAAGGTGGCGTAGGGGTCGTCGACAGTCTGGCCCACATCGCCCACCAGGATCTCCTTGCCCTCCTCCAGGATGATGTTCTTCTTGTCCTCACTCAGGCAGAAGAGCACCGCCTTCTTGCGCTTCTTCACCTCCTCTGGCGTTGAAGACTTACGCACCTTCATGTCGTTGAACACCTTGATGACACCATCAGAGACAGCCACACCGGAGG	9	83	4893126_1	99.0	.	DISC_MAPQ=18;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AGAAGATAAACACCAGATCCTCCTTCTTGCTCTCCTTGGTCTCATAGGTTGCATCATAGAGGGCATAGCGGCAGTCCTTATCTGGCAGCATCTTGACAAAGGTGGCGTAGGGGTCGTCGACAGTCTGGCCCACATCGCCCACCAGGATCTCCTTGCCCTCCTCCAGGATGATGTTCTTCTTGTCCTCACTCAGGCAGAAGAGCACCGCCTTCTTGCGCTTCTTCACCTCCTCTGGCGTTGAAGACTTACGCACCTTCATGTCGTTGAACACCTTGATGACACCATCAGAGACAGCCACACCGGAGG;MAPQ=60;MATEID=4893126_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_65611001_65636001_75C;SPAN=2365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:106 GQ:4.4 PL:[251.9, 0.0, 4.4] SR:83 DR:9 LR:-266.3 LO:266.3);ALT=C[chr11:65625567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65623714	+	chr11	65625567	+	.	195	41	4893129_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=4893129_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_11_65611001_65636001_75C;SPAN=1853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:218 DP:134 GQ:58.9 PL:[646.9, 58.9, 0.0] SR:41 DR:195 LR:-647.0 LO:647.0);ALT=C[chr11:65625567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65647392	+	chr11	65649642	+	.	16	0	4893282_1	22.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4893282_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65647392(+)-11:65649642(-)__11_65635501_65660501D;SPAN=2250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:112 GQ:22.7 PL:[22.7, 0.0, 247.1] SR:0 DR:16 LR:-22.47 LO:33.68);ALT=A[chr11:65649642[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65647456	+	chr11	65648875	+	.	68	0	4893284_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893284_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65647456(+)-11:65648875(-)__11_65635501_65660501D;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:116 GQ:87.5 PL:[193.1, 0.0, 87.5] SR:0 DR:68 LR:-195.1 LO:195.1);ALT=G[chr11:65648875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65647757	+	chr11	65649643	+	AGCATGCTCACCGCCTGGACATCTTTGCCCACAACCTGGCCCAGGCTCAGAGGCTGCAGGAGGAGGACTTGGGCACAGCTGAGTTTGGGGTGACTCCATTCAGTGACCTCA	0	157	4893286_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AGCATGCTCACCGCCTGGACATCTTTGCCCACAACCTGGCCCAGGCTCAGAGGCTGCAGGAGGAGGACTTGGGCACAGCTGAGTTTGGGGTGACTCCATTCAGTGACCTCA;MAPQ=60;MATEID=4893286_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_65635501_65660501_63C;SPAN=1886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:157 DP:109 GQ:42.4 PL:[465.4, 42.4, 0.0] SR:157 DR:0 LR:-465.4 LO:465.4);ALT=G[chr11:65649643[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65767966	+	chr11	65769541	+	.	9	0	4893724_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893724_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65767966(+)-11:65769541(-)__11_65758001_65783001D;SPAN=1575;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:68 GQ:11.3 PL:[11.3, 0.0, 153.2] SR:0 DR:9 LR:-11.29 LO:18.62);ALT=G[chr11:65769541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65820009	+	chr11	65822541	+	.	34	0	4893634_1	85.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893634_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65820009(+)-11:65822541(-)__11_65807001_65832001D;SPAN=2532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:99 GQ:85.4 PL:[85.4, 0.0, 154.7] SR:0 DR:34 LR:-85.41 LO:86.51);ALT=A[chr11:65822541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65820575	+	chr11	65822542	+	.	3	49	4893637_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACAG;MAPQ=60;MATEID=4893637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_65807001_65832001_62C;SPAN=1967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:116 GQ:99 PL:[140.3, 0.0, 140.3] SR:49 DR:3 LR:-140.2 LO:140.2);ALT=G[chr11:65822542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65823057	+	chr11	65824308	+	.	2	8	4893650_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4893650_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_65807001_65832001_226C;SPAN=1251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:8 DR:2 LR:-12.96 LO:20.79);ALT=G[chr11:65824308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65824426	+	chr11	65825784	+	TAGCTGCTCCAGTGGGCCCAGTGGGCCCCACTCCTACAGTTTTGCCCATGGGAGCCCCTGTTCCCCGGCCTCGTGGTCCCCCACCGCCCCCTGGAGATGAGAACAGAGAGATGGATGACCCCTCTGTGGGCCCCAAGATCCCCCAGGCTTTGGAGAAGATCCTGCAGCTGAAGGAGAGCCGCCAGGAAGAGATGAATTCTCAGCAG	2	55	4893653_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TAGCTGCTCCAGTGGGCCCAGTGGGCCCCACTCCTACAGTTTTGCCCATGGGAGCCCCTGTTCCCCGGCCTCGTGGTCCCCCACCGCCCCCTGGAGATGAGAACAGAGAGATGGATGACCCCTCTGTGGGCCCCAAGATCCCCCAGGCTTTGGAGAAGATCCTGCAGCTGAAGGAGAGCCGCCAGGAAGAGATGAATTCTCAGCAG;MAPQ=60;MATEID=4893653_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_65807001_65832001_68C;SPAN=1358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:81 GQ:34.4 PL:[159.8, 0.0, 34.4] SR:55 DR:2 LR:-163.9 LO:163.9);ALT=G[chr11:65825784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65824470	+	chr11	65825522	+	.	10	0	4893654_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4893654_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:65824470(+)-11:65825522(-)__11_65807001_65832001D;SPAN=1052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.34 LO:20.42);ALT=G[chr11:65825522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65829469	+	chr11	65830478	+	.	2	9	4893670_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=4893670_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_65807001_65832001_272C;SPAN=1009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:84 GQ:10.4 PL:[10.4, 0.0, 191.9] SR:9 DR:2 LR:-10.25 LO:20.2);ALT=G[chr11:65830478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65829469	+	chr11	65830865	+	AGCTGTTCCTTTGGGTACCATGCTGGTGGCTGGGGCAAACCTCCAGTGGATGAGACTGGGAAACCGCTCTATGGGGACGTGTTTGGAACCAATGCTGCTGAA	5	20	4893671_1	46.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TTTCAG;INSERTION=AGCTGTTCCTTTGGGTACCATGCTGGTGGCTGGGGCAAACCTCCAGTGGATGAGACTGGGAAACCGCTCTATGGGGACGTGTTTGGAACCAATGCTGCTGAA;MAPQ=60;MATEID=4893671_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_65807001_65832001_272C;SPAN=1396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:86 GQ:46.1 PL:[46.1, 0.0, 161.6] SR:20 DR:5 LR:-46.02 LO:49.68);ALT=G[chr11:65830865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	65831200	+	chr11	65835416	+	.	0	12	4893878_1	26.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=4893878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_65831501_65856501_6C;SPAN=4216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:51 GQ:26 PL:[26.0, 0.0, 95.3] SR:12 DR:0 LR:-25.8 LO:28.16);ALT=G[chr11:65835416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66036199	+	chr11	66039626	+	.	13	0	4894643_1	20.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4894643_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66036199(+)-11:66039626(-)__11_66027501_66052501D;SPAN=3427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:85 GQ:20 PL:[20.0, 0.0, 185.0] SR:0 DR:13 LR:-19.88 LO:27.78);ALT=C[chr11:66039626[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66036203	+	chr11	66039835	+	.	13	0	4894645_1	22.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4894645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66036203(+)-11:66039835(-)__11_66027501_66052501D;SPAN=3632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:0 DR:13 LR:-22.32 LO:28.48);ALT=A[chr11:66039835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66109095	+	chr11	66112443	+	GGAGCTCTCCTCTTCTGACTCTGTCTGGCTGCCGCTCCGCTCCTCCTCACTCTCTTCCTCCTCCCCATTCATCTCAGCAGCAGAATCACCCTCTGCTTCCATCTCTTCTGTGTCTTTGCTTGGAGGCTGGACAGGCATCTGGACT	9	20	4894813_1	53.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGAGCTCTCCTCTTCTGACTCTGTCTGGCTGCCGCTCCGCTCCTCCTCACTCTCTTCCTCCTCCCCATTCATCTCAGCAGCAGAATCACCCTCTGCTTCCATCTCTTCTGTGTCTTTGCTTGGAGGCTGGACAGGCATCTGGACT;MAPQ=60;MATEID=4894813_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_66101001_66126001_10C;SPAN=3348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:73 GQ:53 PL:[53.0, 0.0, 122.3] SR:20 DR:9 LR:-52.84 LO:54.44);ALT=C[chr11:66112443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66109713	+	chr11	66112443	+	.	20	9	4894817_1	45.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4894817_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_66101001_66126001_10C;SPAN=2730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:102 GQ:45.2 PL:[45.2, 0.0, 200.3] SR:9 DR:20 LR:-44.99 LO:50.68);ALT=C[chr11:66112443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66204950	+	chr11	66206208	+	.	29	0	4895066_1	70.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4895066_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66204950(+)-11:66206208(-)__11_66199001_66224001D;SPAN=1258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:93 GQ:70.7 PL:[70.7, 0.0, 153.2] SR:0 DR:29 LR:-70.53 LO:72.28);ALT=C[chr11:66206208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66311452	+	chr11	66313194	+	.	11	12	4895353_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=4895353_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_66297001_66322001_125C;SPAN=1742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:96 GQ:36.8 PL:[36.8, 0.0, 195.2] SR:12 DR:11 LR:-36.71 LO:42.96);ALT=A[chr11:66313194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66360771	+	chr11	66366584	+	TTGGAGTTCGCGGTGCAGATGACCTGTCAGAGCTGTGTGGACGCGGTGCGCAAATCCCTGCAAGGGGTGG	77	103	4895588_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CAGGT;INSERTION=TTGGAGTTCGCGGTGCAGATGACCTGTCAGAGCTGTGTGGACGCGGTGCGCAAATCCCTGCAAGGGGTGG;MAPQ=60;MATEID=4895588_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_66346001_66371001_169C;SPAN=5813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:150 DP:115 GQ:40.6 PL:[445.6, 40.6, 0.0] SR:103 DR:77 LR:-445.6 LO:445.6);ALT=G[chr11:66366584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66711541	+	chr11	66713342	+	.	31	0	4896993_1	89.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=4896993_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66711541(+)-11:66713342(-)__11_66689001_66714001D;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=A[chr11:66713342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	66762769	-	chr11	66763925	+	.	9	0	4896903_1	19.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4896903_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:66762769(-)-11:66763925(-)__11_66738001_66763001D;SPAN=1156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:0 DR:9 LR:-19.68 LO:21.27);ALT=[chr11:66763925[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	67007840	+	chr11	67010478	+	.	5	6	4897828_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4897828_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_66983001_67008001_136C;SPAN=2638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:6 DR:5 LR:-15.57 LO:18.13);ALT=G[chr11:67010478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67167136	+	chr11	67168159	+	.	9	10	4898011_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4898011_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67154501_67179501_195C;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:72 GQ:30.2 PL:[30.2, 0.0, 142.4] SR:10 DR:9 LR:-30.01 LO:34.3);ALT=C[chr11:67168159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67209610	+	chr11	67210877	+	.	16	0	4898144_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4898144_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67209610(+)-11:67210877(-)__11_67203501_67228501D;SPAN=1267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:62 GQ:36.2 PL:[36.2, 0.0, 112.1] SR:0 DR:16 LR:-36.02 LO:38.3);ALT=G[chr11:67210877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67250729	+	chr11	67254475	+	.	40	24	4898541_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=4898541_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67252501_67277501_92C;SPAN=3746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:59 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:24 DR:40 LR:-174.9 LO:174.9);ALT=G[chr11:67254475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67254656	+	chr11	67256736	+	.	0	10	4898552_1	6.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4898552_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67252501_67277501_165C;SPAN=2080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:98 GQ:6.5 PL:[6.5, 0.0, 230.9] SR:10 DR:0 LR:-6.459 LO:19.48);ALT=G[chr11:67256736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67374547	+	chr11	67375866	+	.	75	30	4898795_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4898795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67350501_67375501_24C;SPAN=1319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:44 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:30 DR:75 LR:-254.2 LO:254.2);ALT=G[chr11:67375866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67415053	+	chr11	67418053	+	TATGGG	6	5	4898951_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACC;INSERTION=TATGGG;MAPQ=60;MATEID=4898951_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_11_67399501_67424501_395C;SPAN=3000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:5 DR:6 LR:0.1925 LO:12.92);ALT=T[chr11:67418053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67777863	+	chr11	67782764	+	.	21	4	4899753_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4899753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67767001_67792001_133C;SPAN=4901;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:88 GQ:52.1 PL:[52.1, 0.0, 161.0] SR:4 DR:21 LR:-52.08 LO:55.21);ALT=G[chr11:67782764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67782929	+	chr11	67785995	+	.	0	8	4899761_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4899761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67767001_67792001_274C;SPAN=3066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:8 DR:0 LR:-9.069 LO:16.34);ALT=G[chr11:67785995[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67798253	+	chr11	67800388	+	.	93	0	4900683_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4900683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67798253(+)-11:67800388(-)__11_67791501_67816501D;SPAN=2135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:89 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:93 LR:-274.0 LO:274.0);ALT=G[chr11:67800388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67798276	+	chr11	67799616	+	.	37	0	4900684_1	97.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4900684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67798276(+)-11:67799616(-)__11_67791501_67816501D;SPAN=1340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:91 GQ:97.7 PL:[97.7, 0.0, 120.8] SR:0 DR:37 LR:-97.48 LO:97.65);ALT=G[chr11:67799616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67800751	+	chr11	67803717	+	.	4	25	4900693_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=4900693_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67791501_67816501_196C;SPAN=2966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:124 GQ:62.3 PL:[62.3, 0.0, 237.2] SR:25 DR:4 LR:-62.13 LO:67.97);ALT=G[chr11:67803717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67806587	+	chr11	67808734	+	.	17	3	4900716_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4900716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67791501_67816501_89C;SPAN=2147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:61 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:3 DR:17 LR:-42.89 LO:44.34);ALT=G[chr11:67808734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67806614	+	chr11	67809219	+	.	14	0	4900717_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4900717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:67806614(+)-11:67809219(-)__11_67791501_67816501D;SPAN=2605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:50 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:0 DR:14 LR:-32.67 LO:34.1);ALT=G[chr11:67809219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	67957621	+	chr11	67980943	+	.	7	5	4900994_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4900994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_67963001_67988001_309C;SPAN=23322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:6 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:5 DR:7 LR:-26.41 LO:26.41);ALT=T[chr11:67980943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68580046	+	chr11	68582802	+	.	0	17	4903092_1	34.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4903092_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68575501_68600501_233C;SPAN=2756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:80 GQ:34.4 PL:[34.4, 0.0, 159.8] SR:17 DR:0 LR:-34.44 LO:39.04);ALT=T[chr11:68582802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68580089	+	chr11	68609245	+	.	10	0	4903093_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4903093_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68580089(+)-11:68609245(-)__11_68575501_68600501D;SPAN=29156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:0 DR:10 LR:-22.44 LO:23.91);ALT=C[chr11:68609245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68582956	+	chr11	68609241	+	.	35	6	4903104_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=4903104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68575501_68600501_141C;SPAN=26285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:29 GQ:9.9 PL:[108.9, 9.9, 0.0] SR:6 DR:35 LR:-108.9 LO:108.9);ALT=C[chr11:68609241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68605240	+	chr11	68609241	+	.	27	0	4902963_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4902963_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68605240(+)-11:68609241(-)__11_68600001_68625001D;SPAN=4001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:76 GQ:68.6 PL:[68.6, 0.0, 114.8] SR:0 DR:27 LR:-68.54 LO:69.2);ALT=A[chr11:68609241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68658863	+	chr11	68660358	+	.	2	45	4903512_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;MAPQ=60;MATEID=4903512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68649001_68674001_273C;SPAN=1495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:89 GQ:84.8 PL:[131.0, 0.0, 84.8] SR:45 DR:2 LR:-131.6 LO:131.6);ALT=A[chr11:68660358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68660462	+	chr11	68663981	+	CCTGCTGGTTGGGGCAGACAACTTCACGCTGCTTGGCAAGCCACTCCTCG	2	76	4903517_1	99.0	.	DISC_MAPQ=30;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CCTGCTGGTTGGGGCAGACAACTTCACGCTGCTTGGCAAGCCACTCCTCG;MAPQ=60;MATEID=4903517_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_68649001_68674001_213C;SPAN=3519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:96 GQ:0.5 PL:[231.5, 0.0, 0.5] SR:76 DR:2 LR:-245.5 LO:245.5);ALT=C[chr11:68663981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68664151	+	chr11	68665395	+	.	0	48	4903529_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTGCA;MAPQ=60;MATEID=4903529_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68649001_68674001_362C;SPAN=1244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:93 GQ:90.5 PL:[133.4, 0.0, 90.5] SR:48 DR:0 LR:-133.6 LO:133.6);ALT=A[chr11:68665395[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68664206	+	chr11	68671189	+	.	31	0	4903530_1	80.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4903530_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68664206(+)-11:68671189(-)__11_68649001_68674001D;SPAN=6983;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:79 GQ:80.9 PL:[80.9, 0.0, 110.6] SR:0 DR:31 LR:-80.93 LO:81.18);ALT=T[chr11:68671189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68665480	+	chr11	68668003	+	.	0	25	4903532_1	59.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4903532_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_68649001_68674001_326C;SPAN=2523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:84 GQ:59.9 PL:[59.9, 0.0, 142.4] SR:25 DR:0 LR:-59.77 LO:61.69);ALT=T[chr11:68668003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68665526	+	chr11	68671209	+	.	50	0	4903534_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4903534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68665526(+)-11:68671209(-)__11_68649001_68674001D;SPAN=5683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:82 GQ:53.9 PL:[143.0, 0.0, 53.9] SR:0 DR:50 LR:-144.9 LO:144.9);ALT=G[chr11:68671209[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68668115	+	chr11	68671220	+	.	15	0	4903539_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4903539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:68668115(+)-11:68671220(-)__11_68649001_68674001D;SPAN=3105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:84 GQ:26.9 PL:[26.9, 0.0, 175.4] SR:0 DR:15 LR:-26.76 LO:33.17);ALT=A[chr11:68671220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	68671508	+	chr11	68673534	+	.	6	3	4903547_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=4903547_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_11_68649001_68674001_379C;SPAN=2026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:81 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:3 DR:6 LR:-1.162 LO:13.11);ALT=T[chr11:68673534[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	33386451	+	chr11	76889255	+	GTGGACGGATGGATGGATGGATAGATGGGGGAA	10	31	4925704_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTGGACGGATGGATGGATGGATAGATGGGGGAA;MAPQ=60;MATEID=4925704_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_76881001_76906001_343C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:161 GQ:92 PL:[92.0, 0.0, 296.6] SR:31 DR:10 LR:-91.72 LO:97.87);ALT=]chr22:33386451]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	77103588	+	chr11	77122819	+	.	27	30	4926202_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4926202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77101501_77126501_105C;SPAN=19231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:97 GQ:99 PL:[125.6, 0.0, 109.1] SR:30 DR:27 LR:-125.6 LO:125.6);ALT=T[chr11:77122819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77333719	+	chr11	77336762	+	ATGTGCTTCCACATCATATTCTTCTCCATCGTAGTCATCTGAATCCTCATCCTCAGGATCTGGATGCAAGGCCTGGCATTCGCACATTGCAGTGAACATTGCCTCCA	2	14	4927173_1	26.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATGTGCTTCCACATCATATTCTTCTCCATCGTAGTCATCTGAATCCTCATCCTCAGGATCTGGATGCAAGGCCTGGCATTCGCACATTGCAGTGAACATTGCCTCCA;MAPQ=60;MATEID=4927173_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_77322001_77347001_57C;SPAN=3043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:99 GQ:26 PL:[26.0, 0.0, 214.1] SR:14 DR:2 LR:-25.99 LO:34.61);ALT=C[chr11:77336762[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77333719	+	chr11	77336008	+	.	4	7	4927172_1	12.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=4927172_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTG;SCTG=c_11_77322001_77347001_57C;SPAN=2289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:88 GQ:12.5 PL:[12.5, 0.0, 200.6] SR:7 DR:4 LR:-12.47 LO:22.46);ALT=C[chr11:77336008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77336865	+	chr11	77340808	+	.	0	35	4927183_1	90.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=4927183_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77322001_77347001_168C;SPAN=3943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:94 GQ:90.2 PL:[90.2, 0.0, 136.4] SR:35 DR:0 LR:-90.07 LO:90.62);ALT=T[chr11:77340808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77336903	+	chr11	77348655	+	.	13	0	4927235_1	23.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=4927235_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:77336903(+)-11:77348655(-)__11_77346501_77371501D;SPAN=11752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:71 GQ:23.9 PL:[23.9, 0.0, 146.0] SR:0 DR:13 LR:-23.68 LO:28.9);ALT=T[chr11:77348655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77340946	+	chr11	77348635	+	.	69	108	4927236_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4927236_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77346501_77371501_7C;SPAN=7689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:159 DP:52 GQ:43 PL:[472.0, 43.0, 0.0] SR:108 DR:69 LR:-472.0 LO:472.0);ALT=T[chr11:77348635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77475737	+	chr11	77531574	+	.	0	12	4927465_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CTT;MAPQ=60;MATEID=4927465_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77518001_77543001_48C;SPAN=55837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:40 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:12 DR:0 LR:-28.78 LO:29.66);ALT=T[chr11:77531574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77532287	+	chr11	77553524	+	.	37	5	4927615_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4927615_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77542501_77567501_219C;SPAN=21237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:36 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:5 DR:37 LR:-118.8 LO:118.8);ALT=G[chr11:77553524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77532317	+	chr11	77580765	+	.	8	0	4927544_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4927544_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:77532317(+)-11:77580765(-)__11_77567001_77592001D;SPAN=48448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=G[chr11:77580765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77781084	+	chr11	77784044	+	.	0	92	4928363_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4928363_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_77763001_77788001_42C;SPAN=2960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:101 GQ:27 PL:[297.0, 27.0, 0.0] SR:92 DR:0 LR:-297.1 LO:297.1);ALT=T[chr11:77784044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	77784239	+	chr11	77790677	+	.	39	0	4928397_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=4928397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:77784239(+)-11:77790677(-)__11_77787501_77812501D;SPAN=6438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:104 GQ:99 PL:[100.7, 0.0, 150.2] SR:0 DR:39 LR:-100.6 LO:101.1);ALT=T[chr11:77790677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	82536167	+	chr11	82549429	+	.	4	4	4938526_1	4.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4938526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_82540501_82565501_112C;SPAN=13262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:45 GQ:4.4 PL:[4.4, 0.0, 103.4] SR:4 DR:4 LR:-4.313 LO:9.938);ALT=G[chr11:82549429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	82571161	+	chr11	82611275	+	.	0	26	4938837_1	68.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=4938837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_82589501_82614501_132C;SPAN=40114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:66 GQ:68 PL:[68.0, 0.0, 91.1] SR:26 DR:0 LR:-67.95 LO:68.15);ALT=T[chr11:82611275[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	102213121	-	chr17	886817	+	.	6	17	6280789_1	26.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=TTTTTTTTTTTTTTGAGATGGAGT;MAPQ=60;MATEID=6280789_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=TTTTTTTTTTTTT;SCTG=c_17_882001_907001_11C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:22 DP:28 GQ:2.9 PL:[26.2, 2.9, 0.0] SR:17 DR:6 LR:-26.26 LO:26.26);ALT=[chr17:886817[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	102218107	+	chr11	102219328	+	.	6	5	4981917_1	8.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=4981917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_102214001_102239001_243C;SPAN=1221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:5 DR:6 LR:-8.577 LO:18.05);ALT=G[chr11:102219328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	102272991	+	chr11	102323277	+	.	14	0	4982527_1	33.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4982527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:102272991(+)-11:102323277(-)__11_102312001_102337001D;SPAN=50286;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:46 GQ:33.8 PL:[33.8, 0.0, 76.7] SR:0 DR:14 LR:-33.75 LO:34.71);ALT=T[chr11:102323277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	102319649	+	chr11	102323349	+	.	17	0	4982542_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4982542_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:102319649(+)-11:102323349(-)__11_102312001_102337001D;SPAN=3700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:63 GQ:39.2 PL:[39.2, 0.0, 111.8] SR:0 DR:17 LR:-39.05 LO:41.08);ALT=T[chr11:102323349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	105948621	+	chr11	105950193	+	.	8	13	4990149_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=4990149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_105938001_105963001_103C;SPAN=1572;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:73 GQ:36.5 PL:[36.5, 0.0, 138.8] SR:13 DR:8 LR:-36.34 LO:39.81);ALT=G[chr11:105950193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	106044581	+	chr19	49290023	+	.	8	48	6846481_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6846481_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_49269501_49294501_217C;SECONDARY;SPAN=-1;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:57 GQ:8.7 PL:[155.1, 8.7, 0.0] SR:48 DR:8 LR:-157.7 LO:157.7);ALT=A[chr19:49290023[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr11	111750349	+	chr11	111753087	+	.	34	0	5004468_1	90.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5004468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:111750349(+)-11:111753087(-)__11_111744501_111769501D;SPAN=2738;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:79 GQ:90.8 PL:[90.8, 0.0, 100.7] SR:0 DR:34 LR:-90.83 LO:90.86);ALT=T[chr11:111753087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111753322	+	chr11	111754495	+	TTTGGACACTACTTTGAAACAACATATGATACAAGCTACAACAACAAAATGCCACTTTCAACACATA	0	10	5004477_1	11.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTGGACACTACTTTGAAACAACATATGATACAAGCTACAACAACAAAATGCCACTTTCAACACATA;MAPQ=60;MATEID=5004477_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_111744501_111769501_262C;SPAN=1173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:10 DR:0 LR:-10.79 LO:20.31);ALT=G[chr11:111754495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111949039	+	chr11	111951131	+	.	0	11	5004888_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5004888_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_11_111940501_111965501_328C;SPAN=2092;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:11 DR:0 LR:-16.53 LO:23.43);ALT=G[chr11:111951131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111956197	+	chr11	111957359	+	.	67	0	5004916_1	99.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5004916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:111956197(+)-11:111957359(-)__11_111940501_111965501D;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:77 GQ:14.1 PL:[214.5, 14.1, 0.0] SR:0 DR:67 LR:-216.8 LO:216.8);ALT=A[chr11:111957359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	111957397	-	chrX	133300749	+	.	13	0	7530027_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7530027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:111957397(-)-23:133300749(-)__23_133280001_133305001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:0 DR:13 LR:-33.7 LO:33.85);ALT=[chrX:133300749[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	112020930	+	chr11	112025698	+	ATCATCTTCAG	0	30	5005066_1	75.0	.	EVDNC=ASSMB;INSERTION=ATCATCTTCAG;MAPQ=60;MATEID=5005066_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_112014001_112039001_256C;SPAN=4768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:87 GQ:75.5 PL:[75.5, 0.0, 134.9] SR:30 DR:0 LR:-75.46 LO:76.4);ALT=C[chr11:112025698[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	112020987	+	chr11	112034627	+	.	15	0	5005067_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5005067_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:112020987(+)-11:112034627(-)__11_112014001_112039001D;SPAN=13640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:82 GQ:27.5 PL:[27.5, 0.0, 169.4] SR:0 DR:15 LR:-27.3 LO:33.34);ALT=T[chr11:112034627[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	112025808	+	chr11	112034629	+	.	55	20	5005082_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=5005082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_112014001_112039001_261C;SPAN=8821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:81 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:20 DR:55 LR:-235.6 LO:235.6);ALT=G[chr11:112034629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	112258722	-	chr16	30763574	+	.	12	0	6185727_1	34.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6185727_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:112258722(-)-16:30763574(-)__16_30747501_30772501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:21 GQ:14.3 PL:[34.1, 0.0, 14.3] SR:0 DR:12 LR:-34.22 LO:34.22);ALT=[chr16:30763574[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr22	39916657	+	chr11	113660903	+	.	23	0	7300416_1	61.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=7300416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:113660903(-)-22:39916657(+)__22_39910501_39935501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:54 GQ:61.4 PL:[61.4, 0.0, 68.0] SR:0 DR:23 LR:-61.29 LO:61.32);ALT=]chr22:39916657]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	114310435	+	chr11	114314577	+	.	8	0	5010770_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5010770_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:114310435(+)-11:114314577(-)__11_114292501_114317501D;SPAN=4142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:0 DR:8 LR:2.581 LO:14.46);ALT=A[chr11:114314577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	114311462	+	chr11	114315261	+	GTCCTAACCTGATTATAAAACAACCAGATGAGTTGCTGGACAGCATGTCAGATTGGTGTAAGGAGCATCACGGGA	0	16	5010774_1	28.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GTCCTAACCTGATTATAAAACAACCAGATGAGTTGCTGGACAGCATGTCAGATTGGTGTAAGGAGCATCACGGGA;MAPQ=60;MATEID=5010774_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_114292501_114317501_112C;SPAN=3799;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:91 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:16 DR:0 LR:-28.16 LO:35.26);ALT=G[chr11:114315261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	121498477	+	chr11	121500204	+	.	2	8	5029693_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5029693_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_121495501_121520501_27C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:8 DR:2 LR:-3.971 LO:17.23);ALT=G[chr11:121500204[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	122347584	+	chr11	122349281	+	.	79	60	5031365_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAGAAAG;MAPQ=60;MATEID=5031365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_122328501_122353501_261C;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:42 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:60 DR:79 LR:-346.6 LO:346.6);ALT=G[chr11:122349281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	122931522	+	chr11	122932783	+	.	51	0	5033502_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5033502_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:122931522(+)-11:122932783(-)__11_122916501_122941501D;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:224 GQ:99 PL:[107.8, 0.0, 434.6] SR:0 DR:51 LR:-107.7 LO:118.9);ALT=A[chr11:122932783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124493130	+	chr11	124495565	+	AAAATGCTGCTATTTGTGATGAAATTGCTCGTCTTGAGGAAAAATTTCTTAAAGCAAAAGAAGAAAGA	2	13	5036918_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGGT;INSERTION=AAAATGCTGCTATTTGTGATGAAATTGCTCGTCTTGAGGAAAAATTTCTTAAAGCAAAAGAAGAAAGA;MAPQ=60;MATEID=5036918_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_124484501_124509501_206C;SPAN=2435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:13 DR:2 LR:-26.49 LO:33.08);ALT=G[chr11:124495565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124609932	+	chr11	124615397	+	.	9	0	5037214_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5037214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:124609932(+)-11:124615397(-)__11_124607001_124632001D;SPAN=5465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:0 DR:9 LR:-11.83 LO:18.75);ALT=C[chr11:124615397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124971332	+	chr11	124981440	+	.	10	0	5038162_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5038162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:124971332(+)-11:124981440(-)__11_124974501_124999501D;SPAN=10108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:0 DR:10 LR:-20.55 LO:23.07);ALT=T[chr11:124981440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124972477	+	chr11	124981433	+	.	17	0	5038163_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5038163_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:124972477(+)-11:124981433(-)__11_124974501_124999501D;SPAN=8956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:0 DR:17 LR:-44.2 LO:44.37);ALT=C[chr11:124981433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	124972732	+	chr11	124981433	+	.	9	0	5038164_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5038164_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:124972732(+)-11:124981433(-)__11_124974501_124999501D;SPAN=8701;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=A[chr11:124981433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	125439469	+	chr11	125442353	+	.	13	9	5039416_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5039416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_125440001_125465001_367C;SPAN=2884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:38 GQ:32.6 PL:[32.6, 0.0, 59.0] SR:9 DR:13 LR:-32.62 LO:33.05);ALT=G[chr11:125442353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	125439484	+	chr11	125445158	+	.	8	0	5039417_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5039417_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:125439484(+)-11:125445158(-)__11_125440001_125465001D;SPAN=5674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:32 GQ:17.9 PL:[17.9, 0.0, 57.5] SR:0 DR:8 LR:-17.74 LO:19.02);ALT=A[chr11:125445158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	125465898	+	chr11	125472198	+	CCTTCTCCACTCGTCTGTTTGCTGTCCTGAGATTTGAAAGTGTTATCCATGAGTTTGATCC	0	17	5039500_1	40.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=CCTTCTCCACTCGTCTGTTTGCTGTCCTGAGATTTGAAAGTGTTATCCATGAGTTTGATCC;MAPQ=60;MATEID=5039500_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_11_125464501_125489501_212C;SPAN=6300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:58 GQ:40.4 PL:[40.4, 0.0, 99.8] SR:17 DR:0 LR:-40.4 LO:41.81);ALT=T[chr11:125472198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	125484148	+	chr11	125488266	+	.	8	0	5039556_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5039556_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:125484148(+)-11:125488266(-)__11_125464501_125489501D;SPAN=4118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:0 DR:8 LR:-3.921 LO:15.38);ALT=G[chr11:125488266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	125937458	-	chr12	76478348	+	.	17	0	5252423_1	42.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=5252423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:125937458(-)-12:76478348(-)__12_76464501_76489501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:0 DR:17 LR:-42.84 LO:43.35);ALT=[chr12:76478348[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr11	126117274	-	chr11	126118391	+	.	17	0	5041198_1	34.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=5041198_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:126117274(-)-11:126118391(-)__11_126101501_126126501D;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:79 GQ:34.7 PL:[34.7, 0.0, 156.8] SR:0 DR:17 LR:-34.71 LO:39.14);ALT=[chr11:126118391[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr11	126139186	+	chr11	126141331	+	.	7	3	5041324_1	2.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5041324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_126126001_126151001_14C;SPAN=2145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:3 DR:7 LR:-2.567 LO:15.16);ALT=G[chr11:126141331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	126174178	+	chr11	126176463	+	.	0	13	5041434_1	32.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5041434_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_11_126150501_126175501_280C;SPAN=2285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:41 GQ:32 PL:[32.0, 0.0, 65.0] SR:13 DR:0 LR:-31.81 LO:32.52);ALT=T[chr11:126176463[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	126212228	+	chr11	126225354	+	.	8	0	5041557_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5041557_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:126212228(+)-11:126225354(-)__11_126199501_126224501D;SPAN=13126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=G[chr11:126225354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	126225720	+	chr11	126276367	+	.	10	0	5041670_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5041670_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:126225720(+)-11:126276367(-)__11_126273001_126298001D;SPAN=50647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=C[chr11:126276367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr11	126225740	+	chr11	126275990	+	.	18	12	5041671_1	58.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=5041671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_126273001_126298001_113C;SPAN=50250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:39 GQ:35.6 PL:[58.7, 0.0, 35.6] SR:12 DR:18 LR:-59.05 LO:59.05);ALT=G[chr11:126275990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29447481	+	chr12	145759	+	.	26	0	6362896_1	73.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6362896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:145759(-)-17:29447481(+)__17_29424501_29449501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:47 GQ:40.1 PL:[73.1, 0.0, 40.1] SR:0 DR:26 LR:-73.58 LO:73.58);ALT=]chr17:29447481]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	394830	+	chr12	401923	+	.	5	4	5062912_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5062912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_392001_417001_178C;SPAN=7093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:4 DR:5 LR:-5.818 LO:15.7);ALT=T[chr12:401923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	417172	+	chr12	418967	+	.	3	3	5062980_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=5062980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_416501_441501_27C;SPAN=1795;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:99 GQ:13.5 PL:[0.0, 13.5, 267.3] SR:3 DR:3 LR:13.62 LO:6.133);ALT=C[chr12:418967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	653462	-	chr12	654763	+	CCTCCACACCTCG	4	10	5063818_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCTCCACACCTCG;MAPQ=60;MATEID=5063818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_637001_662001_287C;SPAN=1301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:125 GQ:12.5 PL:[12.5, 0.0, 289.7] SR:10 DR:4 LR:-12.35 LO:27.88);ALT=[chr12:654763[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	653642	+	chr12	654821	-	.	2	6	5063822_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5063822_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_637001_662001_313C;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:124 GQ:6.9 PL:[0.0, 6.9, 313.5] SR:6 DR:2 LR:7.187 LO:13.93);ALT=T]chr12:654821];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	675355	+	chr12	752733	+	.	8	0	5064171_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5064171_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:675355(+)-12:752733(-)__12_735001_760001D;SPAN=77378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:33 GQ:17.6 PL:[17.6, 0.0, 60.5] SR:0 DR:8 LR:-17.47 LO:18.9);ALT=G[chr12:752733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	1857701	+	chr12	785370	+	.	19	44	5064871_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TGGCTCA;MAPQ=60;MATEID=5064871_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_784001_809001_356C;SPAN=1072331;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:28 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:44 DR:19 LR:-174.9 LO:174.9);ALT=]chr12:1857701]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	1194568	+	chr12	1199981	+	.	15	0	5065864_1	39.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=5065864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:1194568(+)-12:1199981(-)__12_1176001_1201001D;SPAN=5413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:38 GQ:39.2 PL:[39.2, 0.0, 52.4] SR:0 DR:15 LR:-39.22 LO:39.33);ALT=G[chr12:1199981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	1195045	+	chr12	1200053	+	.	10	0	5065867_1	25.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=5065867_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:1195045(+)-12:1200053(-)__12_1176001_1201001D;SPAN=5008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:28 GQ:25.4 PL:[25.4, 0.0, 41.9] SR:0 DR:10 LR:-25.42 LO:25.66);ALT=G[chr12:1200053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	1800380	+	chr12	1863423	+	.	11	4	5067817_1	27.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5067817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_1862001_1887001_370C;SPAN=63043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:4 DR:11 LR:-27.42 LO:28.93);ALT=G[chr12:1863423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6041904	+	chr12	6040782	+	.	58	0	5078888_1	99.0	.	DISC_MAPQ=6;EVDNC=DSCRD;IMPRECISE;MAPQ=6;MATEID=5078888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6040782(-)-12:6041904(+)__12_6027001_6052001D;SPAN=1122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:200 GQ:99 PL:[137.3, 0.0, 348.5] SR:0 DR:58 LR:-137.3 LO:142.3);ALT=]chr12:6041904]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	6241438	+	chr12	6248078	+	.	40	49	5079389_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5079389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6247501_6272501_101C;SPAN=6640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:30 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:49 DR:40 LR:-211.3 LO:211.3);ALT=G[chr12:6248078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6309729	+	chr12	6341794	+	.	12	0	5079337_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5079337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6309729(+)-12:6341794(-)__12_6296501_6321501D;SPAN=32065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=T[chr12:6341794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6309731	+	chr12	6334591	+	.	56	58	5079338_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5079338_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6296501_6321501_150C;SPAN=24860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:44 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:58 DR:56 LR:-267.4 LO:267.4);ALT=G[chr12:6334591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6334701	+	chr12	6341795	+	.	0	29	5079275_1	71.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=5079275_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6321001_6346001_6C;SPAN=7094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:92 GQ:71 PL:[71.0, 0.0, 150.2] SR:29 DR:0 LR:-70.8 LO:72.45);ALT=G[chr12:6341795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6345441	+	chr12	6346928	+	.	5	10	5079583_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5079583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6345501_6370501_331C;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:58 GQ:30.5 PL:[30.5, 0.0, 109.7] SR:10 DR:5 LR:-30.5 LO:33.04);ALT=G[chr12:6346928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6443411	+	chr12	6450946	+	AGC	0	12	5079901_1	29.0	.	EVDNC=ASSMB;INSERTION=AGC;MAPQ=60;MATEID=5079901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6419001_6444001_156C;SPAN=7535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:36 GQ:29.9 PL:[29.9, 0.0, 56.3] SR:12 DR:0 LR:-29.86 LO:30.34);ALT=C[chr12:6450946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6547703	-	chr15	40331293	+	.	116	0	5930665_1	99.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=5930665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6547703(-)-15:40331293(-)__15_40327001_40352001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:70 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:0 DR:116 LR:-343.3 LO:343.3);ALT=[chr15:40331293[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	6557359	+	chr12	6560633	+	.	8	0	5080154_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5080154_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6557359(+)-12:6560633(-)__12_6541501_6566501D;SPAN=3274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=A[chr12:6560633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6570104	+	chr12	6571198	+	.	0	6	5080035_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5080035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6566001_6591001_56C;SPAN=1094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:115 GQ:11.1 PL:[0.0, 11.1, 300.3] SR:6 DR:0 LR:11.35 LO:9.877);ALT=G[chr12:6571198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6644055	+	chr12	6645657	+	.	80	0	5080809_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5080809_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6644055(+)-12:6645657(-)__12_6639501_6664501D;SPAN=1602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:80 DP:119 GQ:56.9 PL:[231.8, 0.0, 56.9] SR:0 DR:80 LR:-237.8 LO:237.8);ALT=T[chr12:6645657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6682437	+	chr12	6686951	+	.	3	5	5080745_1	0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5080745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6664001_6689001_298C;SPAN=4514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:5 DR:3 LR:-0.6203 LO:13.03);ALT=T[chr12:6686951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6711665	+	chr12	6715440	+	.	2	8	5081036_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5081036_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_6688501_6713501_87C;SPAN=3775;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:52 GQ:15.8 PL:[15.8, 0.0, 108.2] SR:8 DR:2 LR:-15.62 LO:19.77);ALT=T[chr12:6715440[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6762600	+	chr12	6772227	+	.	31	0	5081197_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5081197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:6762600(+)-12:6772227(-)__12_6737501_6762501D;SPAN=9627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:1 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:31 LR:-89.12 LO:89.12);ALT=G[chr12:6772227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	6859472	+	chr12	6861090	+	ATGTTTCCAATCATGTCATTCATCATCCCAAACATGTCCATGAAACCACCCGACATTCCCAGCATCCCAAAGGGGGAGACAGCTCCAG	6	18	5081538_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=ATGTTTCCAATCATGTCATTCATCATCCCAAACATGTCCATGAAACCACCCGACATTCCCAGCATCCCAAAGGGGGAGACAGCTCCAG;MAPQ=60;MATEID=5081538_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_6860001_6885001_99C;SPAN=1618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:45 GQ:50.6 PL:[57.2, 0.0, 50.6] SR:18 DR:6 LR:-57.14 LO:57.14);ALT=C[chr12:6861090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	7053818	+	chr12	7054932	+	.	18	43	5081934_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=5081934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_7031501_7056501_293C;SPAN=1114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:115 GQ:99 PL:[147.2, 0.0, 130.7] SR:43 DR:18 LR:-147.1 LO:147.1);ALT=G[chr12:7054932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	7075664	+	chr12	7076839	+	GTCTTGGAGATATTCTGGGCTGCTCGAATCTTGCGAAGTTTGATGTAGCCAGGGTTCTTGCTCAGTGCTTCTCCAAG	0	13	5082553_1	22.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTCTTGGAGATATTCTGGGCTGCTCGAATCTTGCGAAGTTTGATGTAGCCAGGGTTCTTGCTCAGTGCTTCTCCAAG;MAPQ=60;MATEID=5082553_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_7056001_7081001_35C;SPAN=1175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:13 DR:0 LR:-22.32 LO:28.48);ALT=C[chr12:7076839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	7080257	+	chr12	7083499	+	.	20	16	5082573_1	64.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTAG;MAPQ=60;MATEID=5082573_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_12_7056001_7081001_87C;SPAN=3242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:44 GQ:41 PL:[64.1, 0.0, 41.0] SR:16 DR:20 LR:-64.23 LO:64.23);ALT=G[chr12:7083499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	7092701	+	chr12	7125576	+	.	0	9	5082593_1	17.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=5082593_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_7105001_7130001_345C;SPAN=32875;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:9 DR:0 LR:-17.79 LO:20.5);ALT=C[chr12:7125576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	7830042	-	chr18	44021851	+	GGGCC	29	36	6610257_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=GGGCC;MAPQ=60;MATEID=6610257_2;MATENM=5;NM=1;NUMPARTS=2;SCTG=c_18_44002001_44027001_84C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:42 GQ:15 PL:[165.0, 15.0, 0.0] SR:36 DR:29 LR:-165.0 LO:165.0);ALT=[chr18:44021851[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	8085795	+	chr12	8088616	+	.	23	0	5085528_1	51.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5085528_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:8085795(+)-12:8088616(-)__12_8085001_8110001D;SPAN=2821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:89 GQ:51.8 PL:[51.8, 0.0, 164.0] SR:0 DR:23 LR:-51.81 LO:55.07);ALT=A[chr12:8088616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	8086500	+	chr12	8088614	+	.	0	31	5085529_1	77.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=57;MATEID=5085529_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_8085001_8110001_2C;SPAN=2114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:94 GQ:77 PL:[77.0, 0.0, 149.6] SR:31 DR:0 LR:-76.86 LO:78.2);ALT=T[chr12:8088614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	8234980	+	chr12	8242530	+	.	12	4	5086009_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5086009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_8232001_8257001_238C;SPAN=7550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:119 GQ:10.7 PL:[10.7, 0.0, 278.0] SR:4 DR:12 LR:-10.67 LO:25.74);ALT=G[chr12:8242530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	8276589	+	chr12	8281859	+	.	9	0	5086163_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5086163_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:8276589(+)-12:8281859(-)__12_8281001_8306001D;SPAN=5270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:0 DR:9 LR:-20.77 LO:21.8);ALT=G[chr12:8281859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9099001	+	chr12	9102083	+	.	0	43	5088552_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5088552_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9089501_9114501_32C;SPAN=3082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:94 GQ:99 PL:[116.6, 0.0, 110.0] SR:43 DR:0 LR:-116.5 LO:116.5);ALT=C[chr12:9102083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9144907	+	chr12	9147714	+	.	9	5	5088859_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5088859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9138501_9163501_18C;SPAN=2807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:81 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:5 DR:9 LR:-20.97 LO:28.08);ALT=G[chr12:9147714[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9632740	+	chr12	31353916	-	.	12	0	5143589_1	28.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=5143589_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:9632740(+)-12:31353916(+)__12_31335501_31360501D;SPAN=21721176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:41 GQ:28.7 PL:[28.7, 0.0, 68.3] SR:0 DR:12 LR:-28.5 LO:29.51);ALT=C]chr12:31353916];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	9697953	+	chr12	31298444	-	.	2	5	5090337_1	9.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=32;MATEID=5090337_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9677501_9702501_18C;SPAN=21600491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:37 GQ:9.8 PL:[9.8, 0.0, 79.1] SR:5 DR:2 LR:-9.782 LO:12.99);ALT=G]chr12:31298444];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	9801529	+	chr12	9806276	+	.	11	27	5090613_1	82.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=5090613_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9800001_9825001_19C;SPAN=4747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:87 GQ:82.1 PL:[82.1, 0.0, 128.3] SR:27 DR:11 LR:-82.06 LO:82.64);ALT=G[chr12:9806276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9906186	+	chr12	9907658	+	AGTTGTTAAATTCTTTGCCATTTGACCACTTCCATGGGTGACCAGGTTCCTTTTTCAGTCCAACCCAGTGTTCCTCTCTACCTGCGTATCGTTTTAGAAAGTT	0	25	5090930_1	55.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGTTGTTAAATTCTTTGCCATTTGACCACTTCCATGGGTGACCAGGTTCCTTTTTCAGTCCAACCCAGTGTTCCTCTCTACCTGCGTATCGTTTTAGAAAGTT;MAPQ=60;MATEID=5090930_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_9898001_9923001_234C;SPAN=1472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:100 GQ:55.4 PL:[55.4, 0.0, 187.4] SR:25 DR:0 LR:-55.43 LO:59.44);ALT=C[chr12:9907658[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9906387	+	chr12	9907513	+	.	11	0	5090932_1	19.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5090932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:9906387(+)-12:9907513(-)__12_9898001_9923001D;SPAN=1126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:64 GQ:19.1 PL:[19.1, 0.0, 134.6] SR:0 DR:11 LR:-18.97 LO:24.12);ALT=A[chr12:9907513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9907908	+	chr12	9913431	+	.	73	0	5090940_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5090940_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:9907908(+)-12:9913431(-)__12_9898001_9923001D;SPAN=5523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:159 GQ:99 PL:[197.9, 0.0, 188.0] SR:0 DR:73 LR:-197.9 LO:197.9);ALT=A[chr12:9913431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	9909015	+	chr12	9913353	+	.	111	36	5090943_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5090943_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TACTAC;SCTG=c_12_9898001_9923001_218C;SPAN=4338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:119 DP:166 GQ:33.3 PL:[264.8, 0.0, 33.3] SR:36 DR:111 LR:-276.8 LO:276.8);ALT=T[chr12:9913353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10007084	+	chr12	10010073	+	.	0	11	5091104_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5091104_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9996001_10021001_261C;SPAN=2989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:82 GQ:14.3 PL:[14.3, 0.0, 182.6] SR:11 DR:0 LR:-14.1 LO:22.83);ALT=C[chr12:10010073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10007132	+	chr12	10021883	+	.	19	0	5091217_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5091217_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:10007132(+)-12:10021883(-)__12_10020501_10045501D;SPAN=14751;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:55 GQ:47.9 PL:[47.9, 0.0, 84.2] SR:0 DR:19 LR:-47.82 LO:48.41);ALT=C[chr12:10021883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10010238	+	chr12	10015098	+	.	2	77	5091116_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5091116_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_9996001_10021001_170C;SPAN=4860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:111 GQ:36.2 PL:[230.9, 0.0, 36.2] SR:77 DR:2 LR:-238.5 LO:238.5);ALT=T[chr12:10015098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10010572	+	chr12	10021800	+	.	84	0	5091219_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5091219_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:10010572(+)-12:10021800(-)__12_10020501_10045501D;SPAN=11228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:53 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=A[chr12:10021800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10015173	+	chr12	10021801	+	.	0	53	5091220_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TACC;MAPQ=60;MATEID=5091220_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_10020501_10045501_10C;SPAN=6628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:53 DR:0 LR:-158.4 LO:158.4);ALT=C[chr12:10021801[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10124286	+	chr12	10131563	+	.	34	46	5091603_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5091603_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_10118501_10143501_313C;SPAN=7277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:91 GQ:54.8 PL:[163.7, 0.0, 54.8] SR:46 DR:34 LR:-166.3 LO:166.3);ALT=G[chr12:10131563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10124286	+	chr12	10131935	+	CACCTCCAGCTCCCTCTCATGTATGGCGTCCAGCAGCCTTGTTTCTGACTCTTCTGTGCCTTCTGTTGCTCATTGGATTGGGAGTCTTGGCAAGCATGT	11	60	5091604_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CACCTCCAGCTCCCTCTCATGTATGGCGTCCAGCAGCCTTGTTTCTGACTCTTCTGTGCCTTCTGTTGCTCATTGGATTGGGAGTCTTGGCAAGCATGT;MAPQ=60;MATEID=5091604_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_10118501_10143501_313C;SPAN=7649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:106 GQ:63.8 PL:[192.5, 0.0, 63.8] SR:60 DR:11 LR:-195.9 LO:195.9);ALT=G[chr12:10131935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10133333	+	chr12	10134618	+	.	2	3	5091628_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5091628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_10118501_10143501_221C;SPAN=1285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:80 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:3 DR:2 LR:5.169 LO:8.632);ALT=G[chr12:10134618[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10280446	+	chr12	10282578	+	.	0	7	5091686_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5091686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_10265501_10290501_70C;SPAN=2132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:7 DR:0 LR:1.818 LO:12.7);ALT=T[chr12:10282578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10760537	+	chr12	10763220	+	CTTATGTGCACAAGAGTGTAATGGAAGAACTGAAGAGAATTATTGATGACAGTGAAATTACAAAAGAAGATGATGCTTTGTGGCCTCCCCCTGATAGGGTTGGCCGAC	0	33	5093200_1	91.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTTATGTGCACAAGAGTGTAATGGAAGAACTGAAGAGAATTATTGATGACAGTGAAATTACAAAAGAAGATGATGCTTTGTGGCCTCCCCCTGATAGGGTTGGCCGAC;MAPQ=60;MATEID=5093200_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_12_10755501_10780501_22C;SPAN=2683;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:65 GQ:65 PL:[91.4, 0.0, 65.0] SR:33 DR:0 LR:-91.53 LO:91.53);ALT=T[chr12:10763220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	10762589	+	chr12	10766036	+	.	11	0	5093207_1	11.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=5093207_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:10762589(+)-12:10766036(-)__12_10755501_10780501D;SPAN=3447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:91 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:0 DR:11 LR:-11.66 LO:22.29);ALT=C[chr12:10766036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	11192447	+	chr12	11218062	+	.	17	21	5094374_1	89.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=CTC;MAPQ=60;MATEID=5094374_2;MATENM=6;NM=2;NUMPARTS=2;SCTG=c_12_11172001_11197001_312C;SPAN=25615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:37 GQ:0 PL:[89.1, 0.0, 0.0] SR:21 DR:17 LR:-94.35 LO:94.35);ALT=C[chr12:11218062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	11199789	+	chr12	11324019	+	.	17	13	5094461_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5094461_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_11319001_11344001_253C;SPAN=124230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:83 GQ:47 PL:[47.0, 0.0, 152.6] SR:13 DR:17 LR:-46.83 LO:50.06);ALT=T[chr12:11324019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	11803094	+	chr12	11905382	+	.	0	7	5095814_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5095814_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_11882501_11907501_139C;SPAN=102288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:47 GQ:10.4 PL:[10.4, 0.0, 102.8] SR:7 DR:0 LR:-10.37 LO:14.87);ALT=G[chr12:11905382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	12022903	+	chr12	12037377	+	.	3	3	5096218_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5096218_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_12029501_12054501_341C;SPAN=14474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:36 GQ:6.8 PL:[6.8, 0.0, 79.4] SR:3 DR:3 LR:-6.752 LO:10.46);ALT=G[chr12:12037377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	12037521	+	chr12	12038858	+	.	2	3	5096241_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5096241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_12029501_12054501_106C;SPAN=1337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:86 GQ:9.9 PL:[0.0, 9.9, 227.7] SR:3 DR:2 LR:10.1 LO:6.381);ALT=G[chr12:12038858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	12544867	+	chr12	12546626	-	.	44	0	5097666_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5097666_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:12544867(+)-12:12546626(+)__12_12519501_12544501D;SPAN=1759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:0 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:0 DR:44 LR:-128.7 LO:128.7);ALT=C]chr12:12546626];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	12871888	+	chr12	12873969	+	.	3	3	5098882_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5098882_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_12862501_12887501_200C;SPAN=2081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:76 GQ:3.9 PL:[0.0, 3.9, 191.4] SR:3 DR:3 LR:4.085 LO:8.747);ALT=G[chr12:12873969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	12966378	+	chr12	12974139	+	.	10	0	5099029_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5099029_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:12966378(+)-12:12974139(-)__12_12960501_12985501D;SPAN=7761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:0 DR:10 LR:-10.79 LO:20.31);ALT=T[chr12:12974139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	13140267	+	chr12	13142210	+	.	4	7	5099715_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5099715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_13132001_13157001_328C;SPAN=1943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:7 DR:4 LR:-4.784 LO:17.36);ALT=C[chr12:13142210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	13142351	+	chr12	13152970	+	.	0	25	5099722_1	56.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5099722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_13132001_13157001_140C;SPAN=10619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:98 GQ:56 PL:[56.0, 0.0, 181.4] SR:25 DR:0 LR:-55.97 LO:59.7);ALT=T[chr12:13152970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48548230	+	chr12	13577390	+	.	3	5	6843159_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGG;MAPQ=60;MATEID=6843159_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48534501_48559501_105C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:55 GQ:1.7 PL:[1.7, 0.0, 130.4] SR:5 DR:3 LR:-1.604 LO:9.478);ALT=]chr19:48548230]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	21654882	+	chr12	21659819	+	.	17	16	5119749_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5119749_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_21633501_21658501_62C;SPAN=4937;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:47 GQ:50 PL:[63.2, 0.0, 50.0] SR:16 DR:17 LR:-63.26 LO:63.26);ALT=A[chr12:21659819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21659912	+	chr12	21661317	+	.	0	7	5119649_1	4.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=5119649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_21658001_21683001_277C;SPAN=1405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:71 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:7 DR:0 LR:-3.871 LO:13.53);ALT=T[chr12:21661317[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21791405	+	chr12	21794886	+	.	13	21	5120072_1	74.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5120072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_21780501_21805501_148C;SPAN=3481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:90 GQ:74.6 PL:[74.6, 0.0, 143.9] SR:21 DR:13 LR:-74.65 LO:75.85);ALT=C[chr12:21794886[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21795061	+	chr12	21796869	+	.	11	30	5120082_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5120082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_21780501_21805501_70C;SPAN=1808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:83 GQ:96.5 PL:[103.1, 0.0, 96.5] SR:30 DR:11 LR:-103.0 LO:103.0);ALT=T[chr12:21796869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21797047	+	chr12	21799833	+	.	7	82	5120086_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTTTA;MAPQ=60;MATEID=5120086_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_21780501_21805501_197C;SPAN=2786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:98 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:82 DR:7 LR:-289.9 LO:289.9);ALT=A[chr12:21799833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21797088	+	chr12	21810684	+	.	28	0	5120203_1	71.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5120203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:21797088(+)-12:21810684(-)__12_21805001_21830001D;SPAN=13596;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:77 GQ:71.6 PL:[71.6, 0.0, 114.5] SR:0 DR:28 LR:-71.57 LO:72.13);ALT=A[chr12:21810684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21800002	+	chr12	21810684	+	.	103	0	5120205_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5120205_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:21800002(+)-12:21810684(-)__12_21805001_21830001D;SPAN=10682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:77 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:0 DR:103 LR:-303.7 LO:303.7);ALT=A[chr12:21810684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	21807612	+	chr12	21810685	+	.	132	33	5120215_1	99.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=C;MAPQ=56;MATEID=5120215_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_21805001_21830001_23C;SPAN=3073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:161 DP:131 GQ:43.3 PL:[475.3, 43.3, 0.0] SR:33 DR:132 LR:-475.3 LO:475.3);ALT=C[chr12:21810685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	45143512	+	chr12	22538398	+	.	17	0	5122025_1	52.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5122025_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:22538398(-)-13:45143512(+)__12_22515501_22540501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:17 DP:20 GQ:2.1 PL:[52.8, 2.1, 0.0] SR:0 DR:17 LR:-54.44 LO:54.44);ALT=]chr13:45143512]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	23720523	-	chr12	23721695	+	.	8	0	5124655_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5124655_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:23720523(-)-12:23721695(-)__12_23716001_23741001D;SPAN=1172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=[chr12:23721695[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	25348332	+	chr12	25356854	+	AAA	3	10	5128831_1	24.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=AAA;MAPQ=41;MATEID=5128831_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_12_25333001_25358001_352C;SPAN=8522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:69 GQ:24.2 PL:[24.2, 0.0, 143.0] SR:10 DR:3 LR:-24.22 LO:29.08);ALT=C[chr12:25356854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	25362848	+	chr12	25378547	+	.	3	2	5128876_1	0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=5128876_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_25357501_25382501_257C;SPAN=15699;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:78 GQ:7.8 PL:[0.0, 7.8, 204.6] SR:2 DR:3 LR:7.928 LO:6.554);ALT=G[chr12:25378547[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	25398331	+	chr12	25403684	+	.	0	22	5128977_1	53.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5128977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_25382001_25407001_33C;SPAN=5353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:71 GQ:53.6 PL:[53.6, 0.0, 116.3] SR:22 DR:0 LR:-53.39 LO:54.76);ALT=T[chr12:25403684[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	25956130	-	chr12	125801147	+	.	36	0	5382534_1	99.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=5382534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:25956130(-)-12:125801147(-)__12_125783001_125808001D;SPAN=99845017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:0 DR:36 LR:-112.2 LO:112.2);ALT=[chr12:125801147[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	104359774	+	chr12	25956218	+	.	20	0	5318092_1	52.0	.	DISC_MAPQ=24;EVDNC=DSCRD;IMPRECISE;MAPQ=24;MATEID=5318092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:25956218(-)-12:104359774(+)__12_104345501_104370501D;SPAN=78403556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:49 GQ:52.7 PL:[52.7, 0.0, 65.9] SR:0 DR:20 LR:-52.75 LO:52.83);ALT=]chr12:104359774]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	27064252	+	chr12	27066390	+	.	6	2	5132772_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5132772_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_27048001_27073001_310C;SPAN=2138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:74 GQ:0 PL:[0.0, 0.0, 178.2] SR:2 DR:6 LR:0.2424 LO:11.06);ALT=T[chr12:27066390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27091643	+	chr12	27107078	+	.	0	31	5133060_1	89.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5133060_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_27097001_27122001_40C;SPAN=15435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:31 DR:0 LR:-89.12 LO:89.12);ALT=A[chr12:27107078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27127161	+	chr12	27128429	+	.	8	8	5133139_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5133139_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_27121501_27146501_305C;SPAN=1268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:89 GQ:25.4 PL:[25.4, 0.0, 190.4] SR:8 DR:8 LR:-25.4 LO:32.75);ALT=C[chr12:27128429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27156324	+	chr12	27167009	+	.	0	10	5133232_1	8.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=5133232_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_27146001_27171001_115C;SPAN=10685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:10 DR:0 LR:-8.898 LO:19.93);ALT=C[chr12:27167009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27175585	+	chr12	27181215	+	.	9	0	5133413_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5133413_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:27175585(+)-12:27181215(-)__12_27170501_27195501D;SPAN=5630;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=T[chr12:27181215[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27175596	+	chr12	27180277	+	.	15	0	5133414_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5133414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:27175596(+)-12:27180277(-)__12_27170501_27195501D;SPAN=4681;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:77 GQ:28.7 PL:[28.7, 0.0, 157.4] SR:0 DR:15 LR:-28.65 LO:33.8);ALT=T[chr12:27180277[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	27339449	-	chr12	27340467	+	.	8	0	5133687_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5133687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:27339449(-)-12:27340467(-)__12_27317501_27342501D;SPAN=1018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=[chr12:27340467[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	27863891	+	chr12	27869221	+	.	37	0	5135005_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5135005_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:27863891(+)-12:27869221(-)__12_27856501_27881501D;SPAN=5330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:84 GQ:99 PL:[99.5, 0.0, 102.8] SR:0 DR:37 LR:-99.38 LO:99.39);ALT=G[chr12:27869221[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	29302591	+	chr12	29324308	+	.	9	0	5138569_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5138569_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:29302591(+)-12:29324308(-)__12_29277501_29302501D;SPAN=21717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:9 DP:2 GQ:2.4 PL:[26.4, 2.4, 0.0] SR:0 DR:9 LR:-26.41 LO:26.41);ALT=C[chr12:29324308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	29523158	+	chr12	29524461	+	.	0	7	5139127_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5139127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_29522501_29547501_18C;SPAN=1303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:69 GQ:4.4 PL:[4.4, 0.0, 162.8] SR:7 DR:0 LR:-4.413 LO:13.62);ALT=G[chr12:29524461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	29844384	+	chr12	29846436	+	.	29	24	5139661_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAC;MAPQ=60;MATEID=5139661_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_29841001_29866001_27C;SPAN=2052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:52 GQ:10.5 PL:[145.2, 10.5, 0.0] SR:24 DR:29 LR:-145.2 LO:145.2);ALT=C[chr12:29846436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	30067279	-	chr12	31704716	+	.	8	0	5140366_1	17.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=5140366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:30067279(-)-12:31704716(-)__12_30061501_30086501D;SPAN=1637437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:0 DR:8 LR:-17.2 LO:18.78);ALT=[chr12:31704716[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	48095389	+	chr12	48096471	+	.	0	7	5177724_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5177724_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_48093501_48118501_189C;SPAN=1082;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:66 GQ:5.3 PL:[5.3, 0.0, 153.8] SR:7 DR:0 LR:-5.226 LO:13.76);ALT=T[chr12:48096471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	48096609	+	chr12	48099734	+	.	9	0	5177729_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5177729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:48096609(+)-12:48099734(-)__12_48093501_48118501D;SPAN=3125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:0 DR:9 LR:-6.951 LO:17.74);ALT=A[chr12:48099734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	48192783	+	chr12	48213608	+	.	12	0	5177928_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5177928_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:48192783(+)-12:48213608(-)__12_48191501_48216501D;SPAN=20825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:63 GQ:22.7 PL:[22.7, 0.0, 128.3] SR:0 DR:12 LR:-22.54 LO:26.91);ALT=A[chr12:48213608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	48358206	+	chr12	48359621	+	AGCAAGTAAATGAGTTGGTGGCTTTGATCCCACACAGTGATCAGAGATTGCGCCCTCAGCGAAC	0	25	5178123_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGCAAGTAAATGAGTTGGTGGCTTTGATCCCACACAGTGATCAGAGATTGCGCCCTCAGCGAAC;MAPQ=60;MATEID=5178123_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_48338501_48363501_328C;SPAN=1415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:96 GQ:56.6 PL:[56.6, 0.0, 175.4] SR:25 DR:0 LR:-56.52 LO:59.96);ALT=G[chr12:48359621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	48545089	+	chr12	48547150	+	.	0	10	5178785_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5178785_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_48534501_48559501_328C;SPAN=2061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:10 DR:0 LR:-9.711 LO:20.09);ALT=C[chr12:48547150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	48725481	+	chr12	48728381	+	.	24	12	5179573_1	89.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GTAATTAAGTTTATT;MAPQ=60;MATEID=5179573_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_48706001_48731001_97C;SPAN=2900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:49 GQ:29.6 PL:[89.0, 0.0, 29.6] SR:12 DR:24 LR:-90.68 LO:90.68);ALT=T[chr12:48728381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49108307	+	chr12	49110298	+	.	0	10	5180510_1	6.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5180510_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_49098001_49123001_36C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:99 GQ:6.2 PL:[6.2, 0.0, 233.9] SR:10 DR:0 LR:-6.189 LO:19.44);ALT=G[chr12:49110298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49239554	+	chr12	49245863	+	.	16	0	5180727_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5180727_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49239554(+)-12:49245863(-)__12_49245001_49270001D;SPAN=6309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.0 LO:39.93);ALT=C[chr12:49245863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49334973	+	chr12	49351092	+	.	44	21	5181180_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5181180_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_49318501_49343501_364C;SPAN=16119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:43 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:21 DR:44 LR:-161.7 LO:161.7);ALT=T[chr12:49351092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49399672	+	chr12	49412512	+	.	18	0	5181251_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5181251_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49399672(+)-12:49412512(-)__12_49392001_49417001D;SPAN=12840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:86 GQ:36.2 PL:[36.2, 0.0, 171.5] SR:0 DR:18 LR:-36.12 LO:41.2);ALT=A[chr12:49412512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49523522	+	chr12	49525104	+	.	133	0	5182092_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=5182092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49523522(+)-12:49525104(-)__12_49514501_49539501D;SPAN=1582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:133 DP:89 GQ:35.7 PL:[392.7, 35.7, 0.0] SR:0 DR:133 LR:-392.8 LO:392.8);ALT=A[chr12:49525104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49580617	+	chr12	49582760	+	.	111	23	5182017_1	99.0	.	DISC_MAPQ=17;EVDNC=ASDIS;HOMSEQ=C;MAPQ=0;MATEID=5182017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_49563501_49588501_187C;SPAN=2143;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:127 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:23 DR:111 LR:-376.3 LO:376.3);ALT=C[chr12:49582760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49658948	+	chr12	49663245	+	.	56	0	5182254_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5182254_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49658948(+)-12:49663245(-)__12_49661501_49686501D;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:65 GQ:10.8 PL:[178.2, 10.8, 0.0] SR:0 DR:56 LR:-180.4 LO:180.4);ALT=C[chr12:49663245[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49960049	+	chr12	49961830	+	.	14	0	5183133_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5183133_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49960049(+)-12:49961830(-)__12_49955501_49980501D;SPAN=1781;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:0 DR:14 LR:-27.52 LO:31.83);ALT=T[chr12:49961830[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	49960669	+	chr12	49961840	+	.	13	0	5183135_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5183135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:49960669(+)-12:49961840(-)__12_49955501_49980501D;SPAN=1171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:80 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:0 DR:13 LR:-21.24 LO:28.16);ALT=G[chr12:49961840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50135426	+	chr12	50146244	+	.	17	0	5183523_1	34.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5183523_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:50135426(+)-12:50146244(-)__12_50127001_50152001D;SPAN=10818;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:82 GQ:34.1 PL:[34.1, 0.0, 162.8] SR:0 DR:17 LR:-33.9 LO:38.83);ALT=G[chr12:50146244[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50135437	+	chr12	50146749	+	.	59	0	5183524_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5183524_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:50135437(+)-12:50146749(-)__12_50127001_50152001D;SPAN=11312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:89 GQ:45.2 PL:[170.6, 0.0, 45.2] SR:0 DR:59 LR:-174.7 LO:174.7);ALT=G[chr12:50146749[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50135437	+	chr12	50149414	+	.	23	0	5183525_1	50.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5183525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:50135437(+)-12:50149414(-)__12_50127001_50152001D;SPAN=13977;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:93 GQ:50.9 PL:[50.9, 0.0, 173.0] SR:0 DR:23 LR:-50.73 LO:54.56);ALT=G[chr12:50149414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50146332	+	chr12	50149415	+	AACCCCGTCAACGCAGCAGCACCTGAAGAAGGTCTATGCAAGTTTTGCCCTTTGTATGTTTGTGGCGGCTGCAGGGGCCTATGTCCATATGGTCACTCATTTCATT	5	118	5183553_1	99.0	.	DISC_MAPQ=48;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=AACCCCGTCAACGCAGCAGCACCTGAAGAAGGTCTATGCAAGTTTTGCCCTTTGTATGTTTGTGGCGGCTGCAGGGGCCTATGTCCATATGGTCACTCATTTCATT;MAPQ=60;MATEID=5183553_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_50127001_50152001_237C;SPAN=3083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:119 DP:100 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:118 DR:5 LR:-353.2 LO:353.2);ALT=T[chr12:50149415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50146865	+	chr12	50149415	+	.	3	58	5183555_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=5183555_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_12_50127001_50152001_237C;SPAN=2550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:112 GQ:98.6 PL:[171.2, 0.0, 98.6] SR:58 DR:3 LR:-172.0 LO:172.0);ALT=G[chr12:50149415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50153105	+	chr12	50155486	+	.	3	40	5184128_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5184128_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_50151501_50176501_208C;SPAN=2381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:120 GQ:99 PL:[106.1, 0.0, 185.3] SR:40 DR:3 LR:-106.1 LO:107.3);ALT=G[chr12:50155486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50155563	+	chr12	50156654	+	.	4	38	5184143_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5184143_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_50151501_50176501_330C;SPAN=1091;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:111 GQ:99 PL:[108.8, 0.0, 158.3] SR:38 DR:4 LR:-108.6 LO:109.1);ALT=G[chr12:50156654[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50506085	+	chr12	50513817	+	.	115	14	5184885_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5184885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_50494501_50519501_396C;SPAN=7732;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:122 DP:123 GQ:33 PL:[363.0, 33.0, 0.0] SR:14 DR:115 LR:-363.1 LO:363.1);ALT=G[chr12:50513817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	50794811	+	chr12	50821543	+	.	11	9	5185639_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5185639_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_50788501_50813501_58C;SPAN=26732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:39 GQ:38.9 PL:[55.4, 0.0, 38.9] SR:9 DR:11 LR:-55.6 LO:55.6);ALT=G[chr12:50821543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51442209	+	chr12	51450130	+	.	8	0	5188382_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5188382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:51442209(+)-12:51450130(-)__12_51425501_51450501D;SPAN=7921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=G[chr12:51450130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51442968	+	chr12	51450131	+	.	0	8	5188386_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5188386_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_51425501_51450501_198C;SPAN=7163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:77 GQ:5.6 PL:[5.6, 0.0, 180.5] SR:8 DR:0 LR:-5.547 LO:15.65);ALT=G[chr12:51450131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51632705	+	chr12	51634125	+	.	68	24	5188897_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5188897_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_51621501_51646501_341C;SPAN=1420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:103 GQ:24.3 PL:[297.0, 24.3, 0.0] SR:24 DR:68 LR:-296.7 LO:296.7);ALT=G[chr12:51634125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51632744	+	chr12	51634652	+	.	58	0	5188898_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5188898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:51632744(+)-12:51634652(-)__12_51621501_51646501D;SPAN=1908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:118 GQ:99 PL:[159.5, 0.0, 126.5] SR:0 DR:58 LR:-159.7 LO:159.7);ALT=T[chr12:51634652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51696573	+	chr12	51717802	+	.	8	0	5189312_1	0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5189312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:51696573(+)-12:51717802(-)__12_51695001_51720001D;SPAN=21229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:0 DR:8 LR:0.1426 LO:14.77);ALT=A[chr12:51717802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	51707689	+	chr12	51717804	+	.	17	13	5189353_1	54.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=0;MATEID=5189353_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=AGAG;SCTG=c_12_51695001_51720001_294C;SECONDARY;SPAN=10115;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:92 GQ:54.5 PL:[54.5, 0.0, 166.7] SR:13 DR:17 LR:-54.3 LO:57.58);ALT=T[chr12:51717804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53492089	+	chr12	53494494	+	.	9	0	5193857_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5193857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53492089(+)-12:53494494(-)__12_53483501_53508501D;SPAN=2405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:82 GQ:7.7 PL:[7.7, 0.0, 189.2] SR:0 DR:9 LR:-7.493 LO:17.84);ALT=A[chr12:53494494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53591736	+	chr12	53594027	+	.	0	8	5194252_1	3.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5194252_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53581501_53606501_31C;SPAN=2291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:8 DR:0 LR:-3.65 LO:15.33);ALT=C[chr12:53594027[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53594271	+	chr12	53600982	+	.	36	0	5194260_1	96.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5194260_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53594271(+)-12:53600982(-)__12_53581501_53606501D;SPAN=6711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:84 GQ:96.2 PL:[96.2, 0.0, 106.1] SR:0 DR:36 LR:-96.08 LO:96.12);ALT=A[chr12:53600982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53595012	+	chr12	53600985	+	.	10	0	5194265_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5194265_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53595012(+)-12:53600985(-)__12_53581501_53606501D;SPAN=5973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:0 DR:10 LR:-10.79 LO:20.31);ALT=C[chr12:53600985[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53689423	+	chr12	53691631	+	.	48	12	5194794_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=0;MATEID=5194794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53679501_53704501_127C;SECONDARY;SPAN=2208;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:174 GQ:99 PL:[141.2, 0.0, 279.8] SR:12 DR:48 LR:-141.0 LO:143.6);ALT=G[chr12:53691631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53690335	+	chr12	53691632	+	.	0	7	5194802_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5194802_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53679501_53704501_49C;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:154 GQ:18.4 PL:[0.0, 18.4, 409.3] SR:7 DR:0 LR:18.62 LO:11.1);ALT=G[chr12:53691632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53835823	+	chr19	40449669	-	.	43	0	6815630_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6815630_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53835823(+)-19:40449669(+)__19_40449501_40474501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:34 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:43 LR:-125.4 LO:125.4);ALT=C]chr19:40449669];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	53846160	+	chr12	53848508	+	.	36	71	5195674_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5195674_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_12_53826501_53851501_26C;SPAN=2348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:121 DP:197 GQ:99 PL:[346.1, 0.0, 131.6] SR:71 DR:36 LR:-351.3 LO:351.3);ALT=G[chr12:53848508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53846199	+	chr12	53849666	+	.	12	0	5195675_1	17.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=5195675_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53846199(+)-12:53849666(-)__12_53826501_53851501D;SPAN=3467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:0 DR:12 LR:-17.67 LO:25.46);ALT=T[chr12:53849666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53853162	+	chr12	53854796	+	.	8	0	5195392_1	2.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=5195392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:53853162(+)-12:53854796(-)__12_53851001_53876001D;SPAN=1634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=G[chr12:53854796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53854927	+	chr12	53856264	+	.	4	12	5195397_1	19.0	.	DISC_MAPQ=34;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5195397_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53851001_53876001_411C;SPAN=1337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:101 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:12 DR:4 LR:-18.85 LO:29.27);ALT=G[chr12:53856264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53856351	+	chr12	53862560	+	TTGACCAAGCTGCACCAGTTGGCAATGCAACAGTCTCATTTTCCCATGACGCATGGCAACACCGGATTCAGTGGCATTGAATCCAGCTCTCCAGAGGTGAAAGGCTATTGG	2	20	5195405_1	38.0	.	DISC_MAPQ=54;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTGACCAAGCTGCACCAGTTGGCAATGCAACAGTCTCATTTTCCCATGACGCATGGCAACACCGGATTCAGTGGCATTGAATCCAGCTCTCCAGAGGTGAAAGGCTATTGG;MAPQ=60;MATEID=5195405_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_53851001_53876001_127C;SPAN=6209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:104 GQ:38 PL:[38.0, 0.0, 212.9] SR:20 DR:2 LR:-37.84 LO:44.94);ALT=G[chr12:53862560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53937235	+	chr12	53946325	+	.	0	12	5195808_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5195808_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_53924501_53949501_111C;SPAN=9090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:12 DR:0 LR:-17.67 LO:25.46);ALT=G[chr12:53946325[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53946424	+	chr12	54020063	+	TCCACAGCCCGGGGCATTGCACACAAACGGTCTGTCGTCTCCCATATTTCATATAGCAGAGAGGAG	13	18	5195945_1	65.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCCACAGCCCGGGGCATTGCACACAAACGGTCTGTCGTCTCCCATATTTCATATAGCAGAGAGGAG;MAPQ=60;MATEID=5195945_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_53998001_54023001_421C;SPAN=73639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:39 GQ:29 PL:[65.3, 0.0, 29.0] SR:18 DR:13 LR:-66.1 LO:66.1);ALT=G[chr12:54020063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	53994806	+	chr12	54020063	+	.	10	8	5195946_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5195946_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_53998001_54023001_421C;SPAN=25257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:8 DR:10 LR:-25.75 LO:26.84);ALT=C[chr12:54020063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54063128	+	chr12	54066356	+	.	47	0	5196112_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5196112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54063128(+)-12:54066356(-)__12_54047001_54072001D;SPAN=3228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:102 GQ:99 PL:[127.7, 0.0, 117.8] SR:0 DR:47 LR:-127.5 LO:127.5);ALT=G[chr12:54066356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54063192	+	chr12	54069834	+	.	18	0	5196113_1	24.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5196113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54063192(+)-12:54069834(-)__12_54047001_54072001D;SPAN=6642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:128 GQ:24.8 PL:[24.8, 0.0, 285.5] SR:0 DR:18 LR:-24.74 LO:37.75);ALT=C[chr12:54069834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54063899	+	chr12	54066360	+	.	6	3	5196118_1	1.0	.	DISC_MAPQ=25;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5196118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_54047001_54072001_371C;SPAN=2461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:3 DR:6 LR:-1.533 LO:16.86);ALT=C[chr12:54066360[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54066457	+	chr12	54069836	+	.	8	0	5196126_1	0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5196126_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54066457(+)-12:54069836(-)__12_54047001_54072001D;SPAN=3379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:143 GQ:12 PL:[0.0, 12.0, 369.6] SR:0 DR:8 LR:12.33 LO:13.42);ALT=C[chr12:54069836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54119020	+	chr12	54121186	+	.	16	0	5196448_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5196448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54119020(+)-12:54121186(-)__12_54096001_54121001D;SPAN=2166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:0 DR:16 LR:-39.54 LO:40.27);ALT=C[chr12:54121186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54646011	+	chr12	54651297	+	.	0	10	5197785_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5197785_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_54635001_54660001_32C;SPAN=5286;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:10 DR:0 LR:-13.77 LO:20.98);ALT=C[chr12:54651297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54651499	+	chr12	54673799	+	.	20	0	5198161_1	54.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5198161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54651499(+)-12:54673799(-)__12_54659501_54684501D;SPAN=22300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:42 GQ:44.9 PL:[54.8, 0.0, 44.9] SR:0 DR:20 LR:-54.67 LO:54.67);ALT=G[chr12:54673799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54668164	+	chr12	54673818	+	.	8	0	5198184_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5198184_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54668164(+)-12:54673818(-)__12_54659501_54684501D;SPAN=5654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=G[chr12:54673818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54687170	+	chr12	54688918	+	.	0	9	5198066_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CCTGCA;MAPQ=60;MATEID=5198066_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_54684001_54709001_104C;SPAN=1748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:92 GQ:5 PL:[5.0, 0.0, 216.2] SR:9 DR:0 LR:-4.784 LO:17.36);ALT=A[chr12:54688918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54689093	+	chr12	54694583	+	.	25	29	5198076_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTGTG;MAPQ=60;MATEID=5198076_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_54684001_54709001_223C;SPAN=5490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:82 GQ:77 PL:[119.9, 0.0, 77.0] SR:29 DR:25 LR:-120.2 LO:120.2);ALT=G[chr12:54694583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54719014	+	chr12	54735987	+	.	30	0	5198485_1	95.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5198485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54719014(+)-12:54735987(-)__12_54708501_54733501D;SPAN=16973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:35 GQ:6 PL:[95.7, 6.0, 0.0] SR:0 DR:30 LR:-96.41 LO:96.41);ALT=G[chr12:54735987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54719017	+	chr12	54737008	+	.	32	0	5198486_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5198486_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54719017(+)-12:54737008(-)__12_54708501_54733501D;SPAN=17991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:35 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:0 DR:32 LR:-102.3 LO:102.3);ALT=G[chr12:54737008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54734399	+	chr12	54737009	+	TACTATGACGACACCTACCCCAGTGTCAAGGAGCAAAAGGCCTTTGAGAAGAACATTTTCAACAAGACCCATCGGACTGACA	2	61	5198247_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=TACTATGACGACACCTACCCCAGTGTCAAGGAGCAAAAGGCCTTTGAGAAGAACATTTTCAACAAGACCCATCGGACTGACA;MAPQ=60;MATEID=5198247_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_54733001_54758001_266C;SPAN=2610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:83 GQ:14 PL:[185.6, 0.0, 14.0] SR:61 DR:2 LR:-193.9 LO:193.9);ALT=G[chr12:54737009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54737100	+	chr12	54741549	+	CTGATGCTTATGGCTGTTCTGAACTGTCTCTTCGACTCATTGAGCCAGATGCTG	2	24	5198254_1	58.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTGATGCTTATGGCTGTTCTGAACTGTCTCTTCGACTCATTGAGCCAGATGCTG;MAPQ=60;MATEID=5198254_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_54733001_54758001_158C;SPAN=4449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:100 GQ:58.7 PL:[58.7, 0.0, 184.1] SR:24 DR:2 LR:-58.73 LO:62.34);ALT=G[chr12:54741549[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54849937	+	chr12	54854161	+	TTGATGAGATAGGTATTCAGTTACTGTGCATTTCCAT	0	23	5198658_1	55.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=TTGATGAGATAGGTATTCAGTTACTGTGCATTTCCAT;MAPQ=60;MATEID=5198658_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_54831001_54856001_252C;SPAN=4224;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:77 GQ:55.1 PL:[55.1, 0.0, 131.0] SR:23 DR:0 LR:-55.06 LO:56.8);ALT=T[chr12:54854161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54854258	+	chr12	54855893	+	.	0	7	5198666_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5198666_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_54831001_54856001_50C;SPAN=1635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:7 DR:0 LR:-0.8912 LO:13.07);ALT=G[chr12:54855893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54857083	+	chr12	54858851	+	.	0	18	5198686_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5198686_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_12_54855501_54880501_176C;SPAN=1768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:78 GQ:38.3 PL:[38.3, 0.0, 150.5] SR:18 DR:0 LR:-38.29 LO:42.07);ALT=T[chr12:54858851[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54857126	+	chr12	54867328	+	.	20	0	5198688_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5198688_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54857126(+)-12:54867328(-)__12_54855501_54880501D;SPAN=10202;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:92 GQ:41.3 PL:[41.3, 0.0, 179.9] SR:0 DR:20 LR:-41.1 LO:46.15);ALT=T[chr12:54867328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54858951	+	chr12	54865017	+	.	3	2	5198690_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5198690_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GG;SCTG=c_12_54855501_54880501_176C;SPAN=6066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:63 GQ:0.3 PL:[0.0, 0.3, 151.8] SR:2 DR:3 LR:0.5633 LO:9.169);ALT=G[chr12:54865017[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54858992	+	chr12	54867329	+	.	13	0	5198691_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5198691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:54858992(+)-12:54867329(-)__12_54855501_54880501D;SPAN=8337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:85 GQ:20 PL:[20.0, 0.0, 185.0] SR:0 DR:13 LR:-19.88 LO:27.78);ALT=G[chr12:54867329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54891675	+	chr12	54894316	+	ACTTGTTCAGACCCCAAATCTAAGCCACCTTTCTTACTGGAAAAGTCCATGGAACCATCTCTCAAGTATATCAACAAGAAATTTCCCAACATAGATGTCCGAAACAGCAC	11	21	5199091_1	63.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACTTGTTCAGACCCCAAATCTAAGCCACCTTTCTTACTGGAAAAGTCCATGGAACCATCTCTCAAGTATATCAACAAGAAATTTCCCAACATAGATGTCCGAAACAGCAC;MAPQ=60;MATEID=5199091_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_54880001_54905001_260C;SPAN=2641;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:94 GQ:63.8 PL:[63.8, 0.0, 162.8] SR:21 DR:11 LR:-63.66 LO:66.13);ALT=G[chr12:54894316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	54891675	+	chr12	54893137	+	.	19	9	5199090_1	31.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5199090_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_12_54880001_54905001_260C;SPAN=1462;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:86 GQ:31.5 PL:[31.5, 0.0, 122.5] SR:9 DR:19 LR:-31.34 LO:35.03);ALT=G[chr12:54893137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56110415	+	chr12	56112873	+	.	81	0	5201743_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5201743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56110415(+)-12:56112873(-)__12_56105001_56130001D;SPAN=2458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:125 GQ:68.6 PL:[233.6, 0.0, 68.6] SR:0 DR:81 LR:-238.4 LO:238.4);ALT=T[chr12:56112873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56110789	+	chr12	56112874	+	.	0	128	5201746_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5201746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56105001_56130001_84C;SPAN=2085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:128 DP:168 GQ:30.4 PL:[377.0, 0.0, 30.4] SR:128 DR:0 LR:-394.4 LO:394.4);ALT=G[chr12:56112874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56120801	+	chr12	56122735	+	.	16	0	5201780_1	22.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5201780_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56120801(+)-12:56122735(-)__12_56105001_56130001D;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:114 GQ:22.1 PL:[22.1, 0.0, 253.1] SR:0 DR:16 LR:-21.93 LO:33.54);ALT=C[chr12:56122735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56121170	+	chr12	56122734	+	.	117	0	5201784_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5201784_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56121170(+)-12:56122734(-)__12_56105001_56130001D;SPAN=1564;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:106 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:0 DR:117 LR:-346.6 LO:346.6);ALT=G[chr12:56122734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56194736	+	chr12	56211447	+	.	40	0	5202113_1	99.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=5202113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56194736(+)-12:56211447(-)__12_56203001_56228001D;SPAN=16711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:68 GQ:50.9 PL:[113.6, 0.0, 50.9] SR:0 DR:40 LR:-114.9 LO:114.9);ALT=T[chr12:56211447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56296139	+	chr12	56297171	+	.	0	7	5202400_1	1.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5202400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56276501_56301501_330C;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:7 DR:0 LR:-0.8912 LO:13.07);ALT=T[chr12:56297171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56297304	+	chr12	56321594	+	.	8	0	5202429_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5202429_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56297304(+)-12:56321594(-)__12_56301001_56326001D;SPAN=24290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=T[chr12:56321594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56308152	+	chr12	56321508	+	.	0	14	5202457_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5202457_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56301001_56326001_273C;SPAN=13356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:100 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:14 DR:0 LR:-19.12 LO:29.33);ALT=T[chr12:56321508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56308152	+	chr12	56309226	+	.	0	10	5202456_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5202456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56301001_56326001_90C;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:10 DR:0 LR:-8.898 LO:19.93);ALT=T[chr12:56309226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56367964	+	chr12	56380697	+	.	9	0	5202771_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5202771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56367964(+)-12:56380697(-)__12_56374501_56399501D;SPAN=12733;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:18 GQ:18.2 PL:[24.8, 0.0, 18.2] SR:0 DR:9 LR:-24.88 LO:24.88);ALT=C[chr12:56380697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56549377	+	chr12	56551251	+	.	0	29	5203568_1	64.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5203568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56546001_56571001_91C;SPAN=1874;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:117 GQ:64.1 PL:[64.1, 0.0, 219.2] SR:29 DR:0 LR:-64.03 LO:68.82);ALT=G[chr12:56551251[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56552242	+	chr12	56553365	+	.	89	0	5203588_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5203588_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56552242(+)-12:56553365(-)__12_56546001_56571001D;SPAN=1123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:89 DP:116 GQ:18.2 PL:[262.4, 0.0, 18.2] SR:0 DR:89 LR:-274.8 LO:274.8);ALT=G[chr12:56553365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56552242	+	chr12	56553757	+	.	53	0	5203589_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5203589_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56552242(+)-12:56553757(-)__12_56546001_56571001D;SPAN=1515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:135 GQ:99 PL:[138.5, 0.0, 188.0] SR:0 DR:53 LR:-138.4 LO:138.8);ALT=G[chr12:56553757[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56552550	+	chr12	56553777	+	.	8	0	5203590_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5203590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56552550(+)-12:56553777(-)__12_56546001_56571001D;SPAN=1227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:218 GQ:32.5 PL:[0.0, 32.5, 594.1] SR:0 DR:8 LR:32.65 LO:11.93);ALT=C[chr12:56553777[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56581092	+	chr12	56583135	+	.	17	7	5203389_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5203389_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56570501_56595501_110C;SPAN=2043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:78 GQ:41.6 PL:[41.6, 0.0, 147.2] SR:7 DR:17 LR:-41.59 LO:44.92);ALT=T[chr12:56583135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56610404	+	chr12	56615588	+	.	14	0	5203507_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5203507_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56610404(+)-12:56615588(-)__12_56595001_56620001D;SPAN=5184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:77 GQ:25.4 PL:[25.4, 0.0, 160.7] SR:0 DR:14 LR:-25.35 LO:31.08);ALT=A[chr12:56615588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	56694049	-	chr19	18141437	+	.	10	0	5203902_1	20.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5203902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:56694049(-)-19:18141437(-)__12_56693001_56718001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:47 GQ:20.3 PL:[20.3, 0.0, 92.9] SR:0 DR:10 LR:-20.28 LO:22.97);ALT=[chr19:18141437[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	56750365	+	chr12	56753842	+	.	8	2	5204112_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=5204112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_56742001_56767001_227C;SPAN=3477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:2 DR:8 LR:0.9554 LO:14.66);ALT=G[chr12:56753842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57032210	+	chr12	57036241	+	CCAAAATCTGCTGGAATCCTTTGATGGTCTCCTTCAGGGGTACCAGCTTCCCCATATGACCTGTGAAGACCTCAGCAACCTGGAATGGCTGAGACAAGAAACGCTGTATTTTCCGTGCACGGGACACGGTCAACTTGTCTTCCTCAGAAAGTTCATCCATACCCAGGATGGCAATGATATCCTGGAGGGATTTGTAGTCCTGCAGGATCTTTTGCACCCCACGGGCAACATCGTAATGCTCACTGCCAACAATGTTGGGATCCATGATACGAGAGGTGGAGTCTAGAGGATCCACAGCTGGATAGATGCCCAGCTCAGCAATGGCACGCGACAGTACAGTGGTAGCATCCAAATGGGCAAACGTAGTAGCAGGGGCAGGGTCAGTCAAGTCATCAGCAGGCACATAGATAG	0	104	5205018_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CCAAAATCTGCTGGAATCCTTTGATGGTCTCCTTCAGGGGTACCAGCTTCCCCATATGACCTGTGAAGACCTCAGCAACCTGGAATGGCTGAGACAAGAAACGCTGTATTTTCCGTGCACGGGACACGGTCAACTTGTCTTCCTCAGAAAGTTCATCCATACCCAGGATGGCAATGATATCCTGGAGGGATTTGTAGTCCTGCAGGATCTTTTGCACCCCACGGGCAACATCGTAATGCTCACTGCCAACAATGTTGGGATCCATGATACGAGAGGTGGAGTCTAGAGGATCCACAGCTGGATAGATGCCCAGCTCAGCAATGGCACGCGACAGTACAGTGGTAGCATCCAAATGGGCAAACGTAGTAGCAGGGGCAGGGTCAGTCAAGTCATCAGCAGGCACATAGATAG;MAPQ=60;MATEID=5205018_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_57011501_57036501_317C;SPAN=4031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:116 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:104 DR:0 LR:-342.1 LO:342.1);ALT=G[chr12:57036241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57033978	+	chr12	57036241	+	.	13	14	5205047_1	65.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=5205047_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_57036001_57061001_414C;SPAN=2263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:37 GQ:23 PL:[65.9, 0.0, 23.0] SR:14 DR:13 LR:-66.98 LO:66.98);ALT=T[chr12:57036241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57037409	+	chr12	57038564	+	.	9	0	5205056_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5205056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57037409(+)-12:57038564(-)__12_57036001_57061001D;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:66 GQ:11.9 PL:[11.9, 0.0, 147.2] SR:0 DR:9 LR:-11.83 LO:18.75);ALT=T[chr12:57038564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57066858	+	chr12	57081845	+	.	45	0	5205323_1	98.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5205323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57066858(+)-12:57081845(-)__12_57060501_57085501D;SPAN=14987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:184 GQ:98.9 PL:[98.9, 0.0, 346.4] SR:0 DR:45 LR:-98.7 LO:106.5);ALT=G[chr12:57081845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57493875	+	chr12	57496072	+	.	3	3	5206657_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5206657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_57477001_57502001_47C;SPAN=2197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:92 GQ:8.1 PL:[0.0, 8.1, 237.6] SR:3 DR:3 LR:8.42 LO:8.321);ALT=T[chr12:57496072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57640684	+	chr12	57642489	+	AGAGATCTTTGACACAAGCGTACTGCTGGTTGCTGTAGAGTGGGGAACTATAGGCCCGATGGAAACCAGGTGG	0	47	5207079_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=AGAGATCTTTGACACAAGCGTACTGCTGGTTGCTGTAGAGTGGGGAACTATAGGCCCGATGGAAACCAGGTGG;MAPQ=60;MATEID=5207079_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_57624001_57649001_366C;SPAN=1805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:109 GQ:99 PL:[125.6, 0.0, 138.8] SR:47 DR:0 LR:-125.6 LO:125.7);ALT=G[chr12:57642489[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57911588	+	chr12	57914200	+	.	42	0	5208090_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5208090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57911588(+)-12:57914200(-)__12_57893501_57918501D;SPAN=2612;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:66 GQ:38.3 PL:[120.8, 0.0, 38.3] SR:0 DR:42 LR:-123.0 LO:123.0);ALT=C[chr12:57914200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57929629	+	chr12	57939810	+	.	0	33	5207875_1	81.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5207875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_57918001_57943001_133C;SPAN=10181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:100 GQ:81.8 PL:[81.8, 0.0, 161.0] SR:33 DR:0 LR:-81.84 LO:83.25);ALT=C[chr12:57939810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	57929679	+	chr12	57940856	+	.	37	0	5207876_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5207876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:57929679(+)-12:57940856(-)__12_57918001_57943001D;SPAN=11177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:110 GQ:92.3 PL:[92.3, 0.0, 174.8] SR:0 DR:37 LR:-92.34 LO:93.73);ALT=A[chr12:57940856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	58109978	+	chr12	58111652	+	GCGAGCCCGACCAAGGATGACAGTAAGGACTCAGATTTCTGGAAGATGCTTAATGAGCCAGAGGACCAGGCCCCAGGAGGGGAGGAGGTGCCGGCTGAGGAGCAGGACCCAAGCCCTGAGGCAGCAGATTCAGCTTCTGGTGCTCCCAAT	2	19	5208570_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=GCGAGCCCGACCAAGGATGACAGTAAGGACTCAGATTTCTGGAAGATGCTTAATGAGCCAGAGGACCAGGCCCCAGGAGGGGAGGAGGTGCCGGCTGAGGAGCAGGACCCAAGCCCTGAGGCAGCAGATTCAGCTTCTGGTGCTCCCAAT;MAPQ=60;MATEID=5208570_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_58089501_58114501_91C;SPAN=1674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:68 GQ:44.3 PL:[44.3, 0.0, 120.2] SR:19 DR:2 LR:-44.3 LO:46.26);ALT=T[chr12:58111652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	58325567	+	chr12	58329644	+	.	12	0	5209551_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5209551_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:58325567(+)-12:58329644(-)__12_58310001_58335001D;SPAN=4077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:209 GQ:16.9 PL:[0.0, 16.9, 541.3] SR:0 DR:12 LR:17.01 LO:20.26);ALT=T[chr12:58329644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	76361973	+	chr12	58469677	+	.	9	0	7454139_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7454139_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:58469677(-)-23:76361973(+)__23_76342001_76367001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:36 GQ:20 PL:[20.0, 0.0, 66.2] SR:0 DR:9 LR:-19.96 LO:21.4);ALT=]chrX:76361973]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	62649095	+	chr12	62652544	+	.	0	12	5218878_1	20.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5218878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_62646501_62671501_175C;SPAN=3449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:73 GQ:20 PL:[20.0, 0.0, 155.3] SR:12 DR:0 LR:-19.83 LO:26.06);ALT=T[chr12:62652544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	62654271	+	chr12	62696568	+	.	20	0	5218990_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5218990_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:62654271(+)-12:62696568(-)__12_62695501_62720501D;SPAN=42297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:46 GQ:53.6 PL:[53.6, 0.0, 56.9] SR:0 DR:20 LR:-53.56 LO:53.57);ALT=A[chr12:62696568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	62654287	+	chr12	62687959	+	.	48	14	5218937_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTA;MAPQ=60;MATEID=5218937_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_62671001_62696001_165C;SPAN=33672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:33 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:14 DR:48 LR:-151.8 LO:151.8);ALT=A[chr12:62687959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	62696703	+	chr12	62708569	+	.	0	9	5218994_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5218994_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_62695501_62720501_233C;SPAN=11866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:9 DR:0 LR:-10.2 LO:18.38);ALT=T[chr12:62708569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	65672646	+	chr12	65720605	+	.	10	10	5227075_1	46.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5227075_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_65709001_65734001_163C;SPAN=47959;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:35 GQ:36.8 PL:[46.7, 0.0, 36.8] SR:10 DR:10 LR:-46.68 LO:46.68);ALT=G[chr12:65720605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	65720714	+	chr12	65722304	+	.	0	12	5227110_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5227110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_65709001_65734001_223C;SPAN=1590;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:71 GQ:20.6 PL:[20.6, 0.0, 149.3] SR:12 DR:0 LR:-20.38 LO:26.22);ALT=G[chr12:65722304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	65847605	+	chr12	65856931	+	.	3	7	5227364_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=5227364_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_65856001_65881001_173C;SPAN=9326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:7 DR:3 LR:-18.6 LO:20.81);ALT=G[chr12:65856931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66522894	+	chr12	66524482	+	.	13	0	5229081_1	17.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=5229081_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:66522894(+)-12:66524482(-)__12_66517501_66542501D;SPAN=1588;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:95 GQ:17.3 PL:[17.3, 0.0, 212.0] SR:0 DR:13 LR:-17.18 LO:27.1);ALT=C[chr12:66524482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66527651	+	chr12	66529877	+	.	70	36	5229088_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GAAAATGGTATTAATA;MAPQ=60;MATEID=5229088_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_66517501_66542501_131C;SPAN=2226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:30 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:36 DR:70 LR:-257.5 LO:257.5);ALT=A[chr12:66529877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66531948	+	chr12	66539620	+	TCAAGAATCCTGACAGGCACAATATCCACAAAAGAGCAAACAG	7	19	5229097_1	61.0	.	DISC_MAPQ=53;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TCAAGAATCCTGACAGGCACAATATCCACAAAAGAGCAAACAG;MAPQ=60;MATEID=5229097_2;MATENM=0;NM=2;NUMPARTS=3;SCTG=c_12_66517501_66542501_324C;SPAN=7672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:66 GQ:61.4 PL:[61.4, 0.0, 97.7] SR:19 DR:7 LR:-61.34 LO:61.82);ALT=T[chr12:66539620[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66539739	+	chr12	66547120	+	AACAACTGCCACAGTCAGAGCTTCCAACAGCGTAAATCCAAAAAGTAGGTACAGGTTAAGGGGATACTTATGTCTGTTTAAAATCAACGCAAAAATCAAACCCAGAGATCCGAGGGCAAACAGCAAAATTAAGGCAGGA	0	65	5228989_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AACAACTGCCACAGTCAGAGCTTCCAACAGCGTAAATCCAAAAAGTAGGTACAGGTTAAGGGGATACTTATGTCTGTTTAAAATCAACGCAAAAATCAAACCCAGAGATCCGAGGGCAAACAGCAAAATTAAGGCAGGA;MAPQ=60;MATEID=5228989_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_66542001_66567001_65C;SPAN=7381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:46 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:65 DR:0 LR:-191.4 LO:191.4);ALT=C[chr12:66547120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66539739	+	chr12	66546051	+	AACAACTGCCACAGTCAGAGCTTCCAACAGCGT	3	23	5229106_1	85.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=AACAACTGCCACAGTCAGAGCTTCCAACAGCGT;MAPQ=60;MATEID=5229106_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_66517501_66542501_190C;SPAN=6312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:29 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:23 DR:3 LR:-85.54 LO:85.54);ALT=C[chr12:66546051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66546210	+	chr12	66563674	+	.	42	0	5229007_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5229007_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:66546210(+)-12:66563674(-)__12_66542001_66567001D;SPAN=17464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:85 GQ:89.3 PL:[115.7, 0.0, 89.3] SR:0 DR:42 LR:-115.8 LO:115.8);ALT=T[chr12:66563674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66547229	+	chr12	66563635	+	.	50	16	5229008_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5229008_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_66542001_66567001_87C;SPAN=16406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:75 GQ:19.4 PL:[161.3, 0.0, 19.4] SR:16 DR:50 LR:-167.5 LO:167.5);ALT=C[chr12:66563635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	66554940	+	chr12	66563677	+	.	13	0	5229023_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5229023_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:66554940(+)-12:66563677(-)__12_66542001_66567001D;SPAN=8737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:0 DR:13 LR:-15.01 LO:26.61);ALT=T[chr12:66563677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69080854	+	chr12	69082740	+	.	4	3	5234917_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5234917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69065501_69090501_278C;SPAN=1886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:3 DR:4 LR:-2.788 LO:13.35);ALT=G[chr12:69082740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69080877	+	chr12	69083310	+	.	9	0	5234918_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5234918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69080877(+)-12:69083310(-)__12_69065501_69090501D;SPAN=2433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:0 DR:9 LR:-6.951 LO:17.74);ALT=A[chr12:69083310[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69633487	+	chr12	69644906	+	.	34	6	5236722_1	98.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5236722_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69629001_69654001_357C;SPAN=11419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:87 GQ:98.6 PL:[98.6, 0.0, 111.8] SR:6 DR:34 LR:-98.57 LO:98.62);ALT=G[chr12:69644906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69649618	+	chr17	4287349	+	.	11	0	5236758_1	23.0	.	DISC_MAPQ=11;EVDNC=DSCRD;IMPRECISE;MAPQ=11;MATEID=5236758_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69649618(+)-17:4287349(-)__12_69629001_69654001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:47 GQ:23.6 PL:[23.6, 0.0, 89.6] SR:0 DR:11 LR:-23.58 LO:25.79);ALT=C[chr17:4287349[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	69653977	+	chr12	69656150	+	.	4	6	5236775_1	4.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAG;MAPQ=60;MATEID=5236775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69653501_69678501_219C;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:81 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:6 DR:4 LR:-4.463 LO:15.47);ALT=G[chr12:69656150[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69742325	+	chr12	69743888	+	.	121	189	5237477_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5237477_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_69727001_69752001_255C;SPAN=1563;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:271 DP:364 GQ:86.4 PL:[796.1, 0.0, 86.4] SR:189 DR:121 LR:-829.0 LO:829.0);ALT=G[chr12:69743888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69742376	+	chr12	69745998	+	.	11	0	5237480_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5237480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69742376(+)-12:69745998(-)__12_69727001_69752001D;SPAN=3622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:134 GQ:0.2 PL:[0.2, 0.0, 323.6] SR:0 DR:11 LR:-0.007112 LO:20.34);ALT=C[chr12:69745998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69744052	+	chr12	69745999	+	.	6	64	5237484_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5237484_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_12_69727001_69752001_255C;SPAN=1947;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:199 GQ:99 PL:[177.2, 0.0, 305.9] SR:64 DR:6 LR:-177.2 LO:179.0);ALT=G[chr12:69745999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69744102	+	chr12	69746931	+	.	14	0	5237485_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5237485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69744102(+)-12:69746931(-)__12_69727001_69752001D;SPAN=2829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:110 GQ:16.4 PL:[16.4, 0.0, 250.7] SR:0 DR:14 LR:-16.41 LO:28.71);ALT=G[chr12:69746931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69979351	+	chr12	69980529	+	.	38	0	5237729_1	98.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5237729_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69979351(+)-12:69980529(-)__12_69972001_69997001D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:98 GQ:98.9 PL:[98.9, 0.0, 138.5] SR:0 DR:38 LR:-98.89 LO:99.26);ALT=C[chr12:69980529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69982042	+	chr12	69983264	+	.	7	4	5237739_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5237739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69972001_69997001_338C;SPAN=1222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:4 DR:7 LR:-7.543 LO:19.68);ALT=G[chr12:69983264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69983468	+	chr12	69985837	+	.	0	19	5237745_1	40.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5237745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69972001_69997001_42C;SPAN=2369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:84 GQ:40.1 PL:[40.1, 0.0, 162.2] SR:19 DR:0 LR:-39.96 LO:44.22);ALT=G[chr12:69985837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69986911	+	chr12	69990933	+	.	8	0	5237758_1	5.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5237758_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:69986911(+)-12:69990933(-)__12_69972001_69997001D;SPAN=4022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:0 DR:8 LR:-5.276 LO:15.61);ALT=T[chr12:69990933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	69993785	+	chr12	69995073	+	.	6	26	5237787_1	70.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5237787_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_69972001_69997001_209C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:94 GQ:70.4 PL:[70.4, 0.0, 156.2] SR:26 DR:6 LR:-70.26 LO:72.12);ALT=G[chr12:69995073[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70594864	+	chr12	70597578	+	.	63	36	5239429_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAAAGTATGACACTTC;MAPQ=60;MATEID=5239429_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_70584501_70609501_34C;SPAN=2714;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:56 GQ:21 PL:[231.0, 21.0, 0.0] SR:36 DR:63 LR:-231.1 LO:231.1);ALT=C[chr12:70597578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70637308	+	chr12	70704672	+	.	11	0	5239514_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5239514_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:70637308(+)-12:70704672(-)__12_70682501_70707501D;SPAN=67364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:0 DR:11 LR:-26.29 LO:27.14);ALT=G[chr12:70704672[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70672056	+	chr12	70704673	+	.	3	14	5239515_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5239515_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_70682501_70707501_222C;SPAN=32617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:37 GQ:39.5 PL:[39.5, 0.0, 49.4] SR:14 DR:3 LR:-39.49 LO:39.56);ALT=T[chr12:70704673[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70738008	+	chr12	70739960	+	.	0	9	5239478_1	9.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5239478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_70731501_70756501_261C;SPAN=1952;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:9 DR:0 LR:-9.661 LO:18.26);ALT=T[chr12:70739960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	70872266	+	chr12	70878218	+	C	0	77	5239796_1	99.0	.	EVDNC=ASSMB;INSERTION=C;MAPQ=60;MATEID=5239796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_70854001_70879001_97C;SPAN=5952;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:38 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:77 DR:0 LR:-227.8 LO:227.8);ALT=G[chr12:70878218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	71602361	+	chr12	71604474	+	.	40	26	5241454_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TACT;MAPQ=60;MATEID=5241454_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_71589001_71614001_136C;SPAN=2113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:43 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:26 DR:40 LR:-151.8 LO:151.8);ALT=T[chr12:71604474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	73239572	-	chr15	94886290	+	ATATATATATATTTTC	20	33	6044573_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;INSERTION=ATATATATATATTTTC;MAPQ=30;MATEID=6044573_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_94864001_94889001_15C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:39 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:33 DR:20 LR:-125.4 LO:125.4);ALT=[chr15:94886290[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr12	73239578	+	chr15	94888547	-	.	71	39	6044574_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=6044574_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_94864001_94889001_17C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:99 DP:40 GQ:26.7 PL:[293.7, 26.7, 0.0] SR:39 DR:71 LR:-293.8 LO:293.8);ALT=G]chr15:94888547];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	75875861	+	chr12	75884182	+	.	15	6	5251112_1	48.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=TCAGGT;MAPQ=60;MATEID=5251112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75876501_75901501_323C;SPAN=8321;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:41 GQ:48.5 PL:[48.5, 0.0, 48.5] SR:6 DR:15 LR:-48.31 LO:48.32);ALT=T[chr12:75884182[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75875901	+	chr12	75889353	+	.	10	0	5250888_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5250888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:75875901(+)-12:75889353(-)__12_75852001_75877001D;SPAN=13452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:40 GQ:22.1 PL:[22.1, 0.0, 74.9] SR:0 DR:10 LR:-22.17 LO:23.78);ALT=G[chr12:75889353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75884298	+	chr12	75889356	+	.	0	45	5251127_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5251127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75876501_75901501_294C;SPAN=5058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:97 GQ:99 PL:[122.3, 0.0, 112.4] SR:45 DR:0 LR:-122.3 LO:122.3);ALT=G[chr12:75889356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75884335	+	chr12	75892603	+	.	8	0	5251128_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5251128_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:75884335(+)-12:75892603(-)__12_75876501_75901501D;SPAN=8268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:0 DR:8 LR:0.6845 LO:14.7);ALT=C[chr12:75892603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75889442	+	chr12	75892604	+	TTAACCGACAGCGAGACCAAGTCAAAC	12	139	5251146_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTAACCGACAGCGAGACCAAGTCAAAC;MAPQ=60;MATEID=5251146_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75876501_75901501_113C;SPAN=3162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:155 GQ:41.8 PL:[458.8, 41.8, 0.0] SR:139 DR:12 LR:-458.8 LO:458.8);ALT=G[chr12:75892604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75900696	+	chr12	75902054	+	.	0	12	5251184_1	27.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5251184_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75876501_75901501_225C;SPAN=1358;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:46 GQ:27.2 PL:[27.2, 0.0, 83.3] SR:12 DR:0 LR:-27.15 LO:28.79);ALT=G[chr12:75902054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	75902228	+	chr12	75905293	+	.	19	4	5250953_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5250953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_75901001_75926001_41C;SPAN=3065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:67 GQ:51.2 PL:[51.2, 0.0, 110.6] SR:4 DR:19 LR:-51.17 LO:52.4);ALT=T[chr12:75905293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	76444480	+	chr12	76446988	+	.	13	0	5252542_1	19.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5252542_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76444480(+)-12:76446988(-)__12_76440001_76465001D;SPAN=2508;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:86 GQ:19.7 PL:[19.7, 0.0, 188.0] SR:0 DR:13 LR:-19.61 LO:27.71);ALT=T[chr12:76446988[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	76447691	+	chr12	76449814	+	.	8	0	5252555_1	2.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=5252555_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76447691(+)-12:76449814(-)__12_76440001_76465001D;SPAN=2123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=T[chr12:76449814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	76454070	+	chr12	76478346	+	.	8	0	5252585_1	18.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=5252585_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76454070(+)-12:76478346(-)__12_76440001_76465001D;SPAN=24276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=A[chr12:76478346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	76461291	+	chr12	76478346	+	.	28	0	5252614_1	82.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5252614_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76461291(+)-12:76478346(-)__12_76440001_76465001D;SPAN=17055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:36 GQ:3.5 PL:[82.7, 0.0, 3.5] SR:0 DR:28 LR:-86.83 LO:86.83);ALT=G[chr12:76478346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	76462802	+	chr12	76478346	+	.	42	0	5252619_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=5252619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:76462802(+)-12:76478346(-)__12_76440001_76465001D;SPAN=15544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:30 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=T[chr12:76478346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	81937176	+	chr19	18553332	+	.	8	0	6756560_1	5.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6756560_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:81937176(+)-19:18553332(-)__19_18546501_18571501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:0 DR:8 LR:-5.818 LO:15.7);ALT=A[chr19:18553332[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr12	82139719	+	chr12	82144320	+	.	31	17	5265170_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AACA;MAPQ=60;MATEID=5265170_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_12_82124001_82149001_249C;SPAN=4601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:69 GQ:50.6 PL:[116.6, 0.0, 50.6] SR:17 DR:31 LR:-118.1 LO:118.1);ALT=A[chr12:82144320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	82751073	+	chr12	82752468	+	.	23	0	5266591_1	58.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5266591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:82751073(+)-12:82752468(-)__12_82736501_82761501D;SPAN=1395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:66 GQ:58.1 PL:[58.1, 0.0, 101.0] SR:0 DR:23 LR:-58.04 LO:58.71);ALT=A[chr12:82752468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	87205881	+	chr12	87204874	+	.	19	0	5275969_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5275969_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:87204874(-)-12:87205881(+)__12_87195501_87220501D;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:52 GQ:48.8 PL:[48.8, 0.0, 75.2] SR:0 DR:19 LR:-48.63 LO:48.99);ALT=]chr12:87205881]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	88440755	+	chr12	88442009	+	.	0	5	5278771_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5278771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_88420501_88445501_279C;SPAN=1254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:83 GQ:5.7 PL:[0.0, 5.7, 211.2] SR:5 DR:0 LR:5.982 LO:8.55);ALT=T[chr12:88442009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	89172969	+	chr12	89184607	+	G	53	33	5280301_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=G;MAPQ=60;MATEID=5280301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_89180001_89205001_73C;SPAN=11638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:21 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:33 DR:53 LR:-214.6 LO:214.6);ALT=A[chr12:89184607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90024424	+	chr12	90028552	+	.	2	12	5282262_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCT;MAPQ=60;MATEID=5282262_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_90013001_90038001_109C;SPAN=4128;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:12 DR:2 LR:-27.52 LO:31.83);ALT=T[chr12:90028552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90036134	+	chr12	90049454	+	.	6	4	5282291_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5282291_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_90013001_90038001_163C;SPAN=13320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:32 GQ:17.9 PL:[17.9, 0.0, 57.5] SR:4 DR:6 LR:-17.74 LO:19.02);ALT=T[chr12:90049454[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90040799	+	chr12	90049456	+	.	0	10	5282126_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5282126_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_90037501_90062501_141C;SPAN=8657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:10 DR:0 LR:-7.272 LO:19.63);ALT=T[chr12:90049456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90049885	+	chr12	90102996	+	.	24	5	5282342_1	72.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5282342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_90086501_90111501_155C;SPAN=53111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:25 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:5 DR:24 LR:-72.62 LO:72.62);ALT=C[chr12:90102996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90049886	+	chr12	90102373	+	.	0	13	5282343_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5282343_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_12_90086501_90111501_184C;SPAN=52487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:20 GQ:11 PL:[37.4, 0.0, 11.0] SR:13 DR:0 LR:-38.29 LO:38.29);ALT=T[chr12:90102373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	90487005	+	chr12	90491695	+	ATATTAATATTAATATATATTATATATTTAATATATATATATATTAAATATATATAATTATATATATATTTAATATACATAAATAT	4	14	5283140_1	49.0	.	DISC_MAPQ=15;EVDNC=TSI_G;HOMSEQ=A;INSERTION=ATATTAATATTAATATATATTATATATTTAATATATATATATATTAAATATATATAATTATATATATATTTAATATACATAAATAT;MAPQ=60;MATEID=5283140_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_12_90478501_90503501_43C;SPAN=4690;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:19 GQ:1.8 PL:[49.5, 1.8, 0.0] SR:14 DR:4 LR:-51.04 LO:51.04);ALT=T[chr12:90491695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104324360	+	chr12	104326052	+	.	9	0	5318210_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5318210_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104324360(+)-12:104326052(-)__12_104321001_104346001D;SPAN=1692;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:0 DR:9 LR:-1.533 LO:16.86);ALT=A[chr12:104326052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104332279	+	chr12	104335184	+	.	11	0	5318235_1	15.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5318235_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104332279(+)-12:104335184(-)__12_104321001_104346001D;SPAN=2905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:0 DR:11 LR:-15.72 LO:23.22);ALT=T[chr12:104335184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104359630	-	chr12	125801148	+	.	18	40	5382537_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;MAPQ=60;MATEID=5382537_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_12_125783001_125808001_400C;SPAN=21441518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:39 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:40 DR:18 LR:-148.5 LO:148.5);ALT=[chr12:125801148[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	104378705	+	chr12	104380725	+	.	9	0	5318322_1	11.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=5318322_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104378705(+)-12:104380725(-)__12_104370001_104395001D;SPAN=2020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=T[chr12:104380725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104379506	+	chr12	104380726	+	.	14	15	5318328_1	68.0	.	DISC_MAPQ=47;EVDNC=ASDIS;MAPQ=60;MATEID=5318328_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_104370001_104395001_240C;SPAN=1220;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:75 GQ:68.9 PL:[68.9, 0.0, 111.8] SR:15 DR:14 LR:-68.81 LO:69.4);ALT=A[chr12:104380726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104680899	+	chr12	104705065	+	.	9	0	5319261_1	18.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5319261_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:104680899(+)-12:104705065(-)__12_104664001_104689001D;SPAN=24166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=G[chr12:104705065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	104707097	+	chr12	104709554	+	.	0	7	5319181_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=5319181_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_104688501_104713501_247C;SPAN=2457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:7 DR:0 LR:-0.6203 LO:13.03);ALT=T[chr12:104709554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105380247	+	chr12	105381943	+	.	11	10	5321050_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5321050_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_105374501_105399501_163C;SPAN=1696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:86 GQ:26.3 PL:[26.3, 0.0, 181.4] SR:10 DR:11 LR:-26.22 LO:33.0);ALT=T[chr12:105381943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105382031	+	chr12	105385490	+	.	0	11	5321052_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5321052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_105374501_105399501_264C;SPAN=3459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:91 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:11 DR:0 LR:-11.66 LO:22.29);ALT=T[chr12:105385490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105385627	+	chr12	105388255	+	.	3	13	5321059_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5321059_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_105374501_105399501_242C;SPAN=2628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:79 GQ:31.4 PL:[31.4, 0.0, 160.1] SR:13 DR:3 LR:-31.41 LO:36.36);ALT=G[chr12:105388255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105501638	+	chr12	105504902	+	.	13	0	5321333_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5321333_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:105501638(+)-12:105504902(-)__12_105497001_105522001D;SPAN=3264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:0 DR:13 LR:-20.7 LO:28.0);ALT=G[chr12:105504902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105556625	+	chr12	105557888	+	.	3	3	5321551_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5321551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_105546001_105571001_215C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:103 GQ:7.8 PL:[0.0, 7.8, 264.0] SR:3 DR:3 LR:8.099 LO:10.17);ALT=T[chr12:105557888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105724716	+	chr12	105761250	+	CCCTGCAGGAGCAGCCAAAGATGTAACAGAAGAATCCGTAACAGAAGATGACAAGAGGAGAAACTATGGAGGAGTATATGTTGGCCTACCATCTGAAGCTGTCAATATGGTGTCCAGTCAAACAAAGACGGTTCGGAAAA	2	22	5322183_1	79.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCCTGCAGGAGCAGCCAAAGATGTAACAGAAGAATCCGTAACAGAAGATGACAAGAGGAGAAACTATGGAGGAGTATATGTTGGCCTACCATCTGAAGCTGTCAATATGGTGTCCAGTCAAACAAAGACGGTTCGGAAAA;MAPQ=60;MATEID=5322183_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_12_105717501_105742501_371C;SPAN=36534;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:27 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:22 DR:2 LR:-78.52 LO:78.52);ALT=G[chr12:105761250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105724716	+	chr12	105759585	+	CCCTGCAGGAGCAGCCAAAGATGT	2	19	5322182_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_L;INSERTION=CCCTGCAGGAGCAGCCAAAGATGT;MAPQ=60;MATEID=5322182_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_12_105717501_105742501_371C;SPAN=34869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:27 GQ:2.6 PL:[62.0, 0.0, 2.6] SR:19 DR:2 LR:-65.13 LO:65.13);ALT=G[chr12:105759585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105724716	+	chr12	105742378	+	.	2	10	5322181_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5322181_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_105717501_105742501_235C;SPAN=17662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:10 DR:2 LR:-20.87 LO:24.74);ALT=G[chr12:105742378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105724727	+	chr12	105764409	+	.	10	0	5322184_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5322184_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:105724727(+)-12:105764409(-)__12_105717501_105742501D;SPAN=39682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:0 DR:10 LR:-26.78 LO:26.78);ALT=G[chr12:105764409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105724767	+	chr12	105760392	+	.	14	0	5322075_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5322075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:105724767(+)-12:105760392(-)__12_105742001_105767001D;SPAN=35625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:38 GQ:35.9 PL:[35.9, 0.0, 55.7] SR:0 DR:14 LR:-35.92 LO:36.17);ALT=G[chr12:105760392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	105761287	+	chr12	105764410	+	CCCTGCAGGAGCAGCCAAAGATGT	2	8	5322124_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;INSERTION=CCCTGCAGGAGCAGCCAAAGATGT;MAPQ=60;MATEID=5322124_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GAGA;SCTG=c_12_105742001_105767001_2C;SPAN=3123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:71 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:8 DR:2 LR:-10.47 LO:18.44);ALT=G[chr12:105764410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112204852	+	chr12	112220959	+	.	14	0	5340513_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5340513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112204852(+)-12:112220959(-)__12_112210001_112235001D;SPAN=16107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:46 GQ:33.8 PL:[33.8, 0.0, 76.7] SR:0 DR:14 LR:-33.75 LO:34.71);ALT=C[chr12:112220959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112204900	+	chr12	112219720	+	.	26	12	5340514_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5340514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_112210001_112235001_3C;SPAN=14820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:40 GQ:12.2 PL:[84.8, 0.0, 12.2] SR:12 DR:26 LR:-88.02 LO:88.02);ALT=G[chr12:112219720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112219827	+	chr12	112220960	+	.	0	24	5340542_1	56.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5340542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_112210001_112235001_187C;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:86 GQ:56 PL:[56.0, 0.0, 151.7] SR:24 DR:0 LR:-55.92 LO:58.42);ALT=G[chr12:112220960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112278283	+	chr12	112279488	+	.	6	7	5340793_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5340793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_112259001_112284001_350C;SPAN=1205;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:7 DR:6 LR:-6.951 LO:17.74);ALT=T[chr12:112279488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112451340	+	chr12	112457557	+	.	44	0	5341325_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5341325_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112451340(+)-12:112457557(-)__12_112430501_112455501D;SPAN=6217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:54 GQ:1.2 PL:[132.0, 1.2, 0.0] SR:0 DR:44 LR:-138.6 LO:138.6);ALT=T[chr12:112457557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	112451340	+	chr20	50727569	-	.	64	0	5341326_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5341326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112451340(+)-20:50727569(+)__12_112430501_112455501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:64 DP:54 GQ:17.1 PL:[188.1, 17.1, 0.0] SR:0 DR:64 LR:-188.1 LO:188.1);ALT=T]chr20:50727569];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	112563447	+	chr12	112572540	+	.	9	0	5341644_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5341644_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:112563447(+)-12:112572540(-)__12_112553001_112578001D;SPAN=9093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:0 DR:9 LR:-5.868 LO:17.54);ALT=C[chr12:112572540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	113019463	+	chr12	113020507	+	.	36	0	5343078_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5343078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:113019463(+)-12:113020507(-)__12_113018501_113043501D;SPAN=1044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:54 GQ:25.1 PL:[104.3, 0.0, 25.1] SR:0 DR:36 LR:-106.8 LO:106.8);ALT=C[chr12:113020507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	113618865	+	chr12	113623083	+	.	0	19	5344768_1	41.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5344768_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_113606501_113631501_10C;SPAN=4218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:77 GQ:41.9 PL:[41.9, 0.0, 144.2] SR:19 DR:0 LR:-41.86 LO:45.05);ALT=T[chr12:113623083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	113860306	+	chr12	113865803	+	.	16	0	5345539_1	26.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5345539_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:113860306(+)-12:113865803(-)__12_113851501_113876501D;SPAN=5497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:99 GQ:26 PL:[26.0, 0.0, 214.1] SR:0 DR:16 LR:-25.99 LO:34.61);ALT=G[chr12:113865803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	114400263	+	chr12	114404069	+	.	12	0	5347153_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5347153_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:114400263(+)-12:114404069(-)__12_114390501_114415501D;SPAN=3806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:0 DR:12 LR:-19.29 LO:25.9);ALT=C[chr12:114404069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	87426048	+	chr12	117013730	+	.	94	0	5353875_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=5353875_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:117013730(-)-16:87426048(+)__12_117012001_117037001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:57 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:0 DR:94 LR:-277.3 LO:277.3);ALT=]chr16:87426048]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	117086884	+	chr12	117088194	+	.	53	28	5354127_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGTGGCTCAGGCCTATAATCCCAGCACTT;MAPQ=60;MATEID=5354127_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_12_117085501_117110501_183C;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:35 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:28 DR:53 LR:-217.9 LO:217.9);ALT=T[chr12:117088194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	117477017	+	chr12	117484363	+	TCAGGAAGTCCTCGAAGGTGATCCCCTCGTACACCTGATCAGGCT	2	23	5355321_1	68.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TCAGGAAGTCCTCGAAGGTGATCCCCTCGTACACCTGATCAGGCT;MAPQ=60;MATEID=5355321_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_117477501_117502501_173C;SPAN=7346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:42 GQ:31.7 PL:[68.0, 0.0, 31.7] SR:23 DR:2 LR:-68.45 LO:68.45);ALT=T[chr12:117484363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	117486965	+	chr12	117494610	+	.	0	10	5355347_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5355347_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_117477501_117502501_95C;SPAN=7645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:10 DR:0 LR:-14.05 LO:21.05);ALT=T[chr12:117494610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	117494740	+	chr12	117537029	+	.	22	0	5355536_1	63.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5355536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:117494740(+)-12:117537029(-)__12_117526501_117551501D;SPAN=42289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:33 GQ:14.3 PL:[63.8, 0.0, 14.3] SR:0 DR:22 LR:-65.24 LO:65.24);ALT=C[chr12:117537029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	117513145	+	chr12	117537030	+	.	0	60	5355633_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5355633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_117502001_117527001_370C;SPAN=23885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:45 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:60 DR:0 LR:-178.2 LO:178.2);ALT=A[chr12:117537030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118454698	+	chr12	118456876	+	.	6	5	5358152_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=5358152_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_12_118433001_118458001_156C;SPAN=2178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:5 DR:6 LR:-3.921 LO:15.38);ALT=G[chr12:118456876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118574063	+	chr12	118575839	+	.	21	0	5358975_1	30.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5358975_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:118574063(+)-12:118575839(-)__12_118555501_118580501D;SPAN=1776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:144 GQ:30.5 PL:[30.5, 0.0, 317.6] SR:0 DR:21 LR:-30.31 LO:44.4);ALT=G[chr12:118575839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118588965	+	chr12	118590032	+	.	0	8	5358575_1	1.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5358575_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118580001_118605001_257C;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:8 DR:0 LR:-1.212 LO:14.96);ALT=T[chr12:118590032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118590215	+	chr12	118597951	+	.	3	4	5358580_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5358580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118580001_118605001_243C;SPAN=7736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:90 GQ:7.8 PL:[0.0, 7.8, 234.3] SR:4 DR:3 LR:7.878 LO:8.37);ALT=C[chr12:118597951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118599834	+	chr12	118610261	+	.	5	5	5358629_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5358629_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118604501_118629501_179C;SPAN=10427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:5 DR:5 LR:-18.6 LO:20.81);ALT=T[chr12:118610261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118610467	+	chr12	118615005	+	.	3	7	5358655_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5358655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118604501_118629501_366C;SPAN=4538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:7 DR:3 LR:-1.754 LO:15.04);ALT=T[chr12:118615005[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118615136	+	chr12	118619175	+	.	4	4	5358666_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5358666_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118604501_118629501_353C;SPAN=4039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:79 GQ:1.7 PL:[1.7, 0.0, 189.8] SR:4 DR:4 LR:-1.704 LO:13.19);ALT=T[chr12:118619175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118639269	+	chr12	118650719	+	.	2	7	5358817_1	1.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5358817_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_12_118629001_118654001_204C;SPAN=11450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:7 DR:2 LR:-1.483 LO:15.0);ALT=C[chr12:118650719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118639269	+	chr12	118651821	+	CTTAATAGTTCTGCTGATGTTGGCCTTTCCTGAGGTATTTTCTGCAAGCAGTAATCAACAAATCTCCTAAAGGAGTCTGT	3	13	5358818_1	24.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CTTAATAGTTCTGCTGATGTTGGCCTTTCCTGAGGTATTTTCTGCAAGCAGTAATCAACAAATCTCCTAAAGGAGTCTGT;MAPQ=60;MATEID=5358818_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_118629001_118654001_204C;SPAN=12552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:93 GQ:24.5 PL:[24.5, 0.0, 199.4] SR:13 DR:3 LR:-24.32 LO:32.44);ALT=C[chr12:118651821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	118693462	+	chr12	118704457	+	.	4	7	5359151_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCT;MAPQ=60;MATEID=5359151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_118678001_118703001_171C;SPAN=10995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:40 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:7 DR:4 LR:-25.47 LO:26.69);ALT=T[chr12:118704457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120639229	+	chr12	120644346	+	.	3	2	5364647_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5364647_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_12_120638001_120663001_278C;SPAN=5117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:72 GQ:6 PL:[0.0, 6.0, 184.8] SR:2 DR:3 LR:6.303 LO:6.696);ALT=G[chr12:120644346[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120639252	+	chr12	120647639	+	.	13	0	5364648_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5364648_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:120639252(+)-12:120647639(-)__12_120638001_120663001D;SPAN=8387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:75 GQ:22.7 PL:[22.7, 0.0, 158.0] SR:0 DR:13 LR:-22.59 LO:28.56);ALT=A[chr12:120647639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120882761	+	chr12	120884029	+	.	0	19	5366168_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5366168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120858501_120883501_516C;SPAN=1268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:38 GQ:39.2 PL:[52.4, 0.0, 39.2] SR:19 DR:0 LR:-52.52 LO:52.52);ALT=G[chr12:120884029[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120884632	+	chr12	120894877	+	.	0	7	5365940_1	1.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5365940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120883001_120908001_295C;SPAN=10245;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:80 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:7 DR:0 LR:-1.433 LO:13.15);ALT=G[chr12:120894877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120901927	+	chr12	120903429	+	.	4	10	5366001_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5366001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120883001_120908001_232C;SPAN=1502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:10 DR:4 LR:-23.73 LO:30.57);ALT=T[chr12:120903429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120903591	+	chr12	120907225	+	.	0	54	5366002_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=39;MATEID=5366002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120883001_120908001_247C;SPAN=3634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:79 GQ:34.7 PL:[156.8, 0.0, 34.7] SR:54 DR:0 LR:-161.2 LO:161.2);ALT=C[chr12:120907225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83360982	+	chr12	120907225	+	.	18	40	6004605_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CGGGGGTCCTCGAAGCGCACGAAGGCGAAGGGCAC;MAPQ=60;MATEID=6004605_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_15_83349001_83374001_26C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:30 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:40 DR:18 LR:-148.5 LO:148.5);ALT=]chr15:83360982]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr12	120934030	+	chr12	120935873	+	.	41	0	5365557_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5365557_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:120934030(+)-12:120935873(-)__12_120932001_120957001D;SPAN=1843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:92 GQ:99 PL:[110.6, 0.0, 110.6] SR:0 DR:41 LR:-110.4 LO:110.4);ALT=C[chr12:120935873[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	120934357	+	chr12	120935874	+	.	7	107	5365559_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5365559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_120932001_120957001_369C;SPAN=1517;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:93 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:107 DR:7 LR:-333.4 LO:333.4);ALT=G[chr12:120935874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121017401	+	chr12	121018916	+	.	0	7	5365769_1	0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=5365769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121005501_121030501_219C;SPAN=1515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:97 GQ:3 PL:[0.0, 3.0, 240.9] SR:7 DR:0 LR:3.173 LO:12.54);ALT=C[chr12:121018916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121017727	+	chr12	121018918	+	.	0	21	5365771_1	42.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5365771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121005501_121030501_370C;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:99 GQ:42.5 PL:[42.5, 0.0, 197.6] SR:21 DR:0 LR:-42.5 LO:48.2);ALT=C[chr12:121018918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121163734	+	chr12	121164827	+	.	37	9	5366604_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5366604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121152501_121177501_365C;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:78 GQ:87.8 PL:[101.0, 0.0, 87.8] SR:9 DR:37 LR:-101.0 LO:101.0);ALT=G[chr12:121164827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121163746	+	chr12	121174785	+	.	8	0	5366605_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5366605_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:121163746(+)-12:121174785(-)__12_121152501_121177501D;SPAN=11039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-2.025 LO:15.08);ALT=G[chr12:121174785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121164996	+	chr12	121174786	+	.	0	17	5366608_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CAGGTGA;MAPQ=60;MATEID=5366608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121152501_121177501_98C;SPAN=9790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:96 GQ:30.2 PL:[30.2, 0.0, 201.8] SR:17 DR:0 LR:-30.11 LO:37.52);ALT=A[chr12:121174786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121448731	+	chr12	121454131	+	GAGGCTCGGTTGGGAGGTTGACAACTGGCTATTTGCAGC	5	9	5367130_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=GAGGCTCGGTTGGGAGGTTGACAACTGGCTATTTGCAGC;MAPQ=60;MATEID=5367130_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_121446501_121471501_71C;SPAN=5400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:81 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:9 DR:5 LR:-14.37 LO:22.89);ALT=T[chr12:121454131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121712391	+	chr12	121734438	+	.	7	2	5368538_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCTG;MAPQ=60;MATEID=5368538_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121691501_121716501_219C;SPAN=22047;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:36 GQ:13.4 PL:[13.4, 0.0, 72.8] SR:2 DR:7 LR:-13.35 LO:15.77);ALT=G[chr12:121734438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121746496	+	chr12	121747504	+	.	8	6	5368715_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5368715_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_121740501_121765501_223C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:6 DR:8 LR:-8.677 LO:21.71);ALT=T[chr12:121747504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	121785687	+	chr12	121789936	+	.	13	28	5368964_1	94.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=5368964_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_121789501_121814501_11C;SPAN=4249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:43 GQ:8.3 PL:[94.1, 0.0, 8.3] SR:28 DR:13 LR:-97.88 LO:97.88);ALT=G[chr12:121789936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122064959	+	chr12	122078946	+	.	14	7	5369907_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=5369907_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122059001_122084001_291C;SPAN=13987;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:77 GQ:25.4 PL:[25.4, 0.0, 160.7] SR:7 DR:14 LR:-25.35 LO:31.08);ALT=G[chr12:122078946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122219144	+	chr12	122231497	+	.	8	0	5370602_1	9.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5370602_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:122219144(+)-12:122231497(-)__12_122206001_122231001D;SPAN=12353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=C[chr12:122231497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122326900	+	chr12	122332645	+	.	0	43	5370852_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5370852_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122328501_122353501_60C;SPAN=5745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:38 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:43 DR:0 LR:-125.4 LO:125.4);ALT=C[chr12:122332645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122326944	+	chr12	122337539	+	.	13	0	5370853_1	29.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5370853_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:122326944(+)-12:122337539(-)__12_122328501_122353501D;SPAN=10595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:0 DR:13 LR:-28.83 LO:30.91);ALT=G[chr12:122337539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122701418	+	chr12	122702812	+	.	0	4	5372085_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5372085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122696001_122721001_306C;SPAN=1394;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:72 GQ:6 PL:[0.0, 6.0, 184.8] SR:4 DR:0 LR:6.303 LO:6.696);ALT=T[chr12:122702812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122702947	+	chr12	122709059	+	.	0	15	5372096_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5372096_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122696001_122721001_230C;SPAN=6112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:83 GQ:27.2 PL:[27.2, 0.0, 172.4] SR:15 DR:0 LR:-27.03 LO:33.26);ALT=G[chr12:122709059[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122702989	+	chr12	122710507	+	.	15	0	5372097_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5372097_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:122702989(+)-12:122710507(-)__12_122696001_122721001D;SPAN=7518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:74 GQ:29.6 PL:[29.6, 0.0, 148.4] SR:0 DR:15 LR:-29.47 LO:34.09);ALT=G[chr12:122710507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122709194	+	chr12	122710508	+	.	13	2	5372119_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTACCTG;MAPQ=60;MATEID=5372119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122696001_122721001_180C;SPAN=1314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:72 GQ:26.9 PL:[26.9, 0.0, 145.7] SR:2 DR:13 LR:-26.71 LO:31.54);ALT=G[chr12:122710508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122748748	+	chr12	122750853	+	.	3	3	5372160_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5372160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122745001_122770001_137C;SPAN=2105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:83 GQ:5.7 PL:[0.0, 5.7, 211.2] SR:3 DR:3 LR:5.982 LO:8.55);ALT=T[chr12:122750853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122862688	-	chr12	122863813	+	.	8	0	5372640_1	1.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5372640_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:122862688(-)-12:122863813(-)__12_122843001_122868001D;SPAN=1125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:0 DR:8 LR:-0.9411 LO:14.92);ALT=[chr12:122863813[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	122991471	+	chr12	122992764	+	.	3	2	5372973_1	0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5372973_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_122990001_123015001_325C;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:78 GQ:7.8 PL:[0.0, 7.8, 204.6] SR:2 DR:3 LR:7.928 LO:6.554);ALT=C[chr12:122992764[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122992999	+	chr12	122995656	+	.	4	11	5372983_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5372983_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122990001_123015001_95C;SPAN=2657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:11 DR:4 LR:-26.49 LO:33.08);ALT=T[chr12:122995656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122999775	+	chr12	123003386	+	GACTCCTACTCCTTGTCCTACTCCTGCTTCTAGTCCTATGCCTGTGTCTTGATCTTGAGCGGGAACGAGACCTGATCCGCCGTTTTCTTTCCCTGCTTCTGGATCTCGATTTCTTCCTCTCTCTGCTTCTGGATCTCGATTTCTTCCGCTCCCTACTCCTGGATCGAGACTTCTTCCGCTCCCTGCTTCTACTACGATGGCGT	0	30	5373014_1	75.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GACTCCTACTCCTTGTCCTACTCCTGCTTCTAGTCCTATGCCTGTGTCTTGATCTTGAGCGGGAACGAGACCTGATCCGCCGTTTTCTTTCCCTGCTTCTGGATCTCGATTTCTTCCTCTCTCTGCTTCTGGATCTCGATTTCTTCCGCTCCCTACTCCTGGATCGAGACTTCTTCCGCTCCCTGCTTCTACTACGATGGCGT;MAPQ=60;MATEID=5373014_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_122990001_123015001_92C;SPAN=3611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:88 GQ:75.2 PL:[75.2, 0.0, 137.9] SR:30 DR:0 LR:-75.19 LO:76.21);ALT=C[chr12:123003386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	122999775	+	chr12	123001774	+	.	8	14	5373013_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5373013_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_12_122990001_123015001_92C;SPAN=1999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:89 GQ:45.2 PL:[45.2, 0.0, 170.6] SR:14 DR:8 LR:-45.21 LO:49.32);ALT=C[chr12:123001774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123001979	+	chr12	123003386	+	.	13	15	5373019_1	53.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5373019_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_122990001_123015001_92C;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:82 GQ:53.9 PL:[53.9, 0.0, 143.0] SR:15 DR:13 LR:-53.71 LO:56.04);ALT=T[chr12:123003386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123003578	+	chr12	123005931	+	.	2	5	5373023_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=5373023_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_12_122990001_123015001_91C;SPAN=2353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:78 GQ:2 PL:[2.0, 0.0, 186.8] SR:5 DR:2 LR:-1.975 LO:13.23);ALT=T[chr12:123005931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123003578	+	chr12	123006690	+	CTTTGCTTCTGCTCCGGCTCCTGTGTTTTCTTCCTTCATTAT	3	20	5373024_1	48.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTTTGCTTCTGCTCCGGCTCCTGTGTTTTCTTCCTTCATTAT;MAPQ=60;MATEID=5373024_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_122990001_123015001_91C;SPAN=3112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:90 GQ:48.2 PL:[48.2, 0.0, 170.3] SR:20 DR:3 LR:-48.24 LO:52.06);ALT=T[chr12:123006690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123006847	+	chr12	123011394	+	.	31	10	5373036_1	85.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5373036_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_122990001_123015001_65C;SPAN=4547;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:101 GQ:85.1 PL:[85.1, 0.0, 157.7] SR:10 DR:31 LR:-84.87 LO:86.14);ALT=C[chr12:123011394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123218034	-	chr12	123219535	+	.	3	5	5373907_1	0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=ATTACAGGTGT;MAPQ=60;MATEID=5373907_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_123210501_123235501_123C;SPAN=1501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:98 GQ:6.6 PL:[0.0, 6.6, 250.8] SR:5 DR:3 LR:6.745 LO:10.3);ALT=[chr12:123219535[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr12	123237484	+	chr20	32834328	-	.	24	0	6985526_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6985526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123237484(+)-20:32834328(+)__20_32830001_32855001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:73 GQ:59.6 PL:[59.6, 0.0, 115.7] SR:0 DR:24 LR:-59.45 LO:60.5);ALT=G]chr20:32834328];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr12	123238354	+	chr12	123247390	+	AAATATTTGTGAATTGTAAATGCTGTATGTATTCGCATCTTGGAAACTTTCAGAAAAATCTGAAGATACAGGACAGTAAAAGGTCTGTTCATTACCAACAG	2	23	5374071_1	56.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TGCAAAGGAGACCCAAGGAACAGTGCCAAGTTAGATGCCGATTACCCACTTCGAGTCCTTTATTGTGGAGAAATATTTGTGAATTGTAAATGCTGTATGTATTCGCATCTTGGAAACTTTCAGAAAAATCTGAAGATACAGGACAGTAAAAGG;INSERTION=AAATATTTGTGAATTGTAAATGCTGTATGTATTCGCATCTTGGAAACTTTCAGAAAAATCTGAAGATACAGGACAGTAAAAGGTCTGTTCATTACCAACAG;MAPQ=38;MATEID=5374071_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_123235001_123260001_267C;SECONDARY;SPAN=9036;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:96 GQ:56.6 PL:[56.6, 0.0, 175.4] SR:23 DR:2 LR:-56.52 LO:59.96);ALT=G[chr12:123247390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123252151	+	chr12	123253328	+	.	3	7	5374106_1	16.0	.	DISC_MAPQ=38;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=5374106_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_12_123235001_123260001_6C;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:7 DR:3 LR:-16.21 LO:21.62);ALT=G[chr12:123253328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123459879	+	chr12	123461198	+	.	8	0	5374728_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5374728_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123459879(+)-12:123461198(-)__12_123455501_123480501D;SPAN=1319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=G[chr12:123461198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123715041	+	chr12	123717620	+	.	10	0	5375531_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5375531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123715041(+)-12:123717620(-)__12_123700501_123725501D;SPAN=2579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.34 LO:20.42);ALT=T[chr12:123717620[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123746351	+	chr12	123749742	+	.	4	7	5375934_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5375934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_123725001_123750001_291C;SPAN=3391;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:93 GQ:4.7 PL:[4.7, 0.0, 219.2] SR:7 DR:4 LR:-4.513 LO:17.32);ALT=C[chr12:123749742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123749894	+	chr12	123752736	+	.	19	0	5375945_1	52.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5375945_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123749894(+)-12:123752736(-)__12_123725001_123750001D;SPAN=2842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:39 GQ:42.2 PL:[52.1, 0.0, 42.2] SR:0 DR:19 LR:-52.2 LO:52.2);ALT=A[chr12:123752736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123900468	+	chr12	123907589	+	.	3	2	5376468_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=5376468_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_123896501_123921501_314C;SPAN=7121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:89 GQ:10.8 PL:[0.0, 10.8, 237.6] SR:2 DR:3 LR:10.91 LO:6.32);ALT=C[chr12:123907589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123915208	+	chr12	123920625	+	.	5	12	5376520_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCACCT;MAPQ=60;MATEID=5376520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_123896501_123921501_160C;SPAN=5417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:104 GQ:21.5 PL:[21.5, 0.0, 229.4] SR:12 DR:5 LR:-21.34 LO:31.64);ALT=T[chr12:123920625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	123942780	+	chr12	123950082	+	.	14	0	5377066_1	34.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5377066_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:123942780(+)-12:123950082(-)__12_123921001_123946001D;SPAN=7302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:45 GQ:34.1 PL:[34.1, 0.0, 73.7] SR:0 DR:14 LR:-34.02 LO:34.88);ALT=T[chr12:123950082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124069363	+	chr12	124071292	+	.	31	57	5376855_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5376855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124068001_124093001_292C;SPAN=1929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:116 GQ:80.9 PL:[199.7, 0.0, 80.9] SR:57 DR:31 LR:-202.3 LO:202.3);ALT=G[chr12:124071292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124074996	+	chr12	124081152	+	.	8	5	5376871_1	16.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=5376871_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124068001_124093001_338C;SPAN=6156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:5 DR:8 LR:-16.31 LO:25.12);ALT=A[chr12:124081152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124086769	+	chr12	124090475	+	.	8	0	5376923_1	6.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5376923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:124086769(+)-12:124090475(-)__12_124068001_124093001D;SPAN=3706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=G[chr12:124090475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124115082	+	chr12	124116891	+	.	0	12	5377260_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5377260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124092501_124117501_136C;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:72 GQ:20.3 PL:[20.3, 0.0, 152.3] SR:12 DR:0 LR:-20.11 LO:26.14);ALT=T[chr12:124116891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124116994	+	chr12	124118092	+	.	14	6	5377268_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5377268_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124092501_124117501_100C;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:23 GQ:13.7 PL:[40.1, 0.0, 13.7] SR:6 DR:14 LR:-40.55 LO:40.55);ALT=C[chr12:124118092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124118470	+	chr12	124129998	+	.	11	0	5377278_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5377278_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:124118470(+)-12:124129998(-)__12_124117001_124142001D;SPAN=11528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:99 GQ:9.5 PL:[9.5, 0.0, 230.6] SR:0 DR:11 LR:-9.49 LO:21.86);ALT=T[chr12:124129998[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	124130108	+	chr12	124132508	+	.	0	8	5377335_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5377335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_124117001_124142001_236C;SPAN=2400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:8 DR:0 LR:-5.276 LO:15.61);ALT=G[chr12:124132508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	131131938	+	chr12	131133868	+	.	90	59	5396285_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=5396285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_131124001_131149001_414C;SPAN=1930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:128 DP:32 GQ:34.5 PL:[379.5, 34.5, 0.0] SR:59 DR:90 LR:-379.6 LO:379.6);ALT=C[chr12:131133868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	132262877	+	chr12	132271006	+	.	4	2	5399335_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=5399335_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_132251001_132276001_268C;SPAN=8129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:83 GQ:9 PL:[0.0, 9.0, 217.8] SR:2 DR:4 LR:9.283 LO:6.444);ALT=T[chr12:132271006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133067447	+	chr12	133084737	+	.	18	45	5401719_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5401719_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_133084001_133109001_158C;SPAN=17290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:35 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:45 DR:18 LR:-151.8 LO:151.8);ALT=G[chr12:133084737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133067489	+	chr12	133085747	+	.	11	0	5401720_1	22.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=5401720_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:133067489(+)-12:133085747(-)__12_133084001_133109001D;SPAN=18258;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:52 GQ:22.4 PL:[22.4, 0.0, 101.6] SR:0 DR:11 LR:-22.22 LO:25.23);ALT=C[chr12:133085747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133141112	+	chr12	133344211	-	.	2	8	5401818_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTGGAGACGGAGTCTC;MAPQ=60;MATEID=5401818_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_12_133133001_133158001_66C;SPAN=203099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:8 DR:2 LR:-21.31 LO:22.09);ALT=C]chr12:133344211];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr12	133175151	+	chr12	133174003	+	.	32	0	5401927_1	87.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5401927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:133174003(-)-12:133175151(+)__12_133157501_133182501D;SPAN=1148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:68 GQ:77.3 PL:[87.2, 0.0, 77.3] SR:0 DR:32 LR:-87.24 LO:87.24);ALT=]chr12:133175151]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr12	133264323	+	chr12	133266845	+	.	20	0	5402494_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5402494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:133264323(+)-12:133266845(-)__12_133255501_133280501D;SPAN=2522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:60 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:0 DR:20 LR:-49.76 LO:50.57);ALT=G[chr12:133266845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133264378	+	chr12	133272469	+	TGGCATTTTGTCAGCACTTGGGAACTTCCTGGCCCAGATGATTGAGAAGAAGCGGAAAAAAGAAAACTCTAGAAGTCTGGATGTCGGTGGGCCTCTGAGATATGCCGTTTACG	0	20	5402496_1	48.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=TGGCATTTTGTCAGCACTTGGGAACTTCCTGGCCCAGATGATTGAGAAGAAGCGGAAAAAAGAAAACTCTAGAAGTCTGGATGTCGGTGGGCCTCTGAGATATGCCGTTTACG;MAPQ=60;MATEID=5402496_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_12_133255501_133280501_334C;SPAN=8091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:65 GQ:48.5 PL:[48.5, 0.0, 107.9] SR:20 DR:0 LR:-48.41 LO:49.71);ALT=G[chr12:133272469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	133331721	+	chr12	133338202	+	.	0	10	5402696_1	17.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=5402696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_133329001_133354001_170C;SPAN=6481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:10 DR:0 LR:-17.84 LO:22.11);ALT=T[chr12:133338202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	19318687	-	chr13	19319694	+	.	9	0	5405014_1	5.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=5405014_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:19318687(-)-13:19319694(-)__13_19306001_19331001D;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:0 DR:9 LR:-5.597 LO:17.5);ALT=[chr13:19319694[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	19694137	+	chr13	19692860	+	.	18	0	5406423_1	40.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5406423_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:19692860(-)-13:19694137(+)__13_19673501_19698501D;SPAN=1277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:71 GQ:40.4 PL:[40.4, 0.0, 129.5] SR:0 DR:18 LR:-40.18 LO:42.93);ALT=]chr13:19694137]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	19766998	+	chr13	21769412	-	.	13	0	5413591_1	32.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5413591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:19766998(+)-13:21769412(+)__13_21756001_21781001D;SPAN=2002414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:40 GQ:32 PL:[32.0, 0.0, 65.0] SR:0 DR:13 LR:-32.08 LO:32.69);ALT=G]chr13:21769412];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr13	20426330	+	chr13	20436537	+	.	0	8	5408838_1	14.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=5408838_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_20433001_20458001_10C;SPAN=10207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:8 DR:0 LR:-14.49 LO:17.76);ALT=C[chr13:20436537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	20426361	+	chr13	20437588	+	.	14	0	5409116_1	37.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5409116_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:20426361(+)-13:20437588(-)__13_20408501_20433501D;SPAN=11227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:32 GQ:37.7 PL:[37.7, 0.0, 37.7] SR:0 DR:14 LR:-37.54 LO:37.55);ALT=C[chr13:20437588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	20532982	+	chr13	20534097	+	.	0	7	5409143_1	4.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5409143_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_20531001_20556001_289C;SPAN=1115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:70 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:7 DR:0 LR:-4.142 LO:13.57);ALT=G[chr13:20534097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	20533251	+	chr13	20567200	+	.	9	0	5409468_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5409468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:20533251(+)-13:20567200(-)__13_20555501_20580501D;SPAN=33949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:0 DR:9 LR:-15.08 LO:19.6);ALT=G[chr13:20567200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21063682	+	chr13	21099892	+	.	17	0	5411083_1	48.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5411083_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:21063682(+)-13:21099892(-)__13_21094501_21119501D;SPAN=36210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:27 GQ:15.8 PL:[48.8, 0.0, 15.8] SR:0 DR:17 LR:-49.67 LO:49.67);ALT=T[chr13:21099892[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21086692	+	chr13	21099893	+	.	10	3	5411229_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=5411229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_21070001_21095001_223C;SPAN=13201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:44 GQ:24.5 PL:[24.5, 0.0, 80.6] SR:3 DR:10 LR:-24.39 LO:26.15);ALT=G[chr13:21099893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21436998	+	chr13	21442735	+	.	0	12	5412168_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5412168_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_21437501_21462501_212C;SPAN=5737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:37 GQ:29.6 PL:[29.6, 0.0, 59.3] SR:12 DR:0 LR:-29.59 LO:30.16);ALT=C[chr13:21442735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21437292	+	chr13	21476807	+	.	28	0	5412244_1	81.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5412244_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:21437292(+)-13:21476807(-)__13_21462001_21487001D;SPAN=39515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:41 GQ:15.5 PL:[81.5, 0.0, 15.5] SR:0 DR:28 LR:-83.57 LO:83.57);ALT=A[chr13:21476807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21442841	+	chr13	21476808	+	.	7	3	5412245_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5412245_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_21462001_21487001_21C;SPAN=33967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:3 DR:7 LR:-15.3 LO:18.03);ALT=C[chr13:21476808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21715134	+	chr13	21719230	+	.	4	6	5413143_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5413143_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_21707001_21732001_322C;SPAN=4096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:110 GQ:0 PL:[0.0, 0.0, 267.3] SR:6 DR:4 LR:0.0927 LO:16.63);ALT=G[chr13:21719230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21715135	+	chr13	21720943	+	.	21	125	5413144_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5413144_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_21707001_21732001_270C;SPAN=5808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:119 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:125 DR:21 LR:-415.9 LO:415.9);ALT=G[chr13:21720943[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21872412	+	chr13	21875556	+	.	8	0	5413724_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5413724_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:21872412(+)-13:21875556(-)__13_21854001_21879001D;SPAN=3144;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=A[chr13:21875556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	21904830	+	chr13	21918882	+	.	9	0	5413845_1	6.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5413845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:21904830(+)-13:21918882(-)__13_21903001_21928001D;SPAN=14052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:0 DR:9 LR:-6.139 LO:17.59);ALT=A[chr13:21918882[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	45168946	-	chr17	38804024	+	.	9	0	6393081_1	12.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=6393081_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:45168946(-)-17:38804024(-)__17_38783501_38808501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=[chr17:38804024[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr13	45694858	+	chr13	45710866	+	ACTCAAGGAAGGACTG	0	17	5480815_1	30.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;INSERTION=ACTCAAGGAAGGACTG;MAPQ=60;MATEID=5480815_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_45692501_45717501_331C;SECONDARY;SPAN=16008;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:94 GQ:30.8 PL:[30.8, 0.0, 195.8] SR:17 DR:0 LR:-30.65 LO:37.69);ALT=T[chr13:45710866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	45841513	+	chr13	45857576	+	.	5	5	5481418_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5481418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_45839501_45864501_170C;SPAN=16063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:96 GQ:0.5 PL:[0.5, 0.0, 231.5] SR:5 DR:5 LR:-0.3992 LO:14.85);ALT=T[chr13:45857576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	45911634	+	chr13	45912793	+	.	19	0	5481685_1	13.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=5481685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:45911634(+)-13:45912793(-)__13_45888501_45913501D;SPAN=1159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:184 GQ:13 PL:[13.0, 0.0, 432.2] SR:0 DR:19 LR:-12.87 LO:37.12);ALT=A[chr13:45912793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46701858	+	chr13	46704949	+	.	14	6	5484045_1	37.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5484045_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46697001_46722001_137C;SPAN=3091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:94 GQ:37.4 PL:[37.4, 0.0, 189.2] SR:6 DR:14 LR:-37.25 LO:43.16);ALT=T[chr13:46704949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46705067	+	chr13	46708261	+	AGGGT	4	5	5484064_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AGGGT;MAPQ=60;MATEID=5484064_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_46697001_46722001_136C;SPAN=3194;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:96 GQ:3.8 PL:[3.8, 0.0, 228.2] SR:5 DR:4 LR:-3.7 LO:17.19);ALT=T[chr13:46708261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46708387	+	chr13	46716424	+	.	3	5	5484076_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCT;MAPQ=60;MATEID=5484076_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_46697001_46722001_87C;SPAN=8037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:75 GQ:2.9 PL:[2.9, 0.0, 177.8] SR:5 DR:3 LR:-2.788 LO:13.35);ALT=T[chr13:46716424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46717542	+	chr13	46718577	+	.	0	7	5484101_1	0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5484101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46697001_46722001_85C;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:7 DR:0 LR:2.902 LO:12.57);ALT=G[chr13:46718577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46721239	+	chr13	46722486	+	.	22	17	5484110_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5484110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46697001_46722001_283C;SPAN=1247;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:59 GQ:53.3 PL:[89.6, 0.0, 53.3] SR:17 DR:22 LR:-90.14 LO:90.14);ALT=C[chr13:46722486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46721268	+	chr13	46725069	+	.	16	0	5484111_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5484111_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:46721268(+)-13:46725069(-)__13_46697001_46722001D;SPAN=3801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:53 GQ:38.6 PL:[38.6, 0.0, 88.1] SR:0 DR:16 LR:-38.46 LO:39.6);ALT=G[chr13:46725069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46722584	+	chr13	46725070	+	.	0	27	5483734_1	64.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5483734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46721501_46746501_259C;SPAN=2486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:93 GQ:64.1 PL:[64.1, 0.0, 159.8] SR:27 DR:0 LR:-63.93 LO:66.28);ALT=T[chr13:46725070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46725215	+	chr13	46726915	+	.	5	12	5483741_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5483741_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_46721501_46746501_60C;SPAN=1700;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:101 GQ:29 PL:[29.0, 0.0, 213.8] SR:12 DR:5 LR:-28.75 LO:37.11);ALT=T[chr13:46726915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46727084	+	chr13	46728939	+	.	5	8	5483744_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTGA;MAPQ=60;MATEID=5483744_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_46721501_46746501_60C;SPAN=1855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:76 GQ:19.1 PL:[19.1, 0.0, 164.3] SR:8 DR:5 LR:-19.02 LO:25.83);ALT=A[chr13:46728939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46727105	+	chr13	46730572	+	.	9	0	5483745_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5483745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:46727105(+)-13:46730572(-)__13_46721501_46746501D;SPAN=3467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=T[chr13:46730572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46729022	+	chr13	46732961	+	AAAGGACAATGCCATCTCCAACAGCATTAAAGAGATCATTCGTGTTTGGGTTCATTGGGATGACATGCCGACAATCAGGATCATTTTCCAGGGCTTTGTTTATCCAGTTGACAAAGGCATACTTTTCTTCCTCTGAATAGGAGTGTTGGGTGCCAACGCTAGACTGCTCTGAAGTACCACCGATTGCACAAATCCCTTCCTTCTTATTGATTGCTTTTCTAAAGGTCTTGGCAACATCTGTGCTTTTTAGGCCATGGAAAAT	0	49	5483750_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AAAGGACAATGCCATCTCCAACAGCATTAAAGAGATCATTCGTGTTTGGGTTCATTGGGATGACATGCCGACAATCAGGATCATTTTCCAGGGCTTTGTTTATCCAGTTGACAAAGGCATACTTTTCTTCCTCTGAATAGGAGTGTTGGGTGCCAACGCTAGACTGCTCTGAAGTACCACCGATTGCACAAATCCCTTCCTTCTTATTGATTGCTTTTCTAAAGGTCTTGGCAACATCTGTGCTTTTTAGGCCATGGAAAAT;MAPQ=60;MATEID=5483750_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_46721501_46746501_37C;SPAN=3939;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:93 GQ:87.2 PL:[136.7, 0.0, 87.2] SR:49 DR:0 LR:-137.1 LO:137.1);ALT=C[chr13:46732961[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46730708	+	chr13	46732657	+	.	16	10	5483753_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=5483753_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_46721501_46746501_37C;SPAN=1949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:80 GQ:47.6 PL:[47.6, 0.0, 146.6] SR:10 DR:16 LR:-47.65 LO:50.45);ALT=G[chr13:46732657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	46733823	+	chr13	46756246	+	.	72	18	5483770_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5483770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_46721501_46746501_155C;SPAN=22423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:48 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:18 DR:72 LR:-237.7 LO:237.7);ALT=T[chr13:46756246[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47345633	+	chr13	47351590	+	.	8	86	5485714_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5485714_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_47334001_47359001_362C;SPAN=5957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:113 GQ:5.9 PL:[266.6, 0.0, 5.9] SR:86 DR:8 LR:-281.3 LO:281.3);ALT=T[chr13:47351590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47351760	+	chr13	47354069	+	.	0	13	5485729_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5485729_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_47334001_47359001_20C;SPAN=2309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:13 DR:0 LR:-19.34 LO:27.64);ALT=T[chr13:47354069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47354168	+	chr13	47355631	+	.	0	7	5485733_1	4.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5485733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_47334001_47359001_221C;SPAN=1463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:70 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:7 DR:0 LR:-4.142 LO:13.57);ALT=A[chr13:47355631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47355752	+	chr13	47356802	+	.	3	6	5485738_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5485738_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_47334001_47359001_17C;SPAN=1050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:6 DR:3 LR:-7.764 LO:17.89);ALT=T[chr13:47356802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47356926	+	chr13	47358385	+	.	5	16	5485742_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=5485742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_47334001_47359001_16C;SPAN=1459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:81 GQ:47.6 PL:[47.6, 0.0, 146.6] SR:16 DR:5 LR:-47.38 LO:50.32);ALT=C[chr13:47358385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47358489	+	chr13	47365481	+	GAGCCAATACAGTGCAGGGCACTTTCCTGTTTCTGCCTTTGGTGGTAAGTAGACAGCAAATTTCATTTTGCAGTTTAGTTCAACA	0	140	5485758_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GAGCCAATACAGTGCAGGGCACTTTCCTGTTTCTGCCTTTGGTGGTAAGTAGACAGCAAATTTCATTTTGCAGTTTAGTTCAACA;MAPQ=60;MATEID=5485758_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_47358501_47383501_189C;SPAN=6992;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:79 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:140 DR:0 LR:-415.9 LO:415.9);ALT=A[chr13:47365481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47358533	+	chr13	47371239	+	.	29	0	5485760_1	62.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5485760_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:47358533(+)-13:47371239(-)__13_47358501_47383501D;SPAN=12706;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:123 GQ:62.6 PL:[62.6, 0.0, 234.2] SR:0 DR:29 LR:-62.41 LO:68.09);ALT=T[chr13:47371239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47361294	+	chr13	47371239	+	.	79	0	5485768_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5485768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:47361294(+)-13:47371239(-)__13_47358501_47383501D;SPAN=9945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:125 GQ:75.2 PL:[227.0, 0.0, 75.2] SR:0 DR:79 LR:-231.0 LO:231.0);ALT=A[chr13:47371239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	47365603	+	chr13	47371239	+	.	42	0	5485783_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5485783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:47365603(+)-13:47371239(-)__13_47358501_47383501D;SPAN=5636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:118 GQ:99 PL:[106.7, 0.0, 179.3] SR:0 DR:42 LR:-106.7 LO:107.7);ALT=A[chr13:47371239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48571144	+	chr13	48575343	+	.	9	0	5488763_1	2.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=5488763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:48571144(+)-13:48575343(-)__13_48559001_48584001D;SPAN=4199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=A[chr13:48575343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48611986	+	chr13	48615054	+	.	9	0	5489019_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5489019_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:48611986(+)-13:48615054(-)__13_48608001_48633001D;SPAN=3068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:0 DR:9 LR:-10.2 LO:18.38);ALT=A[chr13:48615054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48654113	+	chr13	48655780	+	.	0	7	5488975_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5488975_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48632501_48657501_313C;SPAN=1667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:7 DR:0 LR:0.4634 LO:12.88);ALT=T[chr13:48655780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48660591	+	chr13	48664486	+	.	2	8	5489093_1	11.0	.	DISC_MAPQ=30;EVDNC=TSI_L;HOMSEQ=ACCTG;MAPQ=60;MATEID=5489093_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_13_48657001_48682001_145C;SPAN=3895;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:8 DR:2 LR:-11.34 LO:20.42);ALT=G[chr13:48664486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48660620	+	chr13	48669161	+	.	16	0	5489095_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5489095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:48660620(+)-13:48669161(-)__13_48657001_48682001D;SPAN=8541;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:90 GQ:28.4 PL:[28.4, 0.0, 190.1] SR:0 DR:16 LR:-28.43 LO:35.35);ALT=T[chr13:48669161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48664557	+	chr13	48669089	+	.	7	6	5489109_1	2.0	.	DISC_MAPQ=56;EVDNC=TSI_L;HOMSEQ=CCTA;MAPQ=60;MATEID=5489109_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_48657001_48682001_145C;SPAN=4532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:6 DR:7 LR:-1.804 LO:16.9);ALT=A[chr13:48669089[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48807614	+	chr13	48827942	+	.	0	170	5489475_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5489475_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48804001_48829001_210C;SPAN=20328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:184 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:170 DR:0 LR:-544.6 LO:544.6);ALT=G[chr13:48827942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48828072	+	chr13	48830313	+	.	15	22	5489531_1	89.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=5489531_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48828501_48853501_100C;SPAN=2241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:48 GQ:26.6 PL:[89.3, 0.0, 26.6] SR:22 DR:15 LR:-91.16 LO:91.16);ALT=A[chr13:48830313[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48830519	+	chr13	48832931	+	AAACTTACAGCCTATTTAGATCTTAACCTGGATAAGTGCTATGTGATCCCTCTGAACACTTCCATTGTTATGCCACCCAGAAACCTACTGGAGTTACTTATTAACATCA	12	40	5489540_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAACTTACAGCCTATTTAGATCTTAACCTGGATAAGTGCTATGTGATCCCTCTGAACACTTCCATTGTTATGCCACCCAGAAACCTACTGGAGTTACTTATTAACATCA;MAPQ=60;MATEID=5489540_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_48828501_48853501_180C;SPAN=2412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:109 GQ:99 PL:[125.6, 0.0, 138.8] SR:40 DR:12 LR:-125.6 LO:125.7);ALT=G[chr13:48832931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48830519	+	chr13	48832260	+	.	19	18	5489539_1	77.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5489539_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_13_48828501_48853501_180C;SPAN=1741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:93 GQ:77.3 PL:[77.3, 0.0, 146.6] SR:18 DR:19 LR:-77.14 LO:78.38);ALT=G[chr13:48832260[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48833086	+	chr13	48835273	+	.	18	57	5489544_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=5489544_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48828501_48853501_303C;SPAN=2187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:102 GQ:35.3 PL:[210.2, 0.0, 35.3] SR:57 DR:18 LR:-216.9 LO:216.9);ALT=A[chr13:48835273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	48878186	+	chr13	48881414	+	.	0	17	5490009_1	32.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5490009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_48877501_48902501_262C;SPAN=3228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:86 GQ:32.9 PL:[32.9, 0.0, 174.8] SR:17 DR:0 LR:-32.82 LO:38.43);ALT=G[chr13:48881414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49533321	+	chr13	49536621	+	.	10	0	5491619_1	16.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5491619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:49533321(+)-13:49536621(-)__13_49514501_49539501D;SPAN=3300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:61 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.48 LO:21.7);ALT=C[chr13:49536621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49822257	+	chr13	49829973	+	CAGATACCAAGGCTTTCTAAAGTCAACCTTTTCACTCTGCTCAGCCTCTGGATGGAGCTCTTTCCAGCAGAAGCCCAGCGGCAAAAATCTC	0	17	5492331_1	31.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAGATACCAAGGCTTTCTAAAGTCAACCTTTTCACTCTGCTCAGCCTCTGGATGGAGCTCTTTCCAGCAGAAGCCCAGCGGCAAAAATCTC;MAPQ=60;MATEID=5492331_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_49808501_49833501_22C;SPAN=7716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:91 GQ:31.7 PL:[31.7, 0.0, 186.8] SR:17 DR:0 LR:-31.46 LO:37.96);ALT=T[chr13:49829973[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	49951414	+	chr13	49953863	+	.	30	22	5492649_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AAACAAAAACAGT;MAPQ=60;MATEID=5492649_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_49931001_49956001_136C;SPAN=2449;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:67 GQ:57.8 PL:[104.0, 0.0, 57.8] SR:22 DR:30 LR:-104.7 LO:104.7);ALT=T[chr13:49953863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50070235	+	chr13	50080770	+	.	22	8	5493113_1	68.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGT;MAPQ=60;MATEID=5493113_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_13_50078001_50103001_87C;SPAN=10535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:39 GQ:25.7 PL:[68.6, 0.0, 25.7] SR:8 DR:22 LR:-69.71 LO:69.71);ALT=T[chr13:50080770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50070243	+	chr13	50087193	+	.	11	0	5493115_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5493115_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:50070243(+)-13:50087193(-)__13_50078001_50103001D;SPAN=16950;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:52 GQ:22.4 PL:[22.4, 0.0, 101.6] SR:0 DR:11 LR:-22.22 LO:25.23);ALT=G[chr13:50087193[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50080892	+	chr13	50087194	+	.	0	10	5493135_1	8.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5493135_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_50078001_50103001_343C;SPAN=6302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:10 DR:0 LR:-8.627 LO:19.88);ALT=G[chr13:50087194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50087302	+	chr13	50092153	+	.	2	9	5493155_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5493155_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_50078001_50103001_363C;SPAN=4851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:9 DR:2 LR:-15.45 LO:23.15);ALT=G[chr13:50092153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50141492	+	chr13	50159621	+	.	9	0	5493491_1	19.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5493491_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:50141492(+)-13:50159621(-)__13_50151501_50176501D;SPAN=18129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:0 DR:9 LR:-19.68 LO:21.27);ALT=A[chr13:50159621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50202742	+	chr13	50204563	+	.	12	0	5493398_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5493398_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:50202742(+)-13:50204563(-)__13_50200501_50225501D;SPAN=1821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:83 GQ:17.3 PL:[17.3, 0.0, 182.3] SR:0 DR:12 LR:-17.13 LO:25.33);ALT=T[chr13:50204563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50235345	+	chr13	50265389	+	.	29	33	5493823_1	99.0	.	DISC_MAPQ=19;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=24;MATEID=5493823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_50249501_50274501_69C;SPAN=30044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:62 GQ:6.5 PL:[141.8, 0.0, 6.5] SR:33 DR:29 LR:-148.6 LO:148.6);ALT=C[chr13:50265389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50237332	+	chr13	50265389	+	.	0	21	5493824_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5493824_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_50249501_50274501_344C;SPAN=28057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:62 GQ:52.7 PL:[52.7, 0.0, 95.6] SR:21 DR:0 LR:-52.52 LO:53.28);ALT=C[chr13:50265389[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	64294924	+	chr13	50265389	+	.	0	47	6230913_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=55;MATEID=6230913_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_64288001_64313001_250C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:24 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:47 DR:0 LR:-138.6 LO:138.6);ALT=]chr16:64294924]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	64295143	+	chr13	50265515	+	.	26	0	6230914_1	75.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6230914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:50265515(-)-16:64295143(+)__16_64288001_64313001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:37 GQ:13.1 PL:[75.8, 0.0, 13.1] SR:0 DR:26 LR:-78.22 LO:78.22);ALT=]chr16:64295143]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr13	50571290	+	chr13	50586068	+	.	14	0	5494745_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5494745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:50571290(+)-13:50586068(-)__13_50568001_50593001D;SPAN=14778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:99 GQ:19.4 PL:[19.4, 0.0, 220.7] SR:0 DR:14 LR:-19.39 LO:29.4);ALT=C[chr13:50586068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	50571900	+	chr13	50586069	+	.	0	9	5494749_1	3.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5494749_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_50568001_50593001_269C;SPAN=14169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:96 GQ:3.8 PL:[3.8, 0.0, 228.2] SR:9 DR:0 LR:-3.7 LO:17.19);ALT=G[chr13:50586069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51069350	+	chr13	51075079	+	.	103	63	5496294_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCTC;MAPQ=60;MATEID=5496294_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_51058001_51083001_85C;SPAN=5729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:136 DP:33 GQ:36.6 PL:[402.6, 36.6, 0.0] SR:63 DR:103 LR:-402.7 LO:402.7);ALT=C[chr13:51075079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51484276	+	chr13	51501537	+	.	0	11	5497397_1	28.0	.	EVDNC=ASSMB;HOMSEQ=TTTCAG;MAPQ=60;MATEID=5497397_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_51474501_51499501_226C;SPAN=17261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:29 GQ:28.4 PL:[28.4, 0.0, 41.6] SR:11 DR:0 LR:-28.45 LO:28.6);ALT=G[chr13:51501537[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51484620	+	chr13	51503593	+	.	35	0	5497401_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5497401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:51484620(+)-13:51503593(-)__13_51474501_51499501D;SPAN=18973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:35 LR:-115.2 LO:115.2);ALT=T[chr13:51503593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51484917	+	chr13	51501536	+	.	20	0	5497403_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5497403_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:51484917(+)-13:51501536(-)__13_51474501_51499501D;SPAN=16619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:44 GQ:50.9 PL:[54.2, 0.0, 50.9] SR:0 DR:20 LR:-54.1 LO:54.1);ALT=G[chr13:51501536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51501615	+	chr13	51503608	+	.	3	34	5497249_1	91.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5497249_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_51499001_51524001_176C;SPAN=1993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:103 GQ:91.1 PL:[91.1, 0.0, 157.1] SR:34 DR:3 LR:-90.93 LO:91.95);ALT=G[chr13:51503608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51503719	+	chr13	51509019	+	AGGTCTTCTCCATTTTGCCACACCTGTGGATCCTCTATTTCTGCTTCTCCACTACCTCATAAAGGCTGATAAGG	2	32	5497255_1	76.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AGGTCTTCTCCATTTTGCCACACCTGTGGATCCTCTATTTCTGCTTCTCCACTACCTCATAAAGGCTGATAAGG;MAPQ=60;MATEID=5497255_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_51499001_51524001_325C;SPAN=5300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:107 GQ:76.7 PL:[76.7, 0.0, 182.3] SR:32 DR:2 LR:-76.64 LO:79.05);ALT=G[chr13:51509019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51504896	+	chr13	51509019	+	.	2	12	5497261_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=5497261_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGAGGA;SCTG=c_13_51499001_51524001_325C;SPAN=4123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:115 GQ:5.5 PL:[5.5, 0.0, 200.5] SR:12 DR:2 LR:-5.272 LO:18.7);ALT=G[chr13:51509019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	51528121	+	chr13	51530492	+	.	2	24	5497329_1	63.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5497329_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=AAAA;SCTG=c_13_51523501_51548501_53C;SPAN=2371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:83 GQ:63.5 PL:[63.5, 0.0, 136.1] SR:24 DR:2 LR:-63.34 LO:64.87);ALT=G[chr13:51530492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	52330598	+	chr13	52332328	+	.	2	3	5499690_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5499690_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_52307501_52332501_339C;SPAN=1730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:78 GQ:4.5 PL:[0.0, 4.5, 198.0] SR:3 DR:2 LR:4.627 LO:8.689);ALT=A[chr13:52332328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	52373843	+	chr13	52378188	+	.	9	0	5499382_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5499382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:52373843(+)-13:52378188(-)__13_52356501_52381501D;SPAN=4345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:0 DR:9 LR:-8.306 LO:17.99);ALT=G[chr13:52378188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53009019	+	chr13	53010425	+	.	0	16	5501582_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5501582_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_52993501_53018501_142C;SPAN=1406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:92 GQ:28.1 PL:[28.1, 0.0, 193.1] SR:16 DR:0 LR:-27.89 LO:35.18);ALT=T[chr13:53010425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53010541	+	chr13	53024634	+	CTTCCCAATTCCAGCCGCCTGTTCTTCAATGAACACAATTTGGGAAAGGAGAATGGCCATGCAACACTCATGATTTTTCTGATCTCTCCAAATCAGTCGGTGTGTACTAAGAAGGAGAGTCCCAGCATCAAATTTTAT	9	54	5502177_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTTCCCAATTCCAGCCGCCTGTTCTTCAATGAACACAATTTGGGAAAGGAGAATGGCCATGCAACACTCATGATTTTTCTGATCTCTCCAAATCAGTCGGTGTGTACTAAGAAGGAGAGTCCCAGCATCAAATTTTAT;MAPQ=60;MATEID=5502177_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_53018001_53043001_22C;SPAN=14093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:37 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:54 DR:9 LR:-178.2 LO:178.2);ALT=T[chr13:53024634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53013348	+	chr13	53024681	+	.	22	0	5502179_1	60.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5502179_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:53013348(+)-13:53024681(-)__13_53018001_53043001D;SPAN=11333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:44 GQ:44.3 PL:[60.8, 0.0, 44.3] SR:0 DR:22 LR:-60.81 LO:60.81);ALT=C[chr13:53024681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53016582	+	chr13	53024634	+	.	19	14	5502180_1	57.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5502180_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CTCCTC;SCTG=c_13_53018001_53043001_22C;SPAN=8052;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:37 GQ:8.3 PL:[57.7, 0.0, 8.3] SR:14 DR:19 LR:-60.03 LO:60.03);ALT=T[chr13:53024634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53191818	+	chr13	53196121	+	.	0	15	5502022_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=5502022_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_53189501_53214501_347C;SPAN=4303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:106 GQ:20.9 PL:[20.9, 0.0, 235.4] SR:15 DR:0 LR:-20.8 LO:31.5);ALT=G[chr13:53196121[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53227095	+	chr13	53232533	+	TTTTCCAGAGCTTCTCGGATGCCCTAATCGACGAGGACCCCCAGGCGGCGTTAGAGGAGCTGACTAAGGCTTTGGAACAGAAACCAGATGATGCACAGTATTATTGTCAAAGAGCTTATTGTCACATTCTTCTTGGGAATTACTGT	10	43	5502535_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TTTTCCAGAGCTTCTCGGATGCCCTAATCGACGAGGACCCCCAGGCGGCGTTAGAGGAGCTGACTAAGGCTTTGGAACAGAAACCAGATGATGCACAGTATTATTGTCAAAGAGCTTATTGTCACATTCTTCTTGGGAATTACTGT;MAPQ=60;MATEID=5502535_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_53214001_53239001_87C;SPAN=5438;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:94 GQ:96.8 PL:[129.8, 0.0, 96.8] SR:43 DR:10 LR:-129.9 LO:129.9);ALT=T[chr13:53232533[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	53227132	+	chr13	53231664	+	.	14	0	5502536_1	23.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5502536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:53227132(+)-13:53231664(-)__13_53214001_53239001D;SPAN=4532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:85 GQ:23.3 PL:[23.3, 0.0, 181.7] SR:0 DR:14 LR:-23.19 LO:30.41);ALT=C[chr13:53231664[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	74357263	+	chr13	74360260	+	.	0	36	5553853_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GGG;MAPQ=60;MATEID=5553853_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_74333001_74358001_361C;SPAN=2997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:32 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:36 DR:0 LR:-105.6 LO:105.6);ALT=G[chr13:74360260[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	82865266	-	chr13	82866400	+	GTTCTGTCCTGCCTTCTAGCTGTGCCTTCCAATTAGGCCCAAGTTCTCAAGCACATAAAACAAGACGAGAAGGAAACTTG	2	45	5575140_1	54.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ATTTTGGGG;INSERTION=GTTCTGTCCTGCCTTCTAGCTGTGCCTTCCAATTAGGCCCAAGTTCTCAAGCACATAAAACAAGACGAGAAGGAAACTTG;MAPQ=60;MATEID=5575140_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_13_82859001_82884001_38C;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:359 GQ:54.6 PL:[54.6, 0.0, 817.1] SR:45 DR:2 LR:-54.58 LO:94.47);ALT=[chr13:82866400[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	90328232	+	chr13	105798341	+	.	12	28	6027192_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6027192_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_90307001_90332001_201C;SPAN=-1;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:66 GQ:74.6 PL:[84.5, 0.0, 74.6] SR:28 DR:12 LR:-84.47 LO:84.47);ALT=]chr15:90328232]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr13	113223575	+	chr13	113242219	+	.	0	7	5652352_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5652352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_113239001_113264001_166C;SPAN=18644;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:34 GQ:14 PL:[14.0, 0.0, 66.8] SR:7 DR:0 LR:-13.9 LO:15.96);ALT=T[chr13:113242219[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113766676	+	chr13	113765507	+	.	14	0	5653783_1	18.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5653783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:113765507(-)-13:113766676(+)__13_113753501_113778501D;SPAN=1169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:103 GQ:18.5 PL:[18.5, 0.0, 229.7] SR:0 DR:14 LR:-18.31 LO:29.14);ALT=]chr13:113766676]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	113767490	+	chr13	113766059	+	.	13	0	5653784_1	23.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=5653784_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:113766059(-)-13:113767490(+)__13_113753501_113778501D;SPAN=1431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:74 GQ:23 PL:[23.0, 0.0, 155.0] SR:0 DR:13 LR:-22.86 LO:28.64);ALT=]chr13:113767490]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr13	113852626	+	chr13	113862909	+	.	8	0	5654134_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5654134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:113852626(+)-13:113862909(-)__13_113851501_113876501D;SPAN=10283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=A[chr13:113862909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113864403	+	chr13	113873256	+	.	0	10	5654161_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=5654161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_113851501_113876501_83C;SPAN=8853;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:10 DR:0 LR:-12.96 LO:20.79);ALT=G[chr13:113873256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113951810	+	chr13	113963957	+	.	4	3	5654457_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5654457_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_113949501_113974501_232C;SPAN=12147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:3 DR:4 LR:-3.059 LO:13.4);ALT=G[chr13:113963957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113951811	+	chr13	113960799	+	.	0	23	5654458_1	53.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5654458_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_113949501_113974501_43C;SPAN=8988;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:83 GQ:53.6 PL:[53.6, 0.0, 146.0] SR:23 DR:0 LR:-53.44 LO:55.9);ALT=G[chr13:113960799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	113965175	+	chr13	113973782	+	AGGGG	2	4	5654514_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AGGGG;MAPQ=60;MATEID=5654514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_113949501_113974501_116C;SPAN=8607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:97 GQ:9.6 PL:[0.0, 9.6, 254.1] SR:4 DR:2 LR:9.775 LO:8.204);ALT=C[chr13:113973782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114000398	+	chr13	114001703	+	.	16	0	5654874_1	42.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5654874_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:114000398(+)-13:114001703(-)__13_113998501_114023501D;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:38 GQ:42.5 PL:[42.5, 0.0, 49.1] SR:0 DR:16 LR:-42.52 LO:42.55);ALT=C[chr13:114001703[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114050170	+	chr13	114054604	+	.	15	0	5654991_1	35.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5654991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:114050170(+)-13:114054604(-)__13_114047501_114072501D;SPAN=4434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:0 DR:15 LR:-34.89 LO:36.48);ALT=G[chr13:114054604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114145588	+	chr13	114149816	+	.	24	23	5655136_1	96.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5655136_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_114145501_114170501_311C;SPAN=4228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:83 GQ:96.5 PL:[96.5, 0.0, 103.1] SR:23 DR:24 LR:-96.35 LO:96.37);ALT=G[chr13:114149816[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114150341	+	chr13	114152655	+	.	3	5	5655147_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5655147_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_114145501_114170501_47C;SPAN=2314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:100 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:5 DR:3 LR:0.6845 LO:14.7);ALT=G[chr13:114152655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	114239203	+	chr15	79852904	-	.	6	3	5998754_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGGCTGCCCGGTCCGGCCGCGCGGGCGGGG;MAPQ=60;MATEID=5998754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_79845501_79870501_149C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:3 DR:6 LR:-23.75 LO:23.78);ALT=G]chr15:79852904];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr13	114505560	+	chr13	114506636	+	.	26	20	5656155_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GACCC;MAPQ=60;MATEID=5656155_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_114488501_114513501_348C;SPAN=1076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:48 GQ:0.2 PL:[115.7, 0.0, 0.2] SR:20 DR:26 LR:-122.7 LO:122.7);ALT=C[chr13:114506636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	115000607	+	chr13	115002273	+	CAACAGTATCAAAGTGCTCTATTTTGGGCAGATAAAGTAGCTTCACTCTCTCGT	0	9	5657188_1	5.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CAACAGTATCAAAGTGCTCTATTTTGGGCAGATAAAGTAGCTTCACTCTCTCGT;MAPQ=60;MATEID=5657188_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_114978501_115003501_212C;SPAN=1666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:9 DR:0 LR:-5.326 LO:17.45);ALT=G[chr13:115002273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	115000607	+	chr13	115002117	+	.	6	6	5657187_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=5657187_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_13_114978501_115003501_212C;SPAN=1510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:6 DR:6 LR:-13.82 LO:22.76);ALT=G[chr13:115002117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	115097045	+	chr13	115098107	-	.	9	0	5657505_1	8.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5657505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:115097045(+)-13:115098107(+)__13_115076501_115101501D;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:0 DR:9 LR:-8.577 LO:18.05);ALT=T]chr13:115098107];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	29215127	-	chr17	64928552	+	.	2	17	5686089_1	56.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTAATTTAATTTAATTTAATTTAATTT;MAPQ=60;MATEID=5686089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_29204001_29229001_167C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:22 GQ:2.4 PL:[56.1, 2.4, 0.0] SR:17 DR:2 LR:-56.8 LO:56.8);ALT=[chr17:64928552[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	29493717	+	chr14	29492501	+	.	9	0	5686712_1	7.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=5686712_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:29492501(-)-14:29493717(+)__14_29473501_29498501D;SPAN=1216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=]chr14:29493717]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	31091618	+	chr14	31099680	+	.	10	0	5689917_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5689917_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:31091618(+)-14:31099680(-)__14_31090501_31115501D;SPAN=8062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:0 DR:10 LR:-11.34 LO:20.42);ALT=T[chr14:31099680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	31099772	+	chr14	31103153	+	.	0	12	5689940_1	19.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5689940_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_31090501_31115501_276C;SPAN=3381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:12 DR:0 LR:-19.29 LO:25.9);ALT=G[chr14:31103153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	31675163	+	chr14	31676597	+	.	10	5	5691558_1	15.0	.	DISC_MAPQ=56;EVDNC=TSI_L;MAPQ=60;MATEID=5691558_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_31654001_31679001_46C;SPAN=1434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:5 DR:10 LR:-15.45 LO:23.15);ALT=G[chr14:31676597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	31789766	-	chr17	46972515	+	.	75	0	6420812_1	99.0	.	DISC_MAPQ=5;EVDNC=DSCRD;IMPRECISE;MAPQ=5;MATEID=6420812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:31789766(-)-17:46972515(-)__17_46966501_46991501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:55 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:0 DR:75 LR:-221.2 LO:221.2);ALT=[chr17:46972515[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr14	31982787	+	chr20	35270568	+	.	27	0	5692326_1	78.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=5692326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:31982787(+)-20:35270568(-)__14_31972501_31997501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:39 GQ:15.8 PL:[78.5, 0.0, 15.8] SR:0 DR:27 LR:-80.89 LO:80.89);ALT=A[chr20:35270568[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr14	32279042	+	chr14	32087674	+	.	8	0	5693498_1	19.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=5693498_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:32087674(-)-14:32279042(+)__14_32266501_32291501D;SPAN=191368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:27 GQ:19.1 PL:[19.1, 0.0, 45.5] SR:0 DR:8 LR:-19.09 LO:19.72);ALT=]chr14:32279042]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	32953311	+	chr14	32954349	+	.	39	0	5695354_1	99.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=5695354_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:32953311(+)-14:32954349(-)__14_32952501_32977501D;SPAN=1038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:5 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:39 LR:-115.5 LO:115.5);ALT=T[chr14:32954349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	34904510	+	chr14	34931302	+	.	0	11	5699409_1	28.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5699409_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_34912501_34937501_124C;SPAN=26792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:30 GQ:28.1 PL:[28.1, 0.0, 44.6] SR:11 DR:0 LR:-28.18 LO:28.39);ALT=T[chr14:34931302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35002746	+	chr14	35005299	+	.	0	11	5699559_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5699559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_34986001_35011001_352C;SPAN=2553;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:86 GQ:13.1 PL:[13.1, 0.0, 194.6] SR:11 DR:0 LR:-13.01 LO:22.58);ALT=C[chr14:35005299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35005483	+	chr14	35008761	+	.	25	15	5699571_1	81.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5699571_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_34986001_35011001_16C;SPAN=3278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:88 GQ:81.8 PL:[81.8, 0.0, 131.3] SR:15 DR:25 LR:-81.79 LO:82.43);ALT=T[chr14:35008761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35038226	+	chr19	42364392	-	.	17	0	5700297_1	25.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=5700297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35038226(+)-19:42364392(+)__14_35035001_35060001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:113 GQ:25.7 PL:[25.7, 0.0, 246.8] SR:0 DR:17 LR:-25.5 LO:36.2);ALT=A]chr19:42364392];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr14	35048572	-	chr14	35049657	+	.	13	0	5700341_1	24.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5700341_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35048572(-)-14:35049657(-)__14_35035001_35060001D;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:69 GQ:24.2 PL:[24.2, 0.0, 143.0] SR:0 DR:13 LR:-24.22 LO:29.08);ALT=[chr14:35049657[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	35077348	+	chr14	35078844	+	.	0	26	5700228_1	61.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=56;MATEID=5700228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_35059501_35084501_48C;SPAN=1496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:89 GQ:61.7 PL:[61.7, 0.0, 154.1] SR:26 DR:0 LR:-61.71 LO:63.91);ALT=T[chr14:35078844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35077388	+	chr14	35099112	+	.	19	0	5700229_1	51.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5700229_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35077388(+)-14:35099112(-)__14_35059501_35084501D;SPAN=21724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:41 GQ:45.2 PL:[51.8, 0.0, 45.2] SR:0 DR:19 LR:-51.62 LO:51.62);ALT=A[chr14:35099112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35077392	+	chr14	35099314	+	.	15	0	5700230_1	38.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=5700230_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35077392(+)-14:35099314(-)__14_35059501_35084501D;SPAN=21922;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:41 GQ:38.6 PL:[38.6, 0.0, 58.4] SR:0 DR:15 LR:-38.41 LO:38.69);ALT=A[chr14:35099314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35078948	+	chr14	35099113	+	.	4	6	5700235_1	20.0	.	DISC_MAPQ=32;EVDNC=ASDIS;MAPQ=60;MATEID=5700235_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_35059501_35084501_212C;SPAN=20165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:33 GQ:20.9 PL:[20.9, 0.0, 57.2] SR:6 DR:4 LR:-20.77 LO:21.8);ALT=G[chr14:35099113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35078998	+	chr14	35099315	+	.	11	0	5700236_1	29.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=5700236_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35078998(+)-14:35099315(-)__14_35059501_35084501D;SPAN=20317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:26 GQ:29.3 PL:[29.3, 0.0, 32.6] SR:0 DR:11 LR:-29.27 LO:29.29);ALT=T[chr14:35099315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35253136	+	chr14	35254982	+	.	0	12	5701180_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=5701180_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_35231001_35256001_57C;SPAN=1846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:12 DR:0 LR:-18.21 LO:25.61);ALT=G[chr14:35254982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35264127	+	chr14	35269428	+	.	11	0	5700645_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5700645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35264127(+)-14:35269428(-)__14_35255501_35280501D;SPAN=5301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:71 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:0 DR:11 LR:-17.08 LO:23.58);ALT=A[chr14:35269428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35452421	+	chr14	35465882	+	.	6	13	5701562_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5701562_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_35451501_35476501_78C;SPAN=13461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:95 GQ:23.9 PL:[23.9, 0.0, 205.4] SR:13 DR:6 LR:-23.78 LO:32.28);ALT=G[chr14:35465882[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35579187	+	chr14	35591115	+	.	11	0	5701986_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5701986_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35579187(+)-14:35591115(-)__14_35574001_35599001D;SPAN=11928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:0 DR:11 LR:-15.99 LO:23.29);ALT=T[chr14:35591115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35579836	+	chr14	35585816	+	.	3	10	5701987_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5701987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_35574001_35599001_136C;SPAN=5980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:78 GQ:18.5 PL:[18.5, 0.0, 170.3] SR:10 DR:3 LR:-18.48 LO:25.68);ALT=C[chr14:35585816[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35579851	+	chr14	35591107	+	.	14	0	5701988_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5701988_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35579851(+)-14:35591107(-)__14_35574001_35599001D;SPAN=11256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:74 GQ:26.3 PL:[26.3, 0.0, 151.7] SR:0 DR:14 LR:-26.17 LO:31.35);ALT=A[chr14:35591107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35592116	+	chr14	35596683	+	TGTTCCTGGAAAACAATGGAAAGGACAATTCACCACAGTCCGAAAA	0	11	5702025_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGTTCCTGGAAAACAATGGAAAGGACAATTCACCACAGTCCGAAAA;MAPQ=60;MATEID=5702025_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_35574001_35599001_185C;SPAN=4567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:11 DR:0 LR:-17.89 LO:23.8);ALT=C[chr14:35596683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	35761736	+	chr14	35777196	+	.	33	0	5702629_1	96.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=5702629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:35761736(+)-14:35777196(-)__14_35770001_35795001D;SPAN=15460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:47 GQ:17 PL:[96.2, 0.0, 17.0] SR:0 DR:33 LR:-99.25 LO:99.25);ALT=C[chr14:35777196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	36133973	+	chr14	36140594	+	.	0	20	5703660_1	56.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=49;MATEID=5703660_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_36113001_36138001_236C;SPAN=6621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:34 GQ:23.9 PL:[56.9, 0.0, 23.9] SR:20 DR:0 LR:-57.44 LO:57.44);ALT=C[chr14:36140594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67880921	+	chr14	36289080	+	.	28	0	6236824_1	82.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=6236824_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:36289080(-)-16:67880921(+)__16_67865001_67890001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:18 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:0 DR:28 LR:-82.52 LO:82.52);ALT=]chr16:67880921]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr14	36418509	+	chr14	36417419	+	.	11	0	5704359_1	14.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=5704359_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:36417419(-)-14:36418509(+)__14_36407001_36432001D;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:80 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:0 DR:11 LR:-14.64 LO:22.95);ALT=]chr14:36418509]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	44248335	+	chr14	43824277	+	.	64	66	5722667_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAT;MAPQ=60;MATEID=5722667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_44247001_44272001_22C;SPAN=424058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:50 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:66 DR:64 LR:-303.7 LO:303.7);ALT=]chr14:44248335]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	45591219	+	chr14	44835568	+	.	7	14	5724161_1	51.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=TTTTTTTTTTTTTTTTTTT;MAPQ=27;MATEID=5724161_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_44835001_44860001_214C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:42 GQ:48.2 PL:[51.5, 0.0, 48.2] SR:14 DR:7 LR:-51.34 LO:51.34);ALT=]chr19:45591219]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr14	45415133	+	chr14	45431049	+	.	18	3	5725416_1	54.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5725416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_45423001_45448001_246C;SPAN=15916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:32 GQ:21.2 PL:[54.2, 0.0, 21.2] SR:3 DR:18 LR:-54.7 LO:54.7);ALT=T[chr14:45431049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45585455	+	chr14	45587231	+	.	2	11	5725847_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=5725847_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_14_45570001_45595001_229C;SPAN=1776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:11 DR:2 LR:-21.19 LO:26.47);ALT=T[chr14:45587231[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45585455	+	chr14	45590090	+	TTGGCATCAGGCTGTCCTTTCTTTCCGTAAGCCCATTCTGGTTCAATCTCCAGTCGAGCCTTTTCTCCTTTACTCATAGTCAAGAGAGCTTCATCCCA	8	16	5725848_1	52.0	.	DISC_MAPQ=60;EVDNC=TSI_G;INSERTION=TTGGCATCAGGCTGTCCTTTCTTTCCGTAAGCCCATTCTGGTTCAATCTCCAGTCGAGCCTTTTCTCCTTTACTCATAGTCAAGAGAGCTTCATCCCA;MAPQ=60;MATEID=5725848_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_45570001_45595001_229C;SPAN=4635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:75 GQ:52.4 PL:[52.4, 0.0, 128.3] SR:16 DR:8 LR:-52.3 LO:54.12);ALT=T[chr14:45590090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45587370	+	chr14	45590685	+	.	8	0	5725856_1	7.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5725856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:45587370(+)-14:45590685(-)__14_45570001_45595001D;SPAN=3315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.172 LO:15.95);ALT=A[chr14:45590685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45590825	+	chr14	45599902	+	CATCCAGGGTCTCTTCAGACTTGGTTTCTTTGGGTTTATCTTCATTAAGCTTCACATTTTTTACTTGCTCAGACACTTTACTTATACTTTCAGTACCCTTAAAACG	3	46	5726013_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CATCCAGGGTCTCTTCAGACTTGGTTTCTTTGGGTTTATCTTCATTAAGCTTCACATTTTTTACTTGCTCAGACACTTTACTTATACTTTCAGTACCCTTAAAACG;MAPQ=60;MATEID=5726013_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_45594501_45619501_9C;SPAN=9077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:45 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:46 DR:3 LR:-138.6 LO:138.6);ALT=T[chr14:45599902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45599149	+	chr14	45603575	+	.	15	0	5726028_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5726028_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:45599149(+)-14:45603575(-)__14_45594501_45619501D;SPAN=4426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:87 GQ:26 PL:[26.0, 0.0, 184.4] SR:0 DR:15 LR:-25.94 LO:32.91);ALT=C[chr14:45603575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45600004	+	chr14	45603552	+	.	0	12	5726032_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5726032_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_45594501_45619501_281C;SPAN=3548;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:94 GQ:14.3 PL:[14.3, 0.0, 212.3] SR:12 DR:0 LR:-14.15 LO:24.62);ALT=C[chr14:45603552[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	45716582	+	chr14	45722236	+	.	38	10	5726228_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5726228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_45717001_45742001_332C;SPAN=5654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:10 DR:38 LR:-141.4 LO:141.4);ALT=T[chr14:45722236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	47117868	-	chr14	63226284	+	.	40	32	5729177_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=A;MAPQ=0;MATEID=5729177_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GGG;SCTG=c_14_47113501_47138501_134C;SECONDARY;SPAN=16108416;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:51 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:32 DR:40 LR:-191.4 LO:191.4);ALT=[chr14:63226284[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	49331368	+	chr14	49333935	+	.	92	82	5733830_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=GCT;MAPQ=60;MATEID=5733830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_49318501_49343501_217C;SPAN=2567;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:40 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:82 DR:92 LR:-415.9 LO:415.9);ALT=T[chr14:49333935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	50312985	+	chr14	50318281	+	.	0	9	5736191_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5736191_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_50298501_50323501_212C;SPAN=5296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:70 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:9 DR:0 LR:-10.74 LO:18.5);ALT=T[chr14:50318281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	50318383	+	chr14	50319413	+	TTTTGAAGACGAATAAGGTATGTCTTATTATCCACATCATAAACATTGTTTACTCTCATTCCTAGCAAG	0	21	5736212_1	44.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTTTGAAGACGAATAAGGTATGTCTTATTATCCACATCATAAACATTGTTTACTCTCATTCCTAGCAAG;MAPQ=60;MATEID=5736212_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_50298501_50323501_13C;SPAN=1030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:92 GQ:44.6 PL:[44.6, 0.0, 176.6] SR:21 DR:0 LR:-44.4 LO:48.97);ALT=T[chr14:50319413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	50779139	+	chr14	50789228	+	.	9	0	5737908_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5737908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:50779139(+)-14:50789228(-)__14_50788501_50813501D;SPAN=10089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=G[chr14:50789228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	50789437	+	chr14	50790662	+	.	0	4	5737912_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5737912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_50788501_50813501_149C;SPAN=1225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:89 GQ:10.8 PL:[0.0, 10.8, 237.6] SR:4 DR:0 LR:10.91 LO:6.32);ALT=G[chr14:50790662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	50790834	+	chr14	50792325	+	.	5	6	5737916_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5737916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_50788501_50813501_230C;SPAN=1491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:6 DR:5 LR:-9.932 LO:18.32);ALT=G[chr14:50792325[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	51288844	+	chr14	51297793	+	.	13	0	5739285_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5739285_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:51288844(+)-14:51297793(-)__14_51278501_51303501D;SPAN=8949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:66 GQ:25.1 PL:[25.1, 0.0, 134.0] SR:0 DR:13 LR:-25.03 LO:29.37);ALT=C[chr14:51297793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	51404557	+	chr14	51410879	+	.	0	14	5739832_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5739832_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_51401001_51426001_95C;SPAN=6322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:82 GQ:24.2 PL:[24.2, 0.0, 172.7] SR:14 DR:0 LR:-24.0 LO:30.65);ALT=T[chr14:51410879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	51658535	+	chrX	19710867	-	.	9	0	5740337_1	23.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5740337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:51658535(+)-23:19710867(+)__14_51646001_51671001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=A]chrX:19710867];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr14	51707162	+	chr14	51710574	+	.	0	19	5740622_1	35.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5740622_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_51695001_51720001_332C;SPAN=3412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:99 GQ:35.9 PL:[35.9, 0.0, 204.2] SR:19 DR:0 LR:-35.9 LO:42.68);ALT=T[chr14:51710574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	52456418	+	chr14	52460439	+	ATGAAACAGAATTTAGAAACTTCATCGTTTGGCTTGAAGACCAGAAAATCAGGCACTACAAGATTGAAGACAGAGGGAATTTAAGAAACATCCACAGCAGCGACTGGCCCAAGTTCTTTGAAA	12	183	5742363_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=AGTATCTCAGAGATGTTAACTGTCCTTTCAAGATTCAAGATCGACAAGAAGCTATTGACTGGCTTCTTGGTTTAGCTGTTAGACTTGAATATGGAGAT;INSERTION=ATGAAACAGAATTTAGAAACTTCATCGTTTGGCTTGAAGACCAGAAAATCAGGCACTACAAGATTGAAGACAGAGGGAATTTAAGAAACATCCACAGCAGCGACTGGCCCAAGTTCTTTGAAA;MAPQ=60;MATEID=5742363_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_52454501_52479501_323C;SECONDARY;SPAN=4021;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:188 DP:105 GQ:50.8 PL:[557.8, 50.8, 0.0] SR:183 DR:12 LR:-557.8 LO:557.8);ALT=G[chr14:52460439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	52456418	+	chr14	52458033	+	.	71	75	5742362_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5742362_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_52454501_52479501_323C;SPAN=1615;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:104 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:75 DR:71 LR:-389.5 LO:389.5);ALT=G[chr14:52458033[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	53251383	+	chr14	53258146	+	.	5	2	5744517_1	0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5744517_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_53238501_53263501_50C;SPAN=6763;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:72 GQ:0.5 PL:[0.5, 0.0, 172.1] SR:2 DR:5 LR:-0.2994 LO:11.14);ALT=C[chr14:53258146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54655743	+	chrX	121656448	-	.	7	1	5747929_1	9.0	.	DISC_MAPQ=46;EVDNC=TSI_L;HOMSEQ=ACACACACACACACAC;MAPQ=60;MATEID=5747929_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TGTGTGTGTGTGTGTGTGTGTGTGTGTG;SCTG=c_14_54635001_54660001_318C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:8 DP:11 GQ:1.1 PL:[9.6, 1.1, 0.0] SR:1 DR:7 LR:-8.973 LO:8.973);ALT=T]chrX:121656448];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr14	54710349	+	chr14	54713686	+	.	90	61	5748017_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TGA;MAPQ=60;MATEID=5748017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54708501_54733501_165C;SPAN=3337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:123 DP:33 GQ:33 PL:[363.0, 33.0, 0.0] SR:61 DR:90 LR:-363.1 LO:363.1);ALT=A[chr14:54713686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54894560	+	chr14	54896979	+	.	0	9	5748398_1	7.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5748398_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54880001_54905001_220C;SPAN=2419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:9 DR:0 LR:-7.222 LO:17.79);ALT=C[chr14:54896979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54897122	+	chr14	54903084	+	.	0	9	5748405_1	5.0	.	EVDNC=ASSMB;HOMSEQ=TAC;MAPQ=60;MATEID=5748405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54880001_54905001_183C;SPAN=5962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:9 DR:0 LR:-5.868 LO:17.54);ALT=C[chr14:54903084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54897124	+	chr14	54898823	+	.	0	34	5748406_1	87.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=5748406_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54880001_54905001_300C;SPAN=1699;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:92 GQ:87.5 PL:[87.5, 0.0, 133.7] SR:34 DR:0 LR:-87.31 LO:87.89);ALT=T[chr14:54898823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54897171	+	chr14	54907992	+	.	33	0	5748494_1	95.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5748494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54897171(+)-14:54907992(-)__14_54904501_54929501D;SPAN=10821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:48 GQ:20 PL:[95.9, 0.0, 20.0] SR:0 DR:33 LR:-98.67 LO:98.67);ALT=C[chr14:54907992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54898938	+	chr14	54903087	+	.	0	63	5748411_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5748411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54880001_54905001_110C;SPAN=4149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:96 GQ:50 PL:[182.0, 0.0, 50.0] SR:63 DR:0 LR:-186.0 LO:186.0);ALT=G[chr14:54903087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54898987	+	chr14	54907989	+	.	66	0	5748495_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5748495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54898987(+)-14:54907989(-)__14_54904501_54929501D;SPAN=9002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:42 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:0 DR:66 LR:-194.7 LO:194.7);ALT=A[chr14:54907989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54903155	+	chr14	54907965	+	.	36	23	5748496_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5748496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54904501_54929501_119C;SPAN=4810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:28 GQ:12 PL:[132.0, 12.0, 0.0] SR:23 DR:36 LR:-132.0 LO:132.0);ALT=T[chr14:54907965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54950483	+	chr14	54955636	+	.	26	0	5748629_1	72.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5748629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54950483(+)-14:54955636(-)__14_54953501_54978501D;SPAN=5153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:48 GQ:43.1 PL:[72.8, 0.0, 43.1] SR:0 DR:26 LR:-73.21 LO:73.21);ALT=A[chr14:54955636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54976743	+	chr14	54989170	+	.	10	0	5748690_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5748690_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:54976743(+)-14:54989170(-)__14_54953501_54978501D;SPAN=12427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=T[chr14:54989170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	54989311	+	chr14	54996767	+	.	0	9	5748588_1	10.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5748588_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_54978001_55003001_222C;SPAN=7456;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:9 DR:0 LR:-9.932 LO:18.32);ALT=A[chr14:54996767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55518513	+	chr14	55524733	+	.	9	0	5750203_1	4.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5750203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55518513(+)-14:55524733(-)__14_55517001_55542001D;SPAN=6220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:93 GQ:4.7 PL:[4.7, 0.0, 219.2] SR:0 DR:9 LR:-4.513 LO:17.32);ALT=T[chr14:55524733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55518521	+	chr14	55529335	+	.	22	2	5750204_1	50.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5750204_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_14_55517001_55542001_53C;SECONDARY;SPAN=10814;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:96 GQ:50 PL:[50.0, 0.0, 182.0] SR:2 DR:22 LR:-49.91 LO:54.19);ALT=G[chr14:55529335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55596062	+	chr14	55604760	+	.	51	0	5750397_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5750397_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:55596062(+)-14:55604760(-)__14_55590501_55615501D;SPAN=8698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:74 GQ:29.6 PL:[148.4, 0.0, 29.6] SR:0 DR:51 LR:-152.6 LO:152.6);ALT=G[chr14:55604760[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	55609467	+	chr14	55611834	+	.	5	10	5750446_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5750446_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_55590501_55615501_339C;SPAN=2367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:80 GQ:27.8 PL:[27.8, 0.0, 166.4] SR:10 DR:5 LR:-27.84 LO:33.52);ALT=A[chr14:55611834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56047074	+	chr14	56078736	+	.	40	16	5752052_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5752052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56056001_56081001_199C;SPAN=31662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:39 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:16 DR:40 LR:-148.5 LO:148.5);ALT=T[chr14:56078736[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56047074	+	chr14	56068474	+	.	10	8	5752051_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5752051_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56056001_56081001_139C;SPAN=21400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:36 GQ:36.5 PL:[36.5, 0.0, 49.7] SR:8 DR:10 LR:-36.46 LO:36.59);ALT=T[chr14:56068474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56068600	+	chr14	56078735	+	.	0	15	5752091_1	26.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5752091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56056001_56081001_27C;SPAN=10135;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:15 DR:0 LR:-26.49 LO:33.08);ALT=T[chr14:56078735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56079289	+	chr14	56083234	+	.	3	4	5752127_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5752127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56080501_56105501_343C;SPAN=3945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:40 GQ:2.3 PL:[2.3, 0.0, 94.7] SR:4 DR:3 LR:-2.367 LO:7.756);ALT=G[chr14:56083234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56096815	+	chr14	56099951	+	.	2	3	5752161_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5752161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56080501_56105501_352C;SPAN=3136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:63 GQ:0.3 PL:[0.0, 0.3, 151.8] SR:3 DR:2 LR:0.5633 LO:9.169);ALT=G[chr14:56099951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56142637	+	chr14	56145068	+	.	2	4	5752463_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=5752463_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_14_56129501_56154501_94C;SPAN=2431;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:4 DR:2 LR:1.055 LO:10.95);ALT=G[chr14:56145068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	56146403	+	chr14	56150815	+	.	3	5	5752475_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5752475_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_56129501_56154501_206C;SPAN=4412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:81 GQ:1.4 PL:[1.4, 0.0, 192.8] SR:5 DR:3 LR:-1.162 LO:13.11);ALT=G[chr14:56150815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58666995	+	chr14	58674651	+	.	8	0	5758094_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5758094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58666995(+)-14:58674651(-)__14_58653001_58678001D;SPAN=7656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:64 GQ:9.2 PL:[9.2, 0.0, 144.5] SR:0 DR:8 LR:-9.069 LO:16.34);ALT=G[chr14:58674651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58667015	+	chr14	58669573	+	.	10	12	5758095_1	35.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GTG;MAPQ=60;MATEID=5758095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58653001_58678001_106C;SPAN=2558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:65 GQ:35.3 PL:[35.3, 0.0, 121.1] SR:12 DR:10 LR:-35.21 LO:37.92);ALT=G[chr14:58669573[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58669645	+	chr14	58674652	+	.	0	11	5758101_1	16.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5758101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58653001_58678001_199C;SPAN=5007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:11 DR:0 LR:-16.53 LO:23.43);ALT=G[chr14:58674652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58678121	+	chr14	58680349	+	.	0	7	5758641_1	0	.	EVDNC=ASSMB;HOMSEQ=ATAT;MAPQ=60;MATEID=5758641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58677501_58702501_359C;SPAN=2228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:84 GQ:0.5 PL:[0.5, 0.0, 201.8] SR:7 DR:0 LR:-0.3493 LO:12.99);ALT=T[chr14:58680349[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58711659	+	chr14	58718835	+	TATGACCTGTCAGCCTCTACATTCTCTCCTGACGGAAGAGTTTTTCAAGTTGAATATGCTATGAAGGCTGTGGAAAATAGT	41	22	5758570_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TATGACCTGTCAGCCTCTACATTCTCTCCTGACGGAAGAGTTTTTCAAGTTGAATATGCTATGAAGGCTGTGGAAAATAGT;MAPQ=60;MATEID=5758570_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_58702001_58727001_369C;SPAN=7176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:82 GQ:50.6 PL:[146.3, 0.0, 50.6] SR:22 DR:41 LR:-148.5 LO:148.5);ALT=G[chr14:58718835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58711659	+	chr14	58714467	+	.	9	4	5758569_1	13.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5758569_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_14_58702001_58727001_369C;SPAN=2808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:4 DR:9 LR:-13.55 LO:22.7);ALT=G[chr14:58714467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58711707	+	chr14	58724461	+	.	9	0	5758571_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5758571_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58711707(+)-14:58724461(-)__14_58702001_58727001D;SPAN=12754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:85 GQ:6.8 PL:[6.8, 0.0, 198.2] SR:0 DR:9 LR:-6.68 LO:17.69);ALT=T[chr14:58724461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58718961	+	chr14	58724462	+	.	0	24	5758581_1	59.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5758581_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58702001_58727001_149C;SPAN=5501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:74 GQ:59.3 PL:[59.3, 0.0, 118.7] SR:24 DR:0 LR:-59.18 LO:60.32);ALT=G[chr14:58724462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58730488	+	chr14	58737652	+	ATGAAAGAAATGACCTGCCGTGATATCGTTAAAGAAGTTGCAAAAATAATTTACATAGTACATGACGAAGTTAAGGATAAAGCTTTTGAACTAGAACTCAGCTGGGTTGGTGAAT	0	31	5758212_1	78.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATGAAAGAAATGACCTGCCGTGATATCGTTAAAGAAGTTGCAAAAATAATTTACATAGTACATGACGAAGTTAAGGATAAAGCTTTTGAACTAGAACTCAGCTGGGTTGGTGAAT;MAPQ=60;MATEID=5758212_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_14_58726501_58751501_43C;SPAN=7164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:87 GQ:78.8 PL:[78.8, 0.0, 131.6] SR:31 DR:0 LR:-78.76 LO:79.51);ALT=G[chr14:58737652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58734092	+	chr14	58740696	+	.	8	0	5758223_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5758223_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58734092(+)-14:58740696(-)__14_58726501_58751501D;SPAN=6604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:0 DR:8 LR:-6.089 LO:15.75);ALT=T[chr14:58740696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58758427	+	chr14	58764673	+	.	0	20	5758469_1	41.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5758469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58751001_58776001_80C;SPAN=6246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:90 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:20 DR:0 LR:-41.64 LO:46.37);ALT=T[chr14:58764673[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58762531	+	chr14	58764673	+	.	0	9	5758489_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5758489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58751001_58776001_237C;SPAN=2142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:9 DR:0 LR:-1.804 LO:16.9);ALT=T[chr14:58764673[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58877710	+	chr14	58893805	+	.	10	0	5759067_1	14.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5759067_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58877710(+)-14:58893805(-)__14_58873501_58898501D;SPAN=16095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:0 DR:10 LR:-14.59 LO:21.18);ALT=T[chr14:58893805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58878691	+	chr14	58890724	+	.	0	17	5759072_1	32.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=5759072_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_58873501_58898501_203C;SPAN=12033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:88 GQ:32.3 PL:[32.3, 0.0, 180.8] SR:17 DR:0 LR:-32.28 LO:38.24);ALT=T[chr14:58890724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58878731	+	chr14	58893825	+	.	13	0	5759073_1	20.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=5759073_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58878731(+)-14:58893825(-)__14_58873501_58898501D;SPAN=15094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:85 GQ:20 PL:[20.0, 0.0, 185.0] SR:0 DR:13 LR:-19.88 LO:27.78);ALT=A[chr14:58893825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	58890858	+	chr14	58893825	+	.	15	0	5759113_1	28.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5759113_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:58890858(+)-14:58893825(-)__14_58873501_58898501D;SPAN=2967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:79 GQ:28.1 PL:[28.1, 0.0, 163.4] SR:0 DR:15 LR:-28.11 LO:33.61);ALT=A[chr14:58893825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	59655534	+	chr14	59730155	+	.	8	0	5761118_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5761118_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:59655534(+)-14:59730155(-)__14_59706501_59731501D;SPAN=74621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:0 DR:8 LR:-8.527 LO:16.22);ALT=C[chr14:59730155[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	59951350	+	chr14	59953474	+	.	11	0	5761371_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5761371_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:59951350(+)-14:59953474(-)__14_59951501_59976501D;SPAN=2124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:0 DR:11 LR:-26.29 LO:27.14);ALT=G[chr14:59953474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	59953525	+	chr14	59961734	+	TGCCCAAGAGGACAGAGAACGAATGCACAGAAATATTGTCAGCCTTGCACAGAATCTCCTGAACTTTATGATTGGCTCTATCTTGGATTTATGGCAATGCTTCCTCTGGTTTTACATTGGTTCTTCATTGAATGGTACTCGGGGAAAAAG	0	17	5761373_1	34.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TGCCCAAGAGGACAGAGAACGAATGCACAGAAATATTGTCAGCCTTGCACAGAATCTCCTGAACTTTATGATTGGCTCTATCTTGGATTTATGGCAATGCTTCCTCTGGTTTTACATTGGTTCTTCATTGAATGGTACTCGGGGAAAAAG;MAPQ=60;MATEID=5761373_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_59951501_59976501_263C;SPAN=8209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:81 GQ:34.4 PL:[34.4, 0.0, 159.8] SR:17 DR:0 LR:-34.17 LO:38.93);ALT=A[chr14:59961734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	60611732	+	chr14	60616070	+	.	5	8	5762997_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5762997_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_60613001_60638001_266C;SPAN=4338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:8 DR:5 LR:-30.4 LO:30.71);ALT=C[chr14:60616070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	60622872	+	chr14	60631895	+	.	0	38	5763017_1	96.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5763017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_60613001_60638001_264C;SPAN=9023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:106 GQ:96.8 PL:[96.8, 0.0, 159.5] SR:38 DR:0 LR:-96.72 LO:97.59);ALT=T[chr14:60631895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	60913796	-	chr14	60941206	+	.	27	0	5763701_1	79.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=5763701_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:60913796(-)-14:60941206(-)__14_60931501_60956501D;SPAN=27410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:14 GQ:7.2 PL:[79.2, 7.2, 0.0] SR:0 DR:27 LR:-79.22 LO:79.22);ALT=[chr14:60941206[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	60914009	+	chr14	60941074	-	.	28	0	5763703_1	82.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=5763703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:60914009(+)-14:60941074(+)__14_60931501_60956501D;SPAN=27065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:17 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:0 DR:28 LR:-82.52 LO:82.52);ALT=T]chr14:60941074];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	61201669	+	chr14	61262935	+	.	0	7	5764582_1	14.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5764582_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_61250001_61275001_252C;SPAN=61266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:33 GQ:14.3 PL:[14.3, 0.0, 63.8] SR:7 DR:0 LR:-14.17 LO:16.07);ALT=T[chr14:61262935[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	62162558	+	chr14	62187100	+	.	0	13	5767024_1	30.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5767024_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_62181001_62206001_182C;SPAN=24542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:13 DR:0 LR:-30.18 LO:31.58);ALT=G[chr14:62187100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65360396	+	chr14	65363541	+	.	76	52	5775303_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AAGAATTTTC;MAPQ=60;MATEID=5775303_2;MATENM=4;NM=1;NUMPARTS=2;SCTG=c_14_65341501_65366501_300C;SPAN=3145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:33 GQ:27 PL:[297.0, 27.0, 0.0] SR:52 DR:76 LR:-297.1 LO:297.1);ALT=C[chr14:65363541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381253	+	chr14	65390708	+	.	87	8	5775401_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5775401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65390501_65415501_359C;SPAN=9455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:40 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:8 DR:87 LR:-267.4 LO:267.4);ALT=G[chr14:65390708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381279	+	chr14	65398853	+	.	36	0	5775402_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5775402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65381279(+)-14:65398853(-)__14_65390501_65415501D;SPAN=17574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:59 GQ:40.1 PL:[102.8, 0.0, 40.1] SR:0 DR:36 LR:-104.3 LO:104.3);ALT=C[chr14:65398853[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65381282	+	chr14	65392724	+	.	50	0	5775403_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5775403_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65381282(+)-14:65392724(-)__14_65390501_65415501D;SPAN=11442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:50 LR:-161.7 LO:161.7);ALT=G[chr14:65392724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65390844	+	chr14	65392728	+	.	0	83	5775407_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5775407_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65390501_65415501_253C;SPAN=1884;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:83 DP:121 GQ:50 PL:[241.4, 0.0, 50.0] SR:83 DR:0 LR:-248.0 LO:248.0);ALT=C[chr14:65392728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65390845	+	chr14	65398856	+	.	0	28	5775409_1	59.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5775409_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65390501_65415501_334C;SPAN=8011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:120 GQ:59.9 PL:[59.9, 0.0, 231.5] SR:28 DR:0 LR:-59.92 LO:65.6);ALT=G[chr14:65398856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65392799	+	chr14	65398854	+	.	0	82	5775413_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=5775413_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65390501_65415501_200C;SPAN=6055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:122 GQ:56.3 PL:[237.8, 0.0, 56.3] SR:82 DR:0 LR:-243.7 LO:243.7);ALT=G[chr14:65398854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65543383	+	chr14	65544631	+	.	5	7	5775606_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5775606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65537501_65562501_247C;SPAN=1248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:84 GQ:17 PL:[17.0, 0.0, 185.3] SR:7 DR:5 LR:-16.85 LO:25.26);ALT=T[chr14:65544631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65544756	+	chr14	65560425	+	.	0	16	5775607_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5775607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65537501_65562501_224C;SPAN=15669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:83 GQ:30.5 PL:[30.5, 0.0, 169.1] SR:16 DR:0 LR:-30.33 LO:35.97);ALT=T[chr14:65560425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65544790	+	chr14	65569020	+	.	9	0	5775916_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5775916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:65544790(+)-14:65569020(-)__14_65562001_65587001D;SPAN=24230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:45 GQ:17.6 PL:[17.6, 0.0, 90.2] SR:0 DR:9 LR:-17.52 LO:20.4);ALT=T[chr14:65569020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	65560533	+	chr14	65569021	+	.	0	14	5775917_1	34.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5775917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_65562001_65587001_229C;SPAN=8488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:45 GQ:34.1 PL:[34.1, 0.0, 73.7] SR:14 DR:0 LR:-34.02 LO:34.88);ALT=C[chr14:65569021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	797505	+	chr14	65745966	+	.	7	3	5776402_1	15.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=CGGGTCTGCTCTGTGTGCCATGGACGG;MAPQ=18;MATEID=5776402_2;MATENM=0;NM=5;NUMPARTS=2;SCTG=c_14_65733501_65758501_249C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:3 DR:7 LR:-15.3 LO:18.03);ALT=]chr19:797505]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr14	67810157	+	chr14	67812485	+	.	0	7	5781536_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5781536_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_67791501_67816501_136C;SPAN=2328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:7 DR:0 LR:-2.246 LO:13.27);ALT=T[chr14:67812485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	67817409	+	chr14	67819640	+	.	0	9	5781332_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5781332_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_67816001_67841001_251C;SPAN=2231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:9 DR:0 LR:-9.119 LO:18.15);ALT=T[chr14:67819640[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	67819757	+	chr14	67826374	+	.	0	13	5781342_1	19.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5781342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_67816001_67841001_229C;SPAN=6617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:86 GQ:19.7 PL:[19.7, 0.0, 188.0] SR:13 DR:0 LR:-19.61 LO:27.71);ALT=C[chr14:67826374[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	67827210	+	chr14	67831480	+	.	21	0	5781365_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5781365_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:67827210(+)-14:67831480(-)__14_67816001_67841001D;SPAN=4270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:74 GQ:49.4 PL:[49.4, 0.0, 128.6] SR:0 DR:21 LR:-49.27 LO:51.3);ALT=C[chr14:67831480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	68286621	+	chr14	68292178	+	.	8	0	5782820_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5782820_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:68286621(+)-14:68292178(-)__14_68281501_68306501D;SPAN=5557;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:72 GQ:7.1 PL:[7.1, 0.0, 165.5] SR:0 DR:8 LR:-6.901 LO:15.9);ALT=C[chr14:68292178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	69257211	+	chr14	69259598	+	.	0	7	5785073_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5785073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_69237001_69262001_308C;SPAN=2387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:73 GQ:3.5 PL:[3.5, 0.0, 171.8] SR:7 DR:0 LR:-3.33 LO:13.44);ALT=T[chr14:69259598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	69847373	+	chr14	69864947	+	.	15	0	5786812_1	26.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5786812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:69847373(+)-14:69864947(-)__14_69849501_69874501D;SPAN=17574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:84 GQ:26.9 PL:[26.9, 0.0, 175.4] SR:0 DR:15 LR:-26.76 LO:33.17);ALT=G[chr14:69864947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	69853826	+	chr14	69864946	+	.	65	0	5786822_1	99.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=5786822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:69853826(+)-14:69864946(-)__14_69849501_69874501D;SPAN=11120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:114 GQ:91.4 PL:[183.8, 0.0, 91.4] SR:0 DR:65 LR:-185.3 LO:185.3);ALT=A[chr14:69864946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	69861630	+	chr14	69864948	+	.	7	16	5786856_1	40.0	.	DISC_MAPQ=15;EVDNC=ASDIS;HOMSEQ=G;MAPQ=11;MATEID=5786856_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_69849501_69874501_248C;SPAN=3318;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:130 GQ:40.7 PL:[40.7, 0.0, 275.0] SR:16 DR:7 LR:-40.7 LO:50.76);ALT=C[chr14:69864948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70235651	+	chr14	70237181	+	.	10	0	5788233_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5788233_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:70235651(+)-14:70237181(-)__14_70217001_70242001D;SPAN=1530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:108 GQ:3.8 PL:[3.8, 0.0, 257.9] SR:0 DR:10 LR:-3.75 LO:19.04);ALT=G[chr14:70237181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70235969	+	chr14	70237711	+	ATCTCAAAGATTTCATGAGACAAGCTGGGGAAGTAACGTTTGCGGATGCACACCGACCTAAATTAAATGAAG	2	59	5788235_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATCTCAAAGATTTCATGAGACAAGCTGGGGAAGTAACGTTTGCGGATGCACACCGACCTAAATTAAATGAAG;MAPQ=60;MATEID=5788235_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_70217001_70242001_126C;SPAN=1742;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:95 GQ:53.6 PL:[175.7, 0.0, 53.6] SR:59 DR:2 LR:-179.1 LO:179.1);ALT=G[chr14:70237711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70793168	+	chr14	70826236	+	CATATTCCGACTCTAAAGATATTTTATTCTCTTTCAGTTTTTTTTCAAGCTCAGGATCCATTTTACTCTTCACAGCATCATATCGGATTTGAGAAAACTCACGAAGACCAAAAGAACCTCCAACAATCAGCAA	28	82	5789240_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATATTCCGACTCTAAAGATATTTTATTCTCTTTCAGTTTTTTTTCAAGCTCAGGATCCATTTTACTCTTCACAGCATCATATCGGATTTGAGAAAACTCACGAAGACCAAAAGAACCTCCAACAATCAGCAA;MAPQ=60;MATEID=5789240_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_14_70805001_70830001_241C;SPAN=33068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:104 DP:59 GQ:27.9 PL:[306.9, 27.9, 0.0] SR:82 DR:28 LR:-307.0 LO:307.0);ALT=T[chr14:70826236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70793168	+	chr14	70795891	+	.	2	30	5789160_1	82.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5789160_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ATAT;SCTG=c_14_70780501_70805501_335C;SPAN=2723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:85 GQ:82.7 PL:[82.7, 0.0, 122.3] SR:30 DR:2 LR:-82.6 LO:83.05);ALT=T[chr14:70795891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70796006	+	chr14	70826238	+	.	33	0	5789243_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5789243_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:70796006(+)-14:70826238(-)__14_70805001_70830001D;SPAN=30232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:61 GQ:53 PL:[92.6, 0.0, 53.0] SR:0 DR:33 LR:-92.9 LO:92.9);ALT=A[chr14:70826238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	70809487	+	chr14	70826295	+	.	40	0	5789253_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5789253_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:70809487(+)-14:70826295(-)__14_70805001_70830001D;SPAN=16808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:97 GQ:99 PL:[105.8, 0.0, 128.9] SR:0 DR:40 LR:-105.8 LO:105.9);ALT=C[chr14:70826295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	71060097	+	chr14	71064335	+	TGGGCAGGGGACTGCCGCTGTTGCTTCCGAATGATGAAAAGAATGGGCTCTTGAGCATGCAAAAGGATGTACTCGATTCCAACCATCTGA	0	18	5789881_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGGGCAGGGGACTGCCGCTGTTGCTTCCGAATGATGAAAAGAATGGGCTCTTGAGCATGCAAAAGGATGTACTCGATTCCAACCATCTGA;MAPQ=60;MATEID=5789881_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_71050001_71075001_137C;SPAN=4238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:76 GQ:38.9 PL:[38.9, 0.0, 144.5] SR:18 DR:0 LR:-38.83 LO:42.31);ALT=T[chr14:71064335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	71063464	+	chr14	71067332	+	.	11	0	5789891_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5789891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:71063464(+)-14:71067332(-)__14_71050001_71075001D;SPAN=3868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:78 GQ:15.2 PL:[15.2, 0.0, 173.6] SR:0 DR:11 LR:-15.18 LO:23.09);ALT=A[chr14:71067332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73525413	+	chr14	73538334	+	.	44	26	5795961_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5795961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73524501_73549501_277C;SPAN=12921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:96 GQ:79.7 PL:[152.3, 0.0, 79.7] SR:26 DR:44 LR:-153.4 LO:153.4);ALT=G[chr14:73538334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73525418	+	chr14	73543023	+	.	10	0	5795962_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5795962_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:73525418(+)-14:73543023(-)__14_73524501_73549501D;SPAN=17605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:0 DR:10 LR:-7.272 LO:19.63);ALT=G[chr14:73543023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73538456	+	chr14	73544077	+	GACCCCAATGATTCCTGTACCAATGAGCATTATGGCTCCTGCTCCAACT	0	23	5796013_1	56.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=GACCCCAATGATTCCTGTACCAATGAGCATTATGGCTCCTGCTCCAACT;MAPQ=60;MATEID=5796013_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_73524501_73549501_341C;SPAN=5621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:74 GQ:56 PL:[56.0, 0.0, 122.0] SR:23 DR:0 LR:-55.88 LO:57.29);ALT=G[chr14:73544077[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73563808	+	chr14	73566373	+	ATTTTCCGCAGATTTCCAGTGGCCCCACTGATCCCTTATCCACTCATCACTA	3	18	5796279_1	40.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATTTTCCGCAGATTTCCAGTGGCCCCACTGATCCCTTATCCACTCATCACTA;MAPQ=60;MATEID=5796279_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_73549001_73574001_194C;SPAN=2565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:84 GQ:40.1 PL:[40.1, 0.0, 162.2] SR:18 DR:3 LR:-39.96 LO:44.22);ALT=C[chr14:73566373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73563808	+	chr14	73566088	+	.	2	11	5796278_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=5796278_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_14_73549001_73574001_194C;SPAN=2280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:11 DR:2 LR:-17.4 LO:25.39);ALT=C[chr14:73566088[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73570186	+	chr14	73572565	+	.	7	22	5796305_1	58.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5796305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73549001_73574001_255C;SPAN=2379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:113 GQ:58.7 PL:[58.7, 0.0, 213.8] SR:22 DR:7 LR:-58.51 LO:63.58);ALT=G[chr14:73572565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73573041	+	chr14	73576041	+	.	12	0	5796318_1	31.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5796318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:73573041(+)-14:73576041(-)__14_73549001_73574001D;SPAN=3000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:29 GQ:31.7 PL:[31.7, 0.0, 38.3] SR:0 DR:12 LR:-31.76 LO:31.79);ALT=T[chr14:73576041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73576200	+	chr14	73577538	+	.	7	12	5796062_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5796062_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_73573501_73598501_227C;SPAN=1338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:99 GQ:29.3 PL:[29.3, 0.0, 210.8] SR:12 DR:7 LR:-29.3 LO:37.27);ALT=G[chr14:73577538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	73876772	+	chr14	73925198	+	.	9	0	5797544_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5797544_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:73876772(+)-14:73925198(-)__14_73867501_73892501D;SPAN=48426;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.6 LO:20.81);ALT=C[chr14:73925198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	81993310	+	chr14	82000019	+	TGGAATCTAAGGATTCATCCTGGCTGCCTTCTTCAT	0	8	5819459_1	0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TGGAATCTAAGGATTCATCCTGGCTGCCTTCTTCAT;MAPQ=60;MATEID=5819459_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_81977001_82002001_176C;SPAN=6709;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:104 GQ:1.5 PL:[0.0, 1.5, 254.1] SR:8 DR:0 LR:1.768 LO:14.56);ALT=T[chr14:82000019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	89953017	+	chr14	90085372	+	.	9	5	5837473_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5837473_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_90062001_90087001_45C;SPAN=132355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:49 GQ:19.7 PL:[19.7, 0.0, 98.9] SR:5 DR:9 LR:-19.73 LO:22.76);ALT=T[chr14:90085372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	90863578	+	chr14	90867602	+	CTGATCAGCTGACCGAAGAACAGATTGCT	39	211	5839807_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=CTGATCAGCTGACCGAAGAACAGATTGCT;MAPQ=60;MATEID=5839807_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_90846001_90871001_177C;SPAN=4024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:232 DP:135 GQ:62.5 PL:[686.5, 62.5, 0.0] SR:211 DR:39 LR:-686.6 LO:686.6);ALT=G[chr14:90867602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	90867750	+	chr14	90870205	+	.	5	47	5839819_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTAA;MAPQ=60;MATEID=5839819_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_90846001_90871001_282C;SPAN=2455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:113 GQ:99 PL:[134.6, 0.0, 137.9] SR:47 DR:5 LR:-134.4 LO:134.4);ALT=A[chr14:90870205[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	91580628	+	chr14	91626608	+	AGCCAAGTTACACCCTGTTTAACCCTGCCTTCAAAGGGACGACTCTGTA	0	13	5841925_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGCCAAGTTACACCCTGTTTAACCCTGCCTTCAAAGGGACGACTCTGTA;MAPQ=60;MATEID=5841925_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_91605501_91630501_51C;SPAN=45980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:49 GQ:29.6 PL:[29.6, 0.0, 89.0] SR:13 DR:0 LR:-29.64 LO:31.3);ALT=G[chr14:91626608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	91624034	+	chr14	91626608	+	.	2	9	5841985_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5841985_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_14_91605501_91630501_51C;SPAN=2574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:9 DR:2 LR:-4.834 LO:19.21);ALT=G[chr14:91626608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	91929222	+	chr14	91931593	+	.	2	3	5842678_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5842678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_91924001_91949001_267C;SPAN=2371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:3 DR:2 LR:6.574 LO:6.671);ALT=C[chr14:91931593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	91982027	+	chr17	28483267	+	.	20	65	6359574_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6359574_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_17_28469001_28494001_373C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:38 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:65 DR:20 LR:-217.9 LO:217.9);ALT=T[chr17:28483267[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr14	92582606	+	chr14	92587985	+	.	13	0	5844816_1	22.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5844816_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:92582606(+)-14:92587985(-)__14_92585501_92610501D;SPAN=5379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:75 GQ:22.7 PL:[22.7, 0.0, 158.0] SR:0 DR:13 LR:-22.59 LO:28.56);ALT=A[chr14:92587985[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	92584254	+	chr14	92587983	+	.	22	0	5844723_1	60.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=5844723_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:92584254(+)-14:92587983(-)__14_92561001_92586001D;SPAN=3729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:45 GQ:47.3 PL:[60.5, 0.0, 47.3] SR:0 DR:22 LR:-60.5 LO:60.5);ALT=A[chr14:92587983[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	92588472	+	chr14	92597295	+	ATTAATAAAGAACTCTTCAGAATTCCTGGTGTTTCATCATATATACGACTAAGATATCA	6	8	5844840_1	7.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATTAATAAAGAACTCTTCAGAATTCCTGGTGTTTCATCATATATACGACTAAGATATCA;MAPQ=60;MATEID=5844840_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_92585501_92610501_240C;SPAN=8823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:8 DR:6 LR:-7.272 LO:19.63);ALT=G[chr14:92597295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	93651429	+	chr14	93652600	+	.	16	0	5847763_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5847763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:93651429(+)-14:93652600(-)__14_93639001_93664001D;SPAN=1171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:73 GQ:33.2 PL:[33.2, 0.0, 142.1] SR:0 DR:16 LR:-33.04 LO:36.98);ALT=C[chr14:93652600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	93670128	+	chr14	93673171	+	.	0	10	5848003_1	8.0	.	EVDNC=ASSMB;HOMSEQ=TCACC;MAPQ=60;MATEID=5848003_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_93663501_93688501_56C;SPAN=3043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:10 DR:0 LR:-8.898 LO:19.93);ALT=C[chr14:93673171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	94546110	+	chr14	94547464	+	.	50	0	5850020_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5850020_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:94546110(+)-14:94547464(-)__14_94521001_94546001D;SPAN=1354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:0 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=T[chr14:94547464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	94547797	+	chr14	94563233	+	.	12	4	5849898_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=5849898_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_94545501_94570501_151C;SPAN=15436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:4 DR:12 LR:-21.73 LO:26.64);ALT=T[chr14:94563233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	94563312	+	chr14	94568158	+	CAGGGCTGCTGTAGCAGCTGTGGTCGGAGG	0	12	5849928_1	15.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAGGGCTGCTGTAGCAGCTGTGGTCGGAGG;MAPQ=60;MATEID=5849928_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_94545501_94570501_288C;SPAN=4846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:12 DR:0 LR:-15.23 LO:24.87);ALT=G[chr14:94568158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	94849580	+	chr14	94856793	+	.	0	30	5850777_1	71.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5850777_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_94839501_94864501_279C;SPAN=7213;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:102 GQ:71.6 PL:[71.6, 0.0, 173.9] SR:30 DR:0 LR:-71.4 LO:73.85);ALT=T[chr14:94856793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	95591007	+	chr14	95592917	+	.	3	2	5852797_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5852797_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_95574501_95599501_287C;SPAN=1910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:68 GQ:5.1 PL:[0.0, 5.1, 174.9] SR:2 DR:3 LR:5.219 LO:6.798);ALT=T[chr14:95592917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	102411135	-	chr14	102412154	+	.	8	0	5870132_1	0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=5870132_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:102411135(-)-14:102412154(-)__14_102410001_102435001D;SPAN=1019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr14:102412154[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	102822234	+	chr14	102825755	+	.	0	16	5871513_1	34.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5871513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_102802001_102827001_59C;SPAN=3521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:69 GQ:34.1 PL:[34.1, 0.0, 133.1] SR:16 DR:0 LR:-34.12 LO:37.43);ALT=C[chr14:102825755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	102822281	+	chr14	102829181	+	.	11	0	5871515_1	28.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=5871515_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:102822281(+)-14:102829181(-)__14_102802001_102827001D;SPAN=6900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:29 GQ:28.4 PL:[28.4, 0.0, 41.6] SR:0 DR:11 LR:-28.45 LO:28.6);ALT=T[chr14:102829181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	102825915	+	chr14	102829181	+	.	16	0	5871522_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5871522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:102825915(+)-14:102829181(-)__14_102802001_102827001D;SPAN=3266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:40 GQ:41.9 PL:[41.9, 0.0, 55.1] SR:0 DR:16 LR:-41.98 LO:42.08);ALT=A[chr14:102829181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	103334546	+	chr14	103333448	+	.	2	5	5873012_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CCTCTG;MAPQ=60;MATEID=5873012_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_103316501_103341501_148C;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:5 DR:2 LR:1.055 LO:10.95);ALT=]chr14:103334546]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	103388545	+	chr14	103386206	+	.	10	0	5873280_1	7.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5873280_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:103386206(-)-14:103388545(+)__14_103365501_103390501D;SPAN=2339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:0 DR:10 LR:-7.272 LO:19.63);ALT=]chr14:103388545]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	103590289	+	chr14	103592644	+	.	7	15	5873870_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5873870_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_103586001_103611001_72C;SPAN=2355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:58 GQ:47 PL:[47.0, 0.0, 93.2] SR:15 DR:7 LR:-47.01 LO:47.86);ALT=G[chr14:103592644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	103800934	+	chr14	103801989	+	.	32	37	5874493_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5874493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_103782001_103807001_337C;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:37 DR:32 LR:-163.7 LO:163.7);ALT=G[chr14:103801989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	103958371	+	chr14	103969217	+	.	4	3	5875111_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5875111_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_103953501_103978501_282C;SPAN=10846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:3 DR:4 LR:1.547 LO:12.74);ALT=G[chr14:103969217[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104029463	+	chr14	104037959	+	.	29	13	5875491_1	83.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5875491_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_104027001_104052001_207C;SPAN=8496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:84 GQ:83 PL:[83.0, 0.0, 119.3] SR:13 DR:29 LR:-82.88 LO:83.27);ALT=T[chr14:104037959[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104379035	+	chr14	104381403	+	CAAAGCCTTACTTCTTTTAT	0	148	5876589_1	99.0	.	EVDNC=ASSMB;INSERTION=CAAAGCCTTACTTCTTTTAT;MAPQ=60;MATEID=5876589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_104370001_104395001_12C;SPAN=2368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:148 DP:240 GQ:99 PL:[423.5, 0.0, 159.4] SR:148 DR:0 LR:-430.1 LO:430.1);ALT=T[chr14:104381403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104379095	+	chr14	104387803	+	.	75	0	5876590_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5876590_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:104379095(+)-14:104387803(-)__14_104370001_104395001D;SPAN=8708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:176 GQ:99 PL:[200.0, 0.0, 226.4] SR:0 DR:75 LR:-199.9 LO:200.0);ALT=A[chr14:104387803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104381528	+	chr14	104387807	+	.	62	3	5876599_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5876599_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_104370001_104395001_319C;SPAN=6279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:241 GQ:99 PL:[146.2, 0.0, 436.7] SR:3 DR:62 LR:-146.0 LO:154.1);ALT=T[chr14:104387807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	104791597	+	chr14	104790597	+	.	26	0	5877490_1	61.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5877490_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:104790597(-)-14:104791597(+)__14_104786501_104811501D;SPAN=1000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:91 GQ:61.4 PL:[61.4, 0.0, 157.1] SR:0 DR:26 LR:-61.17 LO:63.6);ALT=]chr14:104791597]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	105156041	+	chr14	105167690	+	.	10	0	5878426_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5878426_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105156041(+)-14:105167690(-)__14_105154001_105179001D;SPAN=11649;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:0 DR:10 LR:-18.65 LO:22.38);ALT=G[chr14:105167690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105219656	+	chr14	105221966	+	.	115	62	5878785_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5878785_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_105203001_105228001_34C;SPAN=2310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:81 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:62 DR:115 LR:-422.5 LO:422.5);ALT=G[chr14:105221966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105219688	+	chr14	105222939	+	.	11	0	5878786_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5878786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105219688(+)-14:105222939(-)__14_105203001_105228001D;SPAN=3251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:0 DR:11 LR:-15.99 LO:23.29);ALT=T[chr14:105222939[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105222161	+	chr14	105225765	+	ACCCATCTGGGGTAGCGTCCATTGCCTGTTCCTCATGCGTGCGAGCCGTGGATGGGAAGGCGGTCTGCGGTCAGTGTGAGCGAGCCCTGTGCGGGCAGTGTGTGCGCACCTGCTGGGGCTGCGGCTCCGTGGCCTGTACCCTGTGTGGCCTCGTGGA	0	76	5878793_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACCCATCTGGGGTAGCGTCCATTGCCTGTTCCTCATGCGTGCGAGCCGTGGATGGGAAGGCGGTCTGCGGTCAGTGTGAGCGAGCCCTGTGCGGGCAGTGTGTGCGCACCTGCTGGGGCTGCGGCTCCGTGGCCTGTACCCTGTGTGGCCTCGTGGA;MAPQ=60;MATEID=5878793_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_14_105203001_105228001_112C;SPAN=3604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:76 DP:122 GQ:76.1 PL:[218.0, 0.0, 76.1] SR:76 DR:0 LR:-221.4 LO:221.4);ALT=G[chr14:105225765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105391327	+	chr14	105393476	+	.	45	9	5879068_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5879068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_105374501_105399501_235C;SPAN=2149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:87 GQ:55.7 PL:[154.7, 0.0, 55.7] SR:9 DR:45 LR:-157.2 LO:157.2);ALT=G[chr14:105393476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105417220	+	chr14	105418257	+	.	31	0	5879124_1	92.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=5879124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105417220(+)-14:105418257(-)__14_105399001_105424001D;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=A[chr14:105418257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105478305	+	chr14	105487348	+	.	10	0	5879534_1	18.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5879534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105478305(+)-14:105487348(-)__14_105472501_105497501D;SPAN=9043;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:0 DR:10 LR:-18.65 LO:22.38);ALT=A[chr14:105487348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	105953618	+	chr14	105954996	+	.	22	0	5880804_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5880804_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:105953618(+)-14:105954996(-)__14_105938001_105963001D;SPAN=1378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:22 DP:326 GQ:15.5 PL:[0.0, 15.5, 821.9] SR:0 DR:22 LR:15.7 LO:38.74);ALT=A[chr14:105954996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106227280	+	chr14	106082685	+	AC	35	63	5882176_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=AC;MAPQ=35;MATEID=5882176_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_14_106207501_106232501_108C;SPAN=144595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:107 GQ:7.4 PL:[251.6, 0.0, 7.4] SR:63 DR:35 LR:-265.4 LO:265.4);ALT=]chr14:106227280]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106089348	+	chr14	106133062	+	.	9	15	5881552_1	62.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GTGGGGGACAGCGTCAGGGACAG;MAPQ=60;MATEID=5881552_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_14_106085001_106110001_208C;SPAN=43714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:63 GQ:62.3 PL:[62.3, 0.0, 88.7] SR:15 DR:9 LR:-62.16 LO:62.45);ALT=G[chr14:106133062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106096441	+	chr14	106115536	+	.	12	0	5881613_1	31.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5881613_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106096441(+)-14:106115536(-)__14_106085001_106110001D;SPAN=19095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:29 GQ:31.7 PL:[31.7, 0.0, 38.3] SR:0 DR:12 LR:-31.76 LO:31.79);ALT=A[chr14:106115536[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106115778	+	chr14	106096963	+	.	84	0	5881616_1	99.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5881616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106096963(-)-14:106115778(+)__14_106085001_106110001D;SPAN=18815;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:49 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:0 DR:84 LR:-247.6 LO:247.6);ALT=]chr14:106115778]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	106217127	+	chr14	106315364	-	.	10	0	5882520_1	29.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=5882520_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106217127(+)-14:106315364(+)__14_106305501_106330501D;SPAN=98237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:10 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:10 LR:-29.71 LO:29.71);ALT=A]chr14:106315364];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	106346009	+	chr14	106386922	+	.	41	6	5882731_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=5882731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106379001_106404001_249C;SPAN=40913;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:56 GQ:8 PL:[126.8, 0.0, 8.0] SR:6 DR:41 LR:-132.8 LO:132.8);ALT=A[chr14:106386922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106356056	+	chr14	106361841	+	.	8	3	5882617_1	9.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=G;MAPQ=47;MATEID=5882617_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106354501_106379501_288C;SPAN=5785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:3 DR:8 LR:-9.711 LO:20.09);ALT=G[chr14:106361841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106356069	+	chr14	106362160	+	.	17	0	5882618_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5882618_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106356069(+)-14:106362160(-)__14_106354501_106379501D;SPAN=6091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:84 GQ:33.5 PL:[33.5, 0.0, 168.8] SR:0 DR:17 LR:-33.36 LO:38.63);ALT=T[chr14:106362160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106365505	+	chr14	106386922	+	.	12	4	5882736_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5882736_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106379001_106404001_330C;SECONDARY;SPAN=21417;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:56 GQ:34.4 PL:[34.4, 0.0, 100.4] SR:4 DR:12 LR:-34.34 LO:36.19);ALT=C[chr14:106386922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106374811	+	chr14	106386920	+	.	36	8	5882739_1	99.0	.	DISC_MAPQ=27;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5882739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_106379001_106404001_2C;SPAN=12109;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:53 GQ:0.9 PL:[128.7, 0.9, 0.0] SR:8 DR:36 LR:-135.3 LO:135.3);ALT=G[chr14:106386920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106650158	+	chr14	106841885	+	.	14	0	5884157_1	28.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=5884157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106650158(+)-14:106841885(-)__14_106820001_106845001D;SPAN=191727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:67 GQ:28.1 PL:[28.1, 0.0, 133.7] SR:0 DR:14 LR:-28.06 LO:32.03);ALT=C[chr14:106841885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr14	106842059	+	chr14	106650352	+	.	20	0	5884158_1	51.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=5884158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106650352(-)-14:106842059(+)__14_106820001_106845001D;SPAN=191707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:55 GQ:51.2 PL:[51.2, 0.0, 80.9] SR:0 DR:20 LR:-51.12 LO:51.52);ALT=]chr14:106842059]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr14	107011557	+	chr14	106713111	+	.	10	0	5883646_1	20.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5883646_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=14:106713111(-)-14:107011557(+)__14_106697501_106722501D;SPAN=298446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=]chr14:107011557]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	23671438	+	chr15	23675199	+	.	39	11	5901087_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=GGCACGGTGGCTCACGCCTGTAATCCCAGCACTTTGGGAGGCCAAGG;MAPQ=60;MATEID=5901087_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_23667001_23692001_111C;SPAN=3761;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:77 GQ:45.2 PL:[140.9, 0.0, 45.2] SR:11 DR:39 LR:-143.5 LO:143.5);ALT=G[chr15:23675199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	23685607	-	chr20	37274467	+	.	20	18	5901158_1	90.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=G;MAPQ=28;MATEID=5901158_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_15_23667001_23692001_475C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:56 GQ:44.3 PL:[90.5, 0.0, 44.3] SR:18 DR:20 LR:-91.26 LO:91.26);ALT=[chr20:37274467[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr20	37274667	+	chr15	23706879	+	.	16	16	5902570_1	81.0	.	DISC_MAPQ=38;EVDNC=ASDIS;MAPQ=60;MATEID=5902570_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_23691501_23716501_706C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:53 GQ:45.2 PL:[81.5, 0.0, 45.2] SR:16 DR:16 LR:-81.86 LO:81.86);ALT=]chr20:37274667]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr15	23712660	+	chr15	23717165	+	.	17	0	5902610_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5902610_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:23712660(+)-15:23717165(-)__15_23691501_23716501D;SPAN=4505;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:58 GQ:40.4 PL:[40.4, 0.0, 99.8] SR:0 DR:17 LR:-40.4 LO:41.81);ALT=A[chr15:23717165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	23831701	+	chr15	23992755	-	.	29	0	5902351_1	85.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5902351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:23831701(+)-15:23992755(+)__15_23985501_24010501D;SPAN=161054;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:24 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:0 DR:29 LR:-85.82 LO:85.82);ALT=T]chr15:23992755];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr15	24761591	+	chr15	24454832	+	.	10	0	5903373_1	25.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5903373_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:24454832(-)-15:24761591(+)__15_24451001_24476001D;SPAN=306759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:28 GQ:25.4 PL:[25.4, 0.0, 41.9] SR:0 DR:10 LR:-25.42 LO:25.66);ALT=]chr15:24761591]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	24802670	+	chr15	24588040	+	.	9	1	5904310_1	26.0	.	DISC_MAPQ=19;EVDNC=ASDIS;HOMSEQ=GCCCCAACAGCACATCAACTTCATCCCAGGTCCATG;MAPQ=0;MATEID=5904310_2;MATENM=1;NM=0;NUMPARTS=2;REPSEQ=CCCC;SCTG=c_15_24794001_24819001_61C;SECONDARY;SPAN=214630;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:1 DR:9 LR:-26.78 LO:26.78);ALT=]chr15:24802670]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	24593127	-	chr15	24647420	+	.	4	4	5903936_1	16.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=TCCATGCAGTGA;MAPQ=38;MATEID=5903936_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_24647001_24672001_137C;SPAN=54293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:37 GQ:16.4 PL:[16.4, 0.0, 72.5] SR:4 DR:4 LR:-16.38 LO:18.44);ALT=[chr15:24647420[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	24816543	+	chr15	24643432	+	.	8	0	5903808_1	18.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5903808_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:24643432(-)-15:24816543(+)__15_24622501_24647501D;SPAN=173111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=]chr15:24816543]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	35529517	-	chr15	69113095	+	.	32	0	5979459_1	93.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=5979459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:35529517(-)-15:69113095(-)__15_69090001_69115001D;SPAN=33583578;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:44 GQ:11.3 PL:[93.8, 0.0, 11.3] SR:0 DR:32 LR:-97.22 LO:97.22);ALT=[chr15:69113095[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	35830670	+	chr15	35834614	+	.	0	11	5924605_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5924605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_35819001_35844001_80C;SPAN=3944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:65 GQ:18.8 PL:[18.8, 0.0, 137.6] SR:11 DR:0 LR:-18.7 LO:24.04);ALT=T[chr15:35834614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	35830717	+	chr15	35838319	+	.	15	0	5924606_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5924606_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:35830717(+)-15:35838319(-)__15_35819001_35844001D;SPAN=7602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:0 DR:15 LR:-32.72 LO:35.42);ALT=A[chr15:35838319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	39372395	+	chr15	39373461	+	.	43	34	5929389_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=TTCTCCTGCCTCAGCCTCCCGAGTAGCTGGGATTACAGGCA;MAPQ=60;MATEID=5929389_2;MATENM=5;NM=1;NUMPARTS=2;SCTG=c_15_39371501_39396501_138C;SPAN=1066;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:6 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:34 DR:43 LR:-221.2 LO:221.2);ALT=A[chr15:39373461[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40226471	+	chr15	40231704	+	.	18	0	5930510_1	56.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5930510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:40226471(+)-15:40231704(-)__15_40229001_40254001D;SPAN=5233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:19 GQ:5.1 PL:[56.1, 5.1, 0.0] SR:0 DR:18 LR:-56.11 LO:56.11);ALT=C[chr15:40231704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40231818	+	chr15	40235584	+	.	0	10	5930513_1	17.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5930513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40229001_40254001_90C;SPAN=3766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:10 DR:0 LR:-17.84 LO:22.11);ALT=T[chr15:40235584[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40235688	+	chr15	40241315	+	.	0	33	5930528_1	89.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5930528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40229001_40254001_200C;SPAN=5627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:73 GQ:86 PL:[89.3, 0.0, 86.0] SR:33 DR:0 LR:-89.16 LO:89.16);ALT=T[chr15:40241315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40328700	+	chr15	40331293	+	.	20	0	5930680_1	37.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=5930680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:40328700(+)-15:40331293(-)__15_40327001_40352001D;SPAN=2593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:107 GQ:37.1 PL:[37.1, 0.0, 221.9] SR:0 DR:20 LR:-37.03 LO:44.67);ALT=G[chr15:40331293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40331651	+	chr15	40338159	+	.	6	5	5930691_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=5930691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40327001_40352001_177C;SPAN=6508;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:5 DR:6 LR:-10.97 LO:16.77);ALT=T[chr15:40338159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40596279	+	chr15	40599789	+	.	0	11	5931175_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5931175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40572001_40597001_26C;SPAN=3510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:25 GQ:29.6 PL:[29.6, 0.0, 29.6] SR:11 DR:0 LR:-29.54 LO:29.54);ALT=C[chr15:40599789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40698172	+	chr15	40699835	+	.	0	13	5931390_1	26.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5931390_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_40694501_40719501_259C;SPAN=1663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:13 DR:0 LR:-26.66 LO:29.98);ALT=G[chr15:40699835[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40699927	+	chr15	40702826	+	AATTTTGGAAGCAGCTGGGGAACCTGGGCGTATTGGGCATCACAGCCCCT	0	11	5931400_1	21.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AATTTTGGAAGCAGCTGGGGAACCTGGGCGTATTGGGCATCACAGCCCCT;MAPQ=60;MATEID=5931400_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_40694501_40719501_244C;SPAN=2899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:11 DR:0 LR:-21.68 LO:25.03);ALT=G[chr15:40702826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	40855255	+	chr15	40857131	+	.	18	0	5931772_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5931772_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:40855255(+)-15:40857131(-)__15_40841501_40866501D;SPAN=1876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:50 GQ:45.8 PL:[45.8, 0.0, 75.5] SR:0 DR:18 LR:-45.87 LO:46.27);ALT=A[chr15:40857131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41056415	+	chr15	41058024	+	.	7	4	5932091_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=5932091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41037501_41062501_64C;SPAN=1609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:60 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:4 DR:7 LR:-13.45 LO:19.15);ALT=G[chr15:41058024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41058119	+	chr15	41059424	+	.	0	12	5932093_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5932093_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41037501_41062501_240C;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:58 GQ:23.9 PL:[23.9, 0.0, 116.3] SR:12 DR:0 LR:-23.9 LO:27.4);ALT=T[chr15:41059424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41068826	+	chr15	41071421	+	.	0	9	5932113_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5932113_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41062001_41087001_134C;SPAN=2595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:9 DR:0 LR:-14.27 LO:19.37);ALT=C[chr15:41071421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41072197	+	chr15	41099565	+	.	5	3	5932222_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=5932222_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_15_41086501_41111501_202C;SPAN=27368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:33 GQ:11 PL:[11.0, 0.0, 67.1] SR:3 DR:5 LR:-10.87 LO:13.32);ALT=T[chr15:41099565[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41388553	+	chr15	41408171	+	.	2	2	5932884_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5932884_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41405001_41430001_303C;SPAN=19618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:15 GQ:9.2 PL:[9.2, 0.0, 25.7] SR:2 DR:2 LR:-9.14 LO:9.642);ALT=T[chr15:41408171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41523647	+	chr15	41535865	+	.	7	8	5933145_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=5933145_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_15_41527501_41552501_166C;SPAN=12218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:24 GQ:26.6 PL:[29.9, 0.0, 26.6] SR:8 DR:7 LR:-29.81 LO:29.81);ALT=T[chr15:41535865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41523647	+	chr15	41549105	+	TTTCCCACAGTCAAATCACTCGCCTCTACAGCCGGTTCACCAGCCTGGACAAAGGAGAGAATGGGACTCT	2	11	5933146_1	34.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=TTTCCCACAGTCAAATCACTCGCCTCTACAGCCGGTTCACCAGCCTGGACAAAGGAGAGAATGGGACTCT;MAPQ=60;MATEID=5933146_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_41527501_41552501_166C;SPAN=25458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:30 GQ:34.7 PL:[34.7, 0.0, 38.0] SR:11 DR:2 LR:-34.79 LO:34.79);ALT=T[chr15:41549105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41576309	+	chr15	41577421	+	.	40	14	5933342_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5933342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41576501_41601501_263C;SPAN=1112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:46 DP:31 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:14 DR:40 LR:-135.3 LO:135.3);ALT=G[chr15:41577421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41628510	+	chr15	41621292	+	.	19	22	5933519_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ATAA;MAPQ=60;MATEID=5933519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41601001_41626001_254C;SPAN=7218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:23 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:22 DR:19 LR:-115.5 LO:115.5);ALT=]chr15:41628510]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	41634653	+	chr15	41641292	+	.	0	7	5933424_1	8.0	.	EVDNC=ASSMB;HOMSEQ=TCAGG;MAPQ=60;MATEID=5933424_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41625501_41650501_130C;SPAN=6639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:54 GQ:8.6 PL:[8.6, 0.0, 120.8] SR:7 DR:0 LR:-8.477 LO:14.41);ALT=G[chr15:41641292[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41709512	+	chr15	41730517	+	.	44	56	5933821_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5933821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_41699001_41724001_208C;SPAN=21005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:38 GQ:18 PL:[198.0, 18.0, 0.0] SR:56 DR:44 LR:-198.0 LO:198.0);ALT=G[chr15:41730517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41730629	+	chr15	41745097	+	.	2	9	5933677_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5933677_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_15_41723501_41748501_330C;SPAN=14468;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:9 DR:2 LR:-16.75 LO:21.78);ALT=G[chr15:41745097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41730629	+	chr15	41749868	+	TGGACATTTGGGAGCAATAAAAATAAGAAGAAAGGAAAAGCCAGAAAAATAGAGAAGAAAGGAACCATGAAGAAACAGGCCAACAAAACTGCCTCCTCAGGCAGTTCAGACAAAGACAGTTCAGCTGAGAGCTCAGCCCCTGAGGA	0	55	5933678_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGTGA;INSERTION=TGGACATTTGGGAGCAATAAAAATAAGAAGAAAGGAAAAGCCAGAAAAATAGAGAAGAAAGGAACCATGAAGAAACAGGCCAACAAAACTGCCTCCTCAGGCAGTTCAGACAAAGACAGTTCAGCTGAGAGCTCAGCCCCTGAGGA;MAPQ=60;MATEID=5933678_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_41723501_41748501_330C;SPAN=19239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:31 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:55 DR:0 LR:-161.7 LO:161.7);ALT=G[chr15:41749868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	41745250	+	chr15	41749868	+	.	6	40	5933592_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGTGA;MAPQ=60;MATEID=5933592_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GTGT;SCTG=c_15_41748001_41773001_89C;SPAN=4618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:48 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:40 DR:6 LR:-141.9 LO:141.9);ALT=A[chr15:41749868[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42120398	+	chr15	42126936	+	.	15	0	5934556_1	32.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=5934556_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:42120398(+)-15:42126936(-)__15_42115501_42140501D;SPAN=6538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:63 GQ:32.6 PL:[32.6, 0.0, 118.4] SR:0 DR:15 LR:-32.45 LO:35.29);ALT=T[chr15:42126936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42560230	+	chr15	42565452	+	ACTTCAGGAAGATAGTGGTATTTCTGAAGAGGATCTTTCCAAAACTAAAATAATTTTTCC	0	12	5935319_1	25.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=ACTTCAGGAAGATAGTGGTATTTCTGAAGAGGATCTTTCCAAAACTAAAATAATTTTTCC;MAPQ=60;MATEID=5935319_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_42556501_42581501_255C;SPAN=5222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:12 DR:0 LR:-25.25 LO:27.93);ALT=A[chr15:42565452[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42787911	+	chr15	42804030	+	.	5	3	5935899_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5935899_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_15_42777001_42802001_124C;SPAN=16119;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:42 GQ:5.3 PL:[5.3, 0.0, 94.4] SR:3 DR:5 LR:-5.126 LO:10.1);ALT=G[chr15:42804030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42787961	+	chr15	42807433	+	.	14	0	5935902_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5935902_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:42787961(+)-15:42807433(-)__15_42777001_42802001D;SPAN=19472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:28 GQ:28.7 PL:[38.6, 0.0, 28.7] SR:0 DR:14 LR:-38.7 LO:38.7);ALT=G[chr15:42807433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42805645	+	chr15	42807434	+	.	0	10	5935757_1	17.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5935757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42801501_42826501_282C;SPAN=1789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:10 DR:0 LR:-17.3 LO:21.94);ALT=G[chr15:42807434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42807552	+	chr15	42820456	+	.	4	6	5935762_1	13.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ATAG;MAPQ=60;MATEID=5935762_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42801501_42826501_202C;SPAN=12904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:6 DR:4 LR:-13.67 LO:17.51);ALT=G[chr15:42820456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42841139	+	chr15	42853466	+	.	10	0	5935945_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5935945_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:42841139(+)-15:42853466(-)__15_42850501_42875501D;SPAN=12327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:23 GQ:26.9 PL:[26.9, 0.0, 26.9] SR:0 DR:10 LR:-26.78 LO:26.78);ALT=C[chr15:42853466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42841164	+	chr15	42850394	+	.	9	6	5935946_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5935946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42850501_42875501_19C;SPAN=9230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:0 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:6 DR:9 LR:-29.71 LO:29.71);ALT=G[chr15:42850394[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42851606	+	chr15	42853467	+	.	0	11	5935959_1	21.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5935959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42850501_42875501_267C;SPAN=1861;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:55 GQ:21.5 PL:[21.5, 0.0, 110.6] SR:11 DR:0 LR:-21.41 LO:24.93);ALT=G[chr15:42853467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	42851606	+	chr15	42852979	+	.	0	5	5935958_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5935958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_42850501_42875501_68C;SPAN=1373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:64 GQ:0.6 PL:[0.0, 0.6, 155.1] SR:5 DR:0 LR:0.8342 LO:9.134);ALT=G[chr15:42852979[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	43368155	-	chr20	5268410	+	AGAGGGC	16	29	5936976_1	99.0	.	DISC_MAPQ=6;EVDNC=ASDIS;INSERTION=AGAGGGC;MAPQ=14;MATEID=5936976_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_15_43365001_43390001_64C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:29 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:29 DR:16 LR:-125.4 LO:125.4);ALT=[chr20:5268410[C;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr15	43809939	+	chr15	43813167	+	.	19	0	5937747_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5937747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:43809939(+)-15:43813167(-)__15_43806001_43831001D;SPAN=3228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:52 GQ:48.8 PL:[48.8, 0.0, 75.2] SR:0 DR:19 LR:-48.63 LO:48.99);ALT=T[chr15:43813167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	44084833	+	chr15	44085888	+	.	209	0	5938738_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5938738_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:44084833(+)-15:44085888(-)__15_44075501_44100501D;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:209 DP:77 GQ:56.5 PL:[620.5, 56.5, 0.0] SR:0 DR:209 LR:-620.6 LO:620.6);ALT=G[chr15:44085888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	44109648	+	chr15	44116687	+	.	0	7	5938445_1	7.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=5938445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_44100001_44125001_92C;SPAN=7039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:58 GQ:7.4 PL:[7.4, 0.0, 132.8] SR:7 DR:0 LR:-7.393 LO:14.18);ALT=T[chr15:44116687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	44829435	+	chr15	44843072	+	ACGCCGACGCTTTCTCCGTGGAAGACCCAGTGCGGAAGGTGGGGGGCGGCGGCACTGCCGGCGGGGACCGCTGGGAAGGCGAGGACGAGGACGAGGACGTCA	8	43	5940209_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACGCCGACGCTTTCTCCGTGGAAGACCCAGTGCGGAAGGTGGGGGGCGGCGGCACTGCCGGCGGGGACCGCTGGGAAGGCGAGGACGAGGACGAGGACGTCA;MAPQ=60;MATEID=5940209_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_15_44810501_44835501_250C;SECONDARY;SPAN=13637;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:32 GQ:12 PL:[132.0, 12.0, 0.0] SR:43 DR:8 LR:-132.0 LO:132.0);ALT=G[chr15:44843072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45007899	+	chr15	45009803	+	ATCGAGACATGTAAGCAGCATCATGG	19	90	5940751_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=ATCGAGACATGTAAGCAGCATCATGG;MAPQ=60;MATEID=5940751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_45006501_45031501_235C;SPAN=1904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:101 DP:267 GQ:99 PL:[261.1, 0.0, 386.6] SR:90 DR:19 LR:-261.1 LO:262.4);ALT=G[chr15:45009803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45008609	+	chr15	45009836	+	.	8	0	5940752_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5940752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:45008609(+)-15:45009836(-)__15_45006501_45031501D;SPAN=1227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:229 GQ:35.5 PL:[0.0, 35.5, 627.1] SR:0 DR:8 LR:35.63 LO:11.76);ALT=A[chr15:45009836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45448743	-	chr15	45449776	+	.	8	0	5941337_1	13.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=5941337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:45448743(-)-15:45449776(-)__15_45447501_45472501D;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=[chr15:45449776[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	45879725	+	chr15	45884332	+	.	8	3	5942120_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=5942120_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_45864001_45889001_21C;SPAN=4607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:62 GQ:13.1 PL:[13.1, 0.0, 135.2] SR:3 DR:8 LR:-12.91 LO:19.01);ALT=T[chr15:45884332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45927306	+	chr15	45954151	+	CCTGATCCTGCCTGAAGATGGTGCCACTGGTGGCTGTGGTATCAGGGCCCCGTGCCCAGCTCTTTGCCTGCCTGCTCAGGCTGGGCACTCAGCAGGTCGGCCCCCTTCAGCTGCACACCGGGGCCAGCCATGCGGCCAGGAACCATTATGAGGTGCTGGTGCTGGGTGGGGGCAGTGGCGGAATCACCATGGCTGCCCGCATGAAGAGGAAAGTGGGTGCAGAGAATGTGGCCATTGTTGAGCCCAGTG	3	11	5942279_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCTGATCCTGCCTGAAGATGGTGCCACTGGTGGCTGTGGTATCAGGGCCCCGTGCCCAGCTCTTTGCCTGCCTGCTCAGGCTGGGCACTCAGCAGGTCGGCCCCCTTCAGCTGCACACCGGGGCCAGCCATGCGGCCAGGAACCATTATGAGGTGCTGGTGCTGGGTGGGGGCAGTGGCGGAATCACCATGGCTGCCCGCATGAAGAGGAAAGTGGGTGCAGAGAATGTGGCCATTGTTGAGCCCAGTG;MAPQ=60;MATEID=5942279_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_45913001_45938001_146C;SPAN=26845;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:42 GQ:25.1 PL:[25.1, 0.0, 74.6] SR:11 DR:3 LR:-24.93 LO:26.41);ALT=G[chr15:45954151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45927306	+	chr15	45951104	+	.	46	4	5942278_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5942278_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_15_45913001_45938001_146C;SPAN=23798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:42 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:4 DR:46 LR:-138.6 LO:138.6);ALT=G[chr15:45951104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45951355	+	chr15	45954151	+	.	4	6	5942236_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5942236_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_45937501_45962501_205C;SPAN=2796;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:6 DR:4 LR:-17.03 LO:21.86);ALT=G[chr15:45954151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	45981416	+	chr15	45983169	+	.	9	14	5942388_1	53.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5942388_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_45962001_45987001_72C;SPAN=1753;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:58 GQ:53.6 PL:[53.6, 0.0, 86.6] SR:14 DR:9 LR:-53.61 LO:54.05);ALT=G[chr15:45983169[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55485033	+	chr15	55489006	+	.	79	49	5956087_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=23;MATEID=5956087_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_55468001_55493001_269C;SPAN=3973;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:85 GQ:27 PL:[297.0, 27.0, 0.0] SR:49 DR:79 LR:-297.1 LO:297.1);ALT=T[chr15:55489006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34188507	+	chr15	55489006	+	.	40	26	5956092_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5956092_2;MATENM=4;NM=0;NUMPARTS=2;REPSEQ=CC;SCTG=c_15_55468001_55493001_269C;SECONDARY;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:40 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:26 DR:40 LR:-174.9 LO:174.9);ALT=]chr17:34188507]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr15	55562484	+	chr15	55581914	+	.	7	5	5956137_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=5956137_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_55566001_55591001_134C;SPAN=19430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:19 GQ:21.2 PL:[21.2, 0.0, 24.5] SR:5 DR:7 LR:-21.26 LO:21.28);ALT=T[chr15:55581914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55610067	+	chr15	55611129	+	.	0	10	5956693_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5956693_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_55590501_55615501_41C;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:10 DR:0 LR:-18.65 LO:22.38);ALT=T[chr15:55611129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55677914	+	chr15	55681562	+	.	0	8	5956345_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5956345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_55664001_55689001_98C;SPAN=3648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:8 DR:0 LR:-13.67 LO:17.51);ALT=T[chr15:55681562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	55677956	+	chr15	55700431	+	.	9	0	5956346_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5956346_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:55677956(+)-15:55700431(-)__15_55664001_55689001D;SPAN=22475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=C[chr15:55700431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59009928	+	chr15	59041677	+	.	0	8	5961685_1	17.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=5961685_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59020501_59045501_85C;SPAN=31749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:8 DR:0 LR:-17.2 LO:18.78);ALT=T[chr15:59041677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59186783	+	chr15	59189312	+	.	3	6	5961924_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5961924_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59167501_59192501_167C;SPAN=2529;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:6 DR:3 LR:-14.54 LO:19.45);ALT=T[chr15:59189312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59205898	+	chr15	59224553	+	GATAAAAGCATCATCTTCCACAGAAGCATCTCCACTCAACTCATCTGCTTCATGTTTTTT	0	28	5962091_1	82.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=GATAAAAGCATCATCTTCCACAGAAGCATCTCCACTCAACTCATCTGCTTCATGTTTTTT;MAPQ=60;MATEID=5962091_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_59216501_59241501_94C;SPAN=18655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:28 DR:0 LR:-82.52 LO:82.52);ALT=T[chr15:59224553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59931356	+	chr15	59934335	+	.	3	24	5963427_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5963427_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59927001_59952001_134C;SPAN=2979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:53 GQ:55.1 PL:[71.6, 0.0, 55.1] SR:24 DR:3 LR:-71.55 LO:71.55);ALT=T[chr15:59934335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59934462	+	chr15	59942867	+	.	0	19	5963438_1	46.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5963438_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59927001_59952001_18C;SPAN=8405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:59 GQ:46.7 PL:[46.7, 0.0, 96.2] SR:19 DR:0 LR:-46.73 LO:47.68);ALT=C[chr15:59942867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59934500	+	chr15	59949603	+	.	10	0	5963439_1	17.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=5963439_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:59934500(+)-15:59949603(-)__15_59927001_59952001D;SPAN=15103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:0 DR:10 LR:-17.03 LO:21.86);ALT=T[chr15:59949603[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59942975	+	chr15	59944405	+	.	0	80	5963453_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5963453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59927001_59952001_185C;SPAN=1430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:93 GQ:15 PL:[254.1, 15.0, 0.0] SR:80 DR:0 LR:-257.5 LO:257.5);ALT=G[chr15:59944405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59943023	+	chr15	59949602	+	.	56	0	5963454_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5963454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:59943023(+)-15:59949602(-)__15_59927001_59952001D;SPAN=6579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:61 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:0 DR:56 LR:-178.2 LO:178.2);ALT=A[chr15:59949602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59944527	+	chr15	59949604	+	.	74	7	5963460_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5963460_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59927001_59952001_89C;SPAN=5077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:66 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:7 DR:74 LR:-224.5 LO:224.5);ALT=T[chr15:59949604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59971968	+	chr15	59974607	+	AGGCTGGTCCTCTGGTCCAGTTATAGCTAGTATATCTGCTTCAATACTATCATCTTCTGGTAAAGGT	6	25	5963695_1	79.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AGGCTGGTCCTCTGGTCCAGTTATAGCTAGTATATCTGCTTCAATACTATCATCTTCTGGTAAAGGT;MAPQ=60;MATEID=5963695_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_59951501_59976501_156C;SPAN=2639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:61 GQ:66.2 PL:[79.4, 0.0, 66.2] SR:25 DR:6 LR:-79.24 LO:79.24);ALT=C[chr15:59974607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	59974714	+	chr15	59981333	+	.	0	20	5963707_1	62.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=5963707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_59951501_59976501_284C;SPAN=6619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:22 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:20 DR:0 LR:-62.72 LO:62.72);ALT=C[chr15:59981333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	62327252	+	chr15	62352473	+	AATTTGGCCAGCCTTGACTTTAAAAGGAACATCCAATTCACTCAGGGCATTTTCTTTTATCTGTAGATTATCTAAAGCCACATTT	3	14	5967075_1	40.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AATTTGGCCAGCCTTGACTTTAAAAGGAACATCCAATTCACTCAGGGCATTTTCTTTTATCTGTAGATTATCTAAAGCCACATTT;MAPQ=60;MATEID=5967075_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_15_62352501_62377501_224C;SPAN=25221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:21 GQ:7.7 PL:[40.7, 0.0, 7.7] SR:14 DR:3 LR:-41.52 LO:41.52);ALT=C[chr15:62352473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	62706095	+	chr15	62707793	+	.	73	50	5967651_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ATT;MAPQ=60;MATEID=5967651_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_62695501_62720501_151C;SPAN=1698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:19 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:50 DR:73 LR:-303.7 LO:303.7);ALT=T[chr15:62707793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63446261	+	chr15	63448610	+	TCTGTGAGTCTGGCCTTTCCTCCTGTAGGCTGGCACAACACTGTTGAACAACCTACACAAAGAACCACTGTCTGAGCATGGCTGAAAACCGTGGTGATCTTGTAGCA	6	390	5969019_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=TCTGTGAGTCTGGCCTTTCCTCCTGTAGGCTGGCACAACACTGTTGAACAACCTACACAAAGAACCACTGTCTGAGCATGGCTGAAAACCGTGGTGATCTTGTAGCA;MAPQ=60;MATEID=5969019_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_63430501_63455501_21C;SPAN=2349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:393 DP:99 GQ:99 PL:[1165.0, 106.1, 0.0] SR:390 DR:6 LR:-1165.0 LO:1165.0);ALT=T[chr15:63448610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63446261	+	chr15	63447819	+	.	0	186	5969018_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=5969018_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_63430501_63455501_21C;SPAN=1558;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:186 DP:106 GQ:50.2 PL:[551.2, 50.2, 0.0] SR:186 DR:0 LR:-551.2 LO:551.2);ALT=T[chr15:63447819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63446296	+	chr15	63449598	+	.	15	0	5969021_1	30.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=5969021_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:63446296(+)-15:63449598(-)__15_63430501_63455501D;SPAN=3302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:70 GQ:30.5 PL:[30.5, 0.0, 139.4] SR:0 DR:15 LR:-30.55 LO:34.51);ALT=A[chr15:63449598[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63447972	+	chr15	63449595	+	.	75	0	5969026_1	99.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=5969026_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:63447972(+)-15:63449595(-)__15_63430501_63455501D;SPAN=1623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:70 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:0 DR:75 LR:-221.2 LO:221.2);ALT=G[chr15:63449595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63569935	+	chr15	63571359	+	.	9	4	5969141_1	24.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5969141_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_15_63553001_63578001_27C;SPAN=1424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:4 DR:9 LR:-24.71 LO:27.71);ALT=G[chr15:63571359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	63797029	+	chr15	63824845	+	.	0	7	5969545_1	14.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5969545_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_63822501_63847501_88C;SPAN=27816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:31 GQ:14.9 PL:[14.9, 0.0, 57.8] SR:7 DR:0 LR:-14.71 LO:16.28);ALT=G[chr15:63824845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64067849	+	chr15	64126020	+	.	13	3	5970066_1	46.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5970066_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64116501_64141501_81C;SPAN=58171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:16 DP:16 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:3 DR:13 LR:-46.21 LO:46.21);ALT=C[chr15:64126020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64365227	+	chr15	64367691	+	.	3	5	5970673_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5970673_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64361501_64386501_231C;SPAN=2464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:5 DR:3 LR:-12.59 LO:17.19);ALT=A[chr15:64367691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64381051	+	chr15	64385852	+	ATAAACC	34	44	5970707_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=ATAAACC;MAPQ=60;MATEID=5970707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64361501_64386501_199C;SPAN=4801;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:63 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:44 DR:34 LR:-214.6 LO:214.6);ALT=C[chr15:64385852[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64388371	+	chr15	64404772	+	.	0	12	5970556_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5970556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64386001_64411001_99C;SPAN=16401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:12 DR:0 LR:-22.81 LO:27.0);ALT=C[chr15:64404772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64449110	+	chr15	64452302	+	.	8	45	5970803_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=5970803_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_15_64435001_64460001_159C;SPAN=3192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:70 GQ:23.9 PL:[146.0, 0.0, 23.9] SR:45 DR:8 LR:-151.1 LO:151.1);ALT=T[chr15:64452302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64449143	+	chr15	64455129	+	.	10	0	5970805_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5970805_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64449143(+)-15:64455129(-)__15_64435001_64460001D;SPAN=5986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:156 GQ:9.1 PL:[0.0, 9.1, 396.0] SR:0 DR:10 LR:9.254 LO:17.38);ALT=G[chr15:64455129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64452451	+	chr15	64455048	+	.	112	0	5970813_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5970813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64452451(+)-15:64455048(-)__15_64435001_64460001D;SPAN=2597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:84 GQ:30 PL:[330.0, 30.0, 0.0] SR:0 DR:112 LR:-330.1 LO:330.1);ALT=A[chr15:64455048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64658274	+	chr15	64668942	+	.	0	11	5971160_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=5971160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64655501_64680501_187C;SPAN=10668;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:11 DR:0 LR:-23.85 LO:25.91);ALT=T[chr15:64668942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64658276	+	chr15	64673157	+	.	0	13	5971161_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5971161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64655501_64680501_79C;SPAN=14881;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:69 GQ:24.2 PL:[24.2, 0.0, 143.0] SR:13 DR:0 LR:-24.22 LO:29.08);ALT=T[chr15:64673157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64658315	+	chr15	64673575	+	.	13	0	5971162_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5971162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64658315(+)-15:64673575(-)__15_64655501_64680501D;SPAN=15260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:84 GQ:20.3 PL:[20.3, 0.0, 182.0] SR:0 DR:13 LR:-20.16 LO:27.85);ALT=C[chr15:64673575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64669106	+	chr15	64673157	+	.	0	78	5971194_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5971194_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64655501_64680501_175C;SPAN=4051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:84 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:78 DR:0 LR:-247.6 LO:247.6);ALT=T[chr15:64673157[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64669154	+	chr15	64673556	+	.	86	0	5971195_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5971195_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:64669154(+)-15:64673556(-)__15_64655501_64680501D;SPAN=4402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:55 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:0 DR:86 LR:-254.2 LO:254.2);ALT=C[chr15:64673556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	64983793	+	chr15	64995228	+	.	0	8	5971813_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5971813_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_64974001_64999001_53C;SPAN=11435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:58 GQ:10.7 PL:[10.7, 0.0, 129.5] SR:8 DR:0 LR:-10.69 LO:16.71);ALT=G[chr15:64995228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65247389	+	chr15	65245582	+	.	15	0	5972637_1	41.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=5972637_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:65245582(-)-15:65247389(+)__15_65243501_65268501D;SPAN=1807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:30 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:0 DR:15 LR:-41.46 LO:41.46);ALT=]chr15:65247389]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	65257801	+	chr15	65261590	+	.	2	5	5972661_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=5972661_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_65243501_65268501_221C;SPAN=3789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:59 GQ:7.1 PL:[7.1, 0.0, 135.8] SR:5 DR:2 LR:-7.123 LO:14.13);ALT=C[chr15:65261590[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65273365	+	chr15	65282002	+	TTTTAAGGGGAACTGTACCTCTAAACCAGTTATAATCAGGAGAGACTTTAATCTCTCCCATGATTAGCTGAAATGGAGGTTAAT	25	62	5972695_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=TTTTAAGGGGAACTGTACCTCTAAACCAGTTATAATCAGGAGAGACTTTAATCTCTCCCATGATTAGCTGAAATGGAGGTTAAT;MAPQ=60;MATEID=5972695_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_65268001_65293001_135C;SPAN=8637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:64 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:62 DR:25 LR:-214.6 LO:214.6);ALT=T[chr15:65282002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65273365	+	chr15	65275845	+	.	2	27	5972694_1	80.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5972694_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_15_65268001_65293001_135C;SPAN=2480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:57 GQ:57.2 PL:[80.3, 0.0, 57.2] SR:27 DR:2 LR:-80.48 LO:80.48);ALT=T[chr15:65275845[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65275980	+	chr15	65282054	+	.	24	0	5972704_1	62.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5972704_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:65275980(+)-15:65282054(-)__15_65268001_65293001D;SPAN=6074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:62 GQ:62.6 PL:[62.6, 0.0, 85.7] SR:0 DR:24 LR:-62.43 LO:62.67);ALT=C[chr15:65282054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65412294	+	chr15	65421369	+	.	2	4	5972848_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5972848_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_65415001_65440001_61C;SPAN=9075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:25 GQ:13.1 PL:[13.1, 0.0, 46.1] SR:4 DR:2 LR:-13.03 LO:14.14);ALT=T[chr15:65421369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65804904	+	chr15	65809823	+	.	0	9	5973866_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5973866_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_65807001_65832001_258C;SPAN=4919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:9 DR:0 LR:-21.31 LO:22.09);ALT=T[chr15:65809823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	65823044	+	chr15	65847222	+	.	9	0	5973911_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5973911_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:65823044(+)-15:65847222(-)__15_65807001_65832001D;SPAN=24178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=G[chr15:65847222[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66161963	+	chr15	66169668	+	.	82	13	5974226_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5974226_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_66150001_66175001_191C;SPAN=7705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:68 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:13 DR:82 LR:-260.8 LO:260.8);ALT=G[chr15:66169668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66161987	+	chr15	66170095	+	.	16	0	5974227_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5974227_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:66161987(+)-15:66170095(-)__15_66150001_66175001D;SPAN=8108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:66 GQ:35 PL:[35.0, 0.0, 124.1] SR:0 DR:16 LR:-34.94 LO:37.79);ALT=C[chr15:66170095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66170293	+	chr15	66180036	+	AAAAGAATGGTTTGTCATTCATTGAAACTTCGGCCCTAGACTCTACAAATGTAGAAGCTGCTTTTCAGACAATTTTAA	2	22	5974237_1	69.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AAAAGAATGGTTTGTCATTCATTGAAACTTCGGCCCTAGACTCTACAAATGTAGAAGCTGCTTTTCAGACAATTTTAA;MAPQ=60;MATEID=5974237_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_66150001_66175001_258C;SPAN=9743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:24 GQ:6.3 PL:[69.3, 6.3, 0.0] SR:22 DR:2 LR:-69.32 LO:69.32);ALT=G[chr15:66180036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66172089	+	chr15	66180036	+	.	5	12	5974243_1	46.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=5974243_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_66150001_66175001_258C;SPAN=7947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:23 GQ:7.1 PL:[46.7, 0.0, 7.1] SR:12 DR:5 LR:-48.0 LO:48.0);ALT=G[chr15:66180036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	66786937	+	chr15	66789956	+	.	9	0	5975492_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5975492_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:66786937(+)-15:66789956(-)__15_66787001_66812001D;SPAN=3019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=T[chr15:66789956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	67529167	+	chr15	67546913	+	.	12	0	5976977_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5976977_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:67529167(+)-15:67546913(-)__15_67522001_67547001D;SPAN=17746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:0 DR:12 LR:-22.81 LO:27.0);ALT=A[chr15:67546913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	67811441	+	chr15	67813856	+	.	7	3	5977193_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5977193_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_67791501_67816501_98C;SPAN=2415;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:37 GQ:19.7 PL:[19.7, 0.0, 69.2] SR:3 DR:7 LR:-19.68 LO:21.27);ALT=C[chr15:67813856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	68346740	+	chr15	68378652	+	.	21	0	5978257_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5978257_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:68346740(+)-15:68378652(-)__15_68355001_68380001D;SPAN=31912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:56 GQ:54.2 PL:[54.2, 0.0, 80.6] SR:0 DR:21 LR:-54.15 LO:54.46);ALT=G[chr15:68378652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	68426020	+	chr15	68428928	+	.	56	40	5978453_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGAAATTTAGATTTTTA;MAPQ=60;MATEID=5978453_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_68404001_68429001_49C;SPAN=2908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:33 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:40 DR:56 LR:-237.7 LO:237.7);ALT=A[chr15:68428928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	68510992	+	chr15	68521839	+	.	0	8	5978358_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CCTGG;MAPQ=60;MATEID=5978358_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_68502001_68527001_148C;SPAN=10847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:8 DR:0 LR:-13.95 LO:17.59);ALT=G[chr15:68521839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69080263	+	chr15	69113048	+	.	52	0	5979461_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5979461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:69080263(+)-15:69113048(-)__15_69090001_69115001D;SPAN=32785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:37 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:0 DR:52 LR:-151.8 LO:151.8);ALT=A[chr15:69113048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	69745360	+	chr15	69747508	+	.	39	9	5980559_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=54;MATEID=5980559_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_69727001_69752001_96C;SPAN=2148;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:44 DP:911 GQ:99 PL:[0.0, 101.1, 2413.0] SR:9 DR:39 LR:101.6 LO:70.92);ALT=G[chr15:69747508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	70596153	+	chr15	70594649	+	.	39	0	5981768_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5981768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:70594649(-)-15:70596153(+)__15_70584501_70609501D;SPAN=1504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:69 GQ:57.2 PL:[110.0, 0.0, 57.2] SR:0 DR:39 LR:-110.9 LO:110.9);ALT=]chr15:70596153]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	71708609	+	chr15	71713691	+	ACC	69	42	5983513_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;INSERTION=ACC;MAPQ=60;MATEID=5983513_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_71711501_71736501_121C;SPAN=5082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:14 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:42 DR:69 LR:-267.4 LO:267.4);ALT=A[chr15:71713691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72029089	+	chr15	72027775	+	.	18	0	5984048_1	46.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=5984048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:72027775(-)-15:72029089(+)__15_72005501_72030501D;SPAN=1314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:49 GQ:46.1 PL:[46.1, 0.0, 72.5] SR:0 DR:18 LR:-46.14 LO:46.47);ALT=]chr15:72029089]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	72385978	+	chr15	72388159	+	.	43	32	5984719_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=GCCTGTAATCCCA;MAPQ=60;MATEID=5984719_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72373001_72398001_104C;SPAN=2181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:25 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:32 DR:43 LR:-191.4 LO:191.4);ALT=A[chr15:72388159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72492999	+	chr15	72494793	+	.	6	7	5984846_1	22.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=5984846_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72471001_72496001_272C;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:65 GQ:22.1 PL:[22.1, 0.0, 134.3] SR:7 DR:6 LR:-22.0 LO:26.73);ALT=G[chr15:72494793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72494962	+	chr15	72499069	+	.	8	15	5984886_1	59.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5984886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72495501_72520501_177C;SPAN=4107;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:35 GQ:23.6 PL:[59.9, 0.0, 23.6] SR:15 DR:8 LR:-60.61 LO:60.61);ALT=C[chr15:72499069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72499620	+	chr15	72500961	+	.	12	6	5984901_1	38.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=5984901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72495501_72520501_125C;SPAN=1341;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:64 GQ:38.9 PL:[38.9, 0.0, 114.8] SR:6 DR:12 LR:-38.78 LO:40.95);ALT=T[chr15:72500961[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72502200	+	chr15	72509750	+	GCCCTTGATGAGCCCAGTTCGGATCTCAGGTCCTTTAGTGTCTAGAGCCACAGCAACGGGCCGGTAGAGGATGGGGTCAGAAGCAAAGCTTTCCGTGGCTGTGCGCACATTCTTGATGGTCTCCGCATGGTA	0	49	5984906_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GCCCTTGATGAGCCCAGTTCGGATCTCAGGTCCTTTAGTGTCTAGAGCCACAGCAACGGGCCGGTAGAGGATGGGGTCAGAAGCAAAGCTTTCCGTGGCTGTGCGCACATTCTTGATGGTCTCCGCATGGTA;MAPQ=59;MATEID=5984906_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_72495501_72520501_169C;SPAN=7550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:58 GQ:5.7 PL:[151.8, 5.7, 0.0] SR:49 DR:0 LR:-156.5 LO:156.5);ALT=T[chr15:72509750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72502821	+	chr15	72509750	+	.	2	32	5984907_1	90.0	.	DISC_MAPQ=52;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=5984907_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_72495501_72520501_169C;SPAN=6929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:69 GQ:77 PL:[90.2, 0.0, 77.0] SR:32 DR:2 LR:-90.29 LO:90.29);ALT=T[chr15:72509750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72502856	+	chr15	72523455	+	.	11	0	5984949_1	29.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=5984949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:72502856(+)-15:72523455(-)__15_72520001_72545001D;SPAN=20599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:27 GQ:29 PL:[29.0, 0.0, 35.6] SR:0 DR:11 LR:-29.0 LO:29.04);ALT=A[chr15:72523455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72509842	+	chr15	72511284	+	.	0	95	5984920_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=5984920_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72495501_72520501_56C;SPAN=1442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:96 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:95 DR:0 LR:-283.9 LO:283.9);ALT=C[chr15:72511284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72509880	+	chr15	72523470	+	.	49	0	5984950_1	99.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=5984950_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:72509880(+)-15:72523470(-)__15_72520001_72545001D;SPAN=13590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:60 GQ:0.2 PL:[145.4, 0.0, 0.2] SR:0 DR:49 LR:-154.5 LO:154.5);ALT=T[chr15:72523470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72511453	+	chr15	72523456	+	.	163	30	5984951_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5984951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72520001_72545001_92C;SPAN=12003;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:180 DP:27 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:30 DR:163 LR:-534.7 LO:534.7);ALT=T[chr15:72523456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72636483	+	chr15	72637796	+	CAGCAAC	3	12	5985565_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CAGCAAC;MAPQ=60;MATEID=5985565_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72618001_72643001_64C;SPAN=1313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:77 GQ:25.4 PL:[25.4, 0.0, 160.7] SR:12 DR:3 LR:-25.35 LO:31.08);ALT=T[chr15:72637796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72641602	+	chr15	72642856	+	.	3	11	5985574_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCT;MAPQ=60;MATEID=5985574_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72618001_72643001_185C;SPAN=1254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:11 DR:3 LR:-26.66 LO:29.98);ALT=T[chr15:72642856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72641643	+	chr15	72643472	+	.	10	0	5985575_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5985575_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:72641643(+)-15:72643472(-)__15_72618001_72643001D;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:27 GQ:25.7 PL:[25.7, 0.0, 38.9] SR:0 DR:10 LR:-25.7 LO:25.86);ALT=A[chr15:72643472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	72648960	+	chr15	72668060	+	.	0	21	5985172_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=5985172_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_72667001_72692001_29C;SPAN=19100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:36 GQ:26.6 PL:[59.6, 0.0, 26.6] SR:21 DR:0 LR:-60.19 LO:60.19);ALT=T[chr15:72668060[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74287282	+	chr15	74290343	+	.	11	6	5987914_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=5987914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_74284001_74309001_174C;SPAN=3061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:73 GQ:33.2 PL:[33.2, 0.0, 142.1] SR:6 DR:11 LR:-33.04 LO:36.98);ALT=G[chr15:74290343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74738571	+	chr15	74740819	+	.	0	14	5988784_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=5988784_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_74725001_74750001_19C;SPAN=2248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:68 GQ:27.8 PL:[27.8, 0.0, 136.7] SR:14 DR:0 LR:-27.79 LO:31.93);ALT=G[chr15:74740819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74749013	+	chr15	74751025	+	.	0	20	5988959_1	56.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=5988959_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_74749501_74774501_290C;SPAN=2012;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:36 GQ:29.9 PL:[56.3, 0.0, 29.9] SR:20 DR:0 LR:-56.66 LO:56.66);ALT=C[chr15:74751025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74749060	+	chr15	74753398	+	.	8	0	5988961_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5988961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:74749060(+)-15:74753398(-)__15_74749501_74774501D;SPAN=4338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:28 GQ:18.8 PL:[18.8, 0.0, 48.5] SR:0 DR:8 LR:-18.82 LO:19.57);ALT=A[chr15:74753398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74751238	+	chr15	74753377	+	.	36	5	5988963_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5988963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_74749501_74774501_206C;SPAN=2139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:64 GQ:48.8 PL:[104.9, 0.0, 48.8] SR:5 DR:36 LR:-105.8 LO:105.8);ALT=C[chr15:74753377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	74908289	+	chr15	74912347	+	.	11	0	5989020_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5989020_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:74908289(+)-15:74912347(-)__15_74896501_74921501D;SPAN=4058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:54 GQ:21.8 PL:[21.8, 0.0, 107.6] SR:0 DR:11 LR:-21.68 LO:25.03);ALT=G[chr15:74912347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75075061	+	chr15	75090572	+	.	23	15	5989306_1	64.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5989306_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GAGAGA;SCTG=c_15_75068001_75093001_263C;SPAN=15511;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:51 GQ:25.5 PL:[64.5, 0.0, 25.5] SR:15 DR:23 LR:-65.19 LO:65.19);ALT=G[chr15:75090572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75075061	+	chr15	75090953	+	CTCTAATGGTACCAAGTGACAGGTTGGCTTTACTGTGACTCGGGGACGCCAGAGCTCCTGAGAAGATGTCAGCAATA	10	46	5989307_1	99.0	.	DISC_MAPQ=50;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CTCTAATGGTACCAAGTGACAGGTTGGCTTTACTGTGACTCGGGGACGCCAGAGCTCCTGAGAAGATGTCAGCAATA;MAPQ=60;MATEID=5989307_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_75068001_75093001_263C;SPAN=15892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:46 DR:10 LR:-155.1 LO:155.1);ALT=G[chr15:75090953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75144531	+	chr15	75165539	+	GGGGTCGGCTGGGTTGGTTCCACTGATGGCTGGAGAACCGCTGGCTGTGAGGACCCAGGGAGTTGGGTGACAGGAACTGTTGTCGCTGCATTTGTCTCTGAGAAGGGGTTGAATTCCGCCAGGCCGCCCTGCGGGGCGTTGGTCAGCTGGGTCACAGAGGGAT	0	48	5989627_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=GGGGTCGGCTGGGTTGGTTCCACTGATGGCTGGAGAACCGCTGGCTGTGAGGACCCAGGGAGTTGGGTGACAGGAACTGTTGTCGCTGCATTTGTCTCTGAGAAGGGGTTGAATTCCGCCAGGCCGCCCTGCGGGGCGTTGGTCAGCTGGGTCACAGAGGGAT;MAPQ=60;MATEID=5989627_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_15_75141501_75166501_136C;SPAN=21008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:56 GQ:8.4 PL:[151.8, 8.4, 0.0] SR:48 DR:0 LR:-154.2 LO:154.2);ALT=G[chr15:75165539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75146511	+	chr15	75165601	+	.	28	0	5989632_1	76.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5989632_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75146511(+)-15:75165601(-)__15_75141501_75166501D;SPAN=19090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:60 GQ:69.5 PL:[76.1, 0.0, 69.5] SR:0 DR:28 LR:-76.19 LO:76.19);ALT=T[chr15:75165601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75147037	+	chr15	75165604	+	.	31	0	5989635_1	87.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5989635_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75147037(+)-15:75165604(-)__15_75141501_75166501D;SPAN=18567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:56 GQ:47.6 PL:[87.2, 0.0, 47.6] SR:0 DR:31 LR:-87.74 LO:87.74);ALT=G[chr15:75165604[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75182482	+	chr15	75183717	+	.	13	0	5989855_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5989855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75182482(+)-15:75183717(-)__15_75166001_75191001D;SPAN=1235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:71 GQ:23.9 PL:[23.9, 0.0, 146.0] SR:0 DR:13 LR:-23.68 LO:28.9);ALT=G[chr15:75183717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75197572	+	chr15	75198926	+	.	0	6	5989757_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=5989757_2;MATENM=3;NM=0;NUMPARTS=2;SCTG=c_15_75190501_75215501_252C;SPAN=1354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:55 GQ:5 PL:[5.0, 0.0, 127.1] SR:6 DR:0 LR:-4.905 LO:11.87);ALT=C[chr15:75198926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75197574	+	chr15	75198616	+	.	0	5	5989758_1	3.0	.	EVDNC=ASSMB;HOMSEQ=GACCT;MAPQ=60;MATEID=5989758_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_75190501_75215501_32C;SPAN=1042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:5 DR:0 LR:-3.23 LO:9.742);ALT=T[chr15:75198616[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75212784	+	chr15	75215989	+	.	3	177	5989994_1	99.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5989994_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_75215001_75240001_71C;SPAN=3205;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:180 DP:52 GQ:48.7 PL:[534.7, 48.7, 0.0] SR:177 DR:3 LR:-534.7 LO:534.7);ALT=C[chr15:75215989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75216113	+	chr15	75219106	+	.	5	63	5990002_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5990002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_75215001_75240001_252C;SPAN=2993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:68 DP:77 GQ:17.4 PL:[221.1, 17.4, 0.0] SR:63 DR:5 LR:-221.7 LO:221.7);ALT=T[chr15:75219106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75221619	+	chr15	75230314	+	.	131	0	5990015_1	99.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=5990015_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75221619(+)-15:75230314(-)__15_75215001_75240001D;SPAN=8695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:131 DP:119 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:0 DR:131 LR:-386.2 LO:386.2);ALT=T[chr15:75230314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75320794	+	chr15	75335781	+	.	2	3	5989891_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5989891_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GGG;SCTG=c_15_75313001_75338001_166C;SPAN=14987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:58 GQ:0.8 PL:[0.8, 0.0, 139.4] SR:3 DR:2 LR:-0.7914 LO:9.357);ALT=G[chr15:75335781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75335877	+	chr15	75340894	+	ATGTGGAAGAGCCGCTCTGACCCAGTTCTGCACATTGACCTGCGGAGGTGGGCAGACCTCCTGCTGGTGGCTCCTCTTGATGCCAACACTCTGGGGAAGGTGGCCAGTGGCATCTGTGACAACTTGCTT	4	11	5990066_1	30.0	.	DISC_MAPQ=56;EVDNC=TSI_G;INSERTION=ATGTGGAAGAGCCGCTCTGACCCAGTTCTGCACATTGACCTGCGGAGGTGGGCAGACCTCCTGCTGGTGGCTCCTCTTGATGCCAACACTCTGGGGAAGGTGGCCAGTGGCATCTGTGACAACTTGCTT;MAPQ=60;MATEID=5990066_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_75337501_75362501_176C;SPAN=5017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:11 DR:4 LR:-30.67 LO:30.91);ALT=G[chr15:75340894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75624710	+	chr15	78240417	-	.	23	0	5995616_1	66.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=5995616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75624710(+)-15:78240417(+)__15_78228501_78253501D;SPAN=2615707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:15 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:23 LR:-66.02 LO:66.02);ALT=C]chr15:78240417];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr15	75628486	+	chr15	75631324	+	.	8	0	5991032_1	10.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=5991032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:75628486(+)-15:75631324(-)__15_75607001_75632001D;SPAN=2838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:0 DR:8 LR:-10.15 LO:16.58);ALT=G[chr15:75631324[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	75909893	+	chr15	75913235	+	.	2	11	5991502_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5991502_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_75901001_75926001_145C;SPAN=3342;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:59 GQ:20.3 PL:[20.3, 0.0, 122.6] SR:11 DR:2 LR:-20.33 LO:24.55);ALT=G[chr15:75913235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76028206	+	chr15	78161176	-	.	12	0	5995362_1	32.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=5995362_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:76028206(+)-15:78161176(+)__15_78155001_78180001D;SPAN=2132970;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:27 GQ:32.3 PL:[32.3, 0.0, 32.3] SR:0 DR:12 LR:-32.3 LO:32.3);ALT=T]chr15:78161176];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr15	76028395	-	chr15	78161017	+	.	10	0	5995363_1	27.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=5995363_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:76028395(-)-15:78161017(-)__15_78155001_78180001D;SPAN=2132622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:22 GQ:23.9 PL:[27.2, 0.0, 23.9] SR:0 DR:10 LR:-27.05 LO:27.05);ALT=[chr15:78161017[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	76235995	+	chr15	76248271	+	.	0	24	5992209_1	71.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=5992209_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76244001_76269001_261C;SPAN=12276;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:31 GQ:1.7 PL:[71.0, 0.0, 1.7] SR:24 DR:0 LR:-74.32 LO:74.32);ALT=C[chr15:76248271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76248355	+	chr15	76254168	+	.	0	19	5992218_1	47.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=5992218_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76244001_76269001_250C;SPAN=5813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:56 GQ:47.6 PL:[47.6, 0.0, 87.2] SR:19 DR:0 LR:-47.55 LO:48.22);ALT=G[chr15:76254168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76301636	+	chr15	76303562	+	.	0	30	5992264_1	83.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=5992264_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76293001_76318001_214C;SPAN=1926;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:58 GQ:56.9 PL:[83.3, 0.0, 56.9] SR:30 DR:0 LR:-83.57 LO:83.57);ALT=T[chr15:76303562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76301683	+	chr15	76304363	+	.	19	0	5992266_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5992266_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:76301683(+)-15:76304363(-)__15_76293001_76318001D;SPAN=2680;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:46 GQ:50.3 PL:[50.3, 0.0, 60.2] SR:0 DR:19 LR:-50.26 LO:50.32);ALT=C[chr15:76304363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76303629	+	chr15	76344405	+	.	0	7	5992395_1	16.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=5992395_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76342001_76367001_52C;SPAN=40776;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:26 GQ:16.1 PL:[16.1, 0.0, 45.8] SR:7 DR:0 LR:-16.06 LO:16.91);ALT=T[chr15:76344405[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76344569	+	chr15	76349293	+	.	20	0	5992406_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=5992406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:76344569(+)-15:76349293(-)__15_76342001_76367001D;SPAN=4724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:53 GQ:51.8 PL:[51.8, 0.0, 74.9] SR:0 DR:20 LR:-51.66 LO:51.93);ALT=A[chr15:76349293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76578825	+	chr15	76584772	+	CATAAATAGTTCTCACAAATGTGTCAGGTGACTTGATTGCAATGATGTCAGAAATCGGGGCAACCTCAAGTTTGGCTGCTACTCTGGGCAAAAGGTT	2	32	5992796_1	93.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CATAAATAGTTCTCACAAATGTGTCAGGTGACTTGATTGCAATGATGTCAGAAATCGGGGCAACCTCAAGTTTGGCTGCTACTCTGGGCAAAAGGTT;MAPQ=60;MATEID=5992796_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_76562501_76587501_234C;SPAN=5947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:56 GQ:41 PL:[93.8, 0.0, 41.0] SR:32 DR:2 LR:-94.82 LO:94.82);ALT=G[chr15:76584772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76578825	+	chr15	76580186	+	.	0	11	5992795_1	21.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=5992795_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_76562501_76587501_234C;SPAN=1361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:11 DR:0 LR:-21.14 LO:24.83);ALT=G[chr15:76580186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76580327	+	chr15	76603686	+	.	16	0	5992865_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5992865_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:76580327(+)-15:76603686(-)__15_76587001_76612001D;SPAN=23359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:43 GQ:41.3 PL:[41.3, 0.0, 61.1] SR:0 DR:16 LR:-41.17 LO:41.42);ALT=T[chr15:76603686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76585042	+	chr15	76603688	+	.	46	2	5992866_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=5992866_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_76587001_76612001_276C;SPAN=18646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:44 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:2 DR:46 LR:-138.6 LO:138.6);ALT=C[chr15:76603688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	76588079	+	chr15	76603690	+	.	32	7	5992872_1	92.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=5992872_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_15_76587001_76612001_30C;SPAN=15611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:73 GQ:82.7 PL:[92.6, 0.0, 82.7] SR:7 DR:32 LR:-92.47 LO:92.47);ALT=C[chr15:76603690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	77287950	+	chr15	77310488	+	.	0	8	5994016_1	20.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5994016_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_77297501_77322501_295C;SPAN=22538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:8 DR:0 LR:-19.91 LO:20.23);ALT=G[chr15:77310488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	77328276	+	chr15	77329383	+	.	2	4	5993989_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=5993989_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_77322001_77347001_134C;SPAN=1107;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:43 GQ:8.3 PL:[8.3, 0.0, 94.1] SR:4 DR:2 LR:-8.156 LO:12.56);ALT=G[chr15:77329383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	77348598	+	chr15	77363233	+	.	23	15	5994059_1	61.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=5994059_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AGAAGA;SCTG=c_15_77346501_77371501_171C;SPAN=14635;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:43 GQ:14.6 PL:[61.4, 0.0, 14.6] SR:15 DR:23 LR:-62.93 LO:62.93);ALT=C[chr15:77363233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78241309	-	chr15	79039378	+	.	16	0	5995641_1	41.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=5995641_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78241309(-)-15:79039378(-)__15_78228501_78253501D;SPAN=798069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:42 GQ:41.6 PL:[41.6, 0.0, 58.1] SR:0 DR:16 LR:-41.44 LO:41.63);ALT=[chr15:79039378[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	78346531	+	chr15	78369634	+	.	6	6	5995838_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=5995838_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78351001_78376001_16C;SPAN=23103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:27 GQ:19.1 PL:[19.1, 0.0, 45.5] SR:6 DR:6 LR:-19.09 LO:19.72);ALT=T[chr15:78369634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78441817	+	chr15	78452433	+	.	12	0	5995944_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5995944_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78441817(+)-15:78452433(-)__15_78449001_78474001D;SPAN=10616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:32 GQ:31.1 PL:[31.1, 0.0, 44.3] SR:0 DR:12 LR:-30.94 LO:31.12);ALT=G[chr15:78452433[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78456122	+	chr15	78457331	+	.	0	4	5995960_1	0	.	EVDNC=ASSMB;HOMSEQ=TAG;MAPQ=60;MATEID=5995960_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78449001_78474001_98C;SPAN=1209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:56 GQ:1.8 PL:[0.0, 1.8, 138.6] SR:4 DR:0 LR:1.968 LO:7.145);ALT=G[chr15:78457331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78575866	+	chr15	78577601	+	.	0	9	5996071_1	15.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=5996071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78571501_78596501_144C;SPAN=1735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:9 DR:0 LR:-15.35 LO:19.68);ALT=G[chr15:78577601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78585189	+	chr15	78591903	+	.	23	0	5996093_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5996093_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78585189(+)-15:78591903(-)__15_78571501_78596501D;SPAN=6714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:66 GQ:58.1 PL:[58.1, 0.0, 101.0] SR:0 DR:23 LR:-58.04 LO:58.71);ALT=T[chr15:78591903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78585673	+	chr15	78591902	+	.	43	0	5996096_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5996096_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78585673(+)-15:78591902(-)__15_78571501_78596501D;SPAN=6229;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:70 GQ:47 PL:[122.9, 0.0, 47.0] SR:0 DR:43 LR:-124.8 LO:124.8);ALT=G[chr15:78591902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78730699	+	chr15	78732134	+	.	3	3	5996521_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=5996521_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78718501_78743501_198C;SPAN=1435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:57 GQ:4.4 PL:[4.4, 0.0, 133.1] SR:3 DR:3 LR:-4.363 LO:11.78);ALT=G[chr15:78732134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78730739	+	chr15	78755262	+	.	11	0	5996522_1	27.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5996522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78730739(+)-15:78755262(-)__15_78718501_78743501D;SPAN=24523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:33 GQ:27.5 PL:[27.5, 0.0, 50.6] SR:0 DR:11 LR:-27.37 LO:27.81);ALT=C[chr15:78755262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78832882	+	chr15	78834518	+	AACTATATAAAGTTCAGAAAACAT	22	45	5996828_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AACTATATAAAGTTCAGAAAACAT;MAPQ=60;MATEID=5996828_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78816501_78841501_207C;SPAN=1636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:86 GQ:79.1 PL:[128.6, 0.0, 79.1] SR:45 DR:22 LR:-129.1 LO:129.1);ALT=G[chr15:78834518[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78832908	+	chr15	78834820	+	.	118	0	5996829_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5996829_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:78832908(+)-15:78834820(-)__15_78816501_78841501D;SPAN=1912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:85 GQ:31.8 PL:[349.8, 31.8, 0.0] SR:0 DR:118 LR:-349.9 LO:349.9);ALT=C[chr15:78834820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78834988	+	chr15	78836532	+	.	7	28	5996833_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=5996833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_78816501_78841501_273C;SPAN=1544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:65 GQ:58.4 PL:[98.0, 0.0, 58.4] SR:28 DR:7 LR:-98.42 LO:98.42);ALT=G[chr15:78836532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78836613	+	chr15	78837974	+	TTATTACAGTATCAGGAGCCAATACCTTGTGAGCAGTTGGTTACAGCGCTGTGTGATATCAAACAAGCTTATACACAATTTGG	5	42	5996840_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TTATTACAGTATCAGGAGCCAATACCTTGTGAGCAGTTGGTTACAGCGCTGTGTGATATCAAACAAGCTTATACACAATTTGG;MAPQ=60;MATEID=5996840_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_78816501_78841501_83C;SPAN=1361;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:64 GQ:22.4 PL:[131.3, 0.0, 22.4] SR:42 DR:5 LR:-135.4 LO:135.4);ALT=T[chr15:78837974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78838107	+	chr15	78841130	+	CAGCTGTGTCAATGTTGAAACAAGACTATAAAGAAGGAGAAATGACCTTGAAGTCAGCACTTGCTTTAGCTATCAAAGTACTAAATAAGACCATGGATGTTAGTAAACTCTCTGCTGAAAA	4	112	5996905_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAGCTGTGTCAATGTTGAAACAAGACTATAAAGAAGGAGAAATGACCTTGAAGTCAGCACTTGCTTTAGCTATCAAAGTACTAAATAAGACCATGGATGTTAGTAAACTCTCTGCTGAAAA;MAPQ=60;MATEID=5996905_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_78841001_78866001_140C;SPAN=3023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:35 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:112 DR:4 LR:-340.0 LO:340.0);ALT=G[chr15:78841130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78839040	+	chr15	78841130	+	.	3	53	5996906_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=5996906_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_15_78841001_78866001_140C;SPAN=2090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:35 GQ:15 PL:[165.0, 15.0, 0.0] SR:53 DR:3 LR:-165.0 LO:165.0);ALT=G[chr15:78841130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	78892128	+	chr22	31416873	+	.	10	26	7265638_1	98.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAATCCTAGCACTTTGGGAGGCCAAGGC;MAPQ=60;MATEID=7265638_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_31409001_31434001_100C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:49 GQ:19.7 PL:[98.9, 0.0, 19.7] SR:26 DR:10 LR:-101.9 LO:101.9);ALT=C[chr22:31416873[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr15	79229767	+	chr15	79237233	+	TAGACATCCATGACTTGAAGTGAAACTTCT	0	20	5997950_1	62.0	.	EVDNC=ASSMB;INSERTION=TAGACATCCATGACTTGAAGTGAAACTTCT;MAPQ=60;MATEID=5997950_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_15_79233001_79258001_248C;SPAN=7466;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:22 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:20 DR:0 LR:-62.72 LO:62.72);ALT=T[chr15:79237233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	79603761	+	chr15	79606096	+	.	0	28	5998307_1	74.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=5998307_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_79600501_79625501_42C;SPAN=2335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:68 GQ:74 PL:[74.0, 0.0, 90.5] SR:28 DR:0 LR:-74.01 LO:74.1);ALT=T[chr15:79606096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80181726	+	chr15	80189281	+	.	14	0	5999227_1	39.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=5999227_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:80181726(+)-15:80189281(-)__15_80188501_80213501D;SPAN=7555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:26 GQ:22.7 PL:[39.2, 0.0, 22.7] SR:0 DR:14 LR:-39.37 LO:39.37);ALT=T[chr15:80189281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80253517	+	chr15	80263041	+	.	3	6	5999419_1	18.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=5999419_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_80237501_80262501_89C;SPAN=9524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:30 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:6 DR:3 LR:-18.28 LO:19.28);ALT=C[chr15:80263041[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80445457	+	chr15	80452095	+	.	17	0	5999900_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5999900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:80445457(+)-15:80452095(-)__15_80433501_80458501D;SPAN=6638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:75 GQ:35.9 PL:[35.9, 0.0, 144.8] SR:0 DR:17 LR:-35.8 LO:39.58);ALT=G[chr15:80452095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80445477	+	chr15	80450402	+	.	28	19	5999901_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=5999901_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_80433501_80458501_213C;SPAN=4925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:73 GQ:86 PL:[89.3, 0.0, 86.0] SR:19 DR:28 LR:-89.16 LO:89.16);ALT=C[chr15:80450402[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80450512	+	chr15	80452096	+	.	0	21	5999909_1	51.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=5999909_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_80433501_80458501_276C;SPAN=1584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:66 GQ:51.5 PL:[51.5, 0.0, 107.6] SR:21 DR:0 LR:-51.44 LO:52.57);ALT=G[chr15:80452096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	80473502	+	chr15	80478469	+	.	0	32	5999855_1	86.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=5999855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_80458001_80483001_48C;SPAN=4967;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:70 GQ:83.3 PL:[86.6, 0.0, 83.3] SR:32 DR:0 LR:-86.67 LO:86.67);ALT=G[chr15:80478469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	81271820	+	chr15	81274289	+	.	0	11	6001017_1	20.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6001017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_81266501_81291501_50C;SPAN=2469;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:11 DR:0 LR:-20.87 LO:24.74);ALT=T[chr15:81274289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	81274567	+	chr15	81282081	+	.	9	0	6001025_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6001025_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:81274567(+)-15:81282081(-)__15_81266501_81291501D;SPAN=7514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=T[chr15:81282081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	81589471	+	chr15	81591730	+	.	10	0	6001642_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6001642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:81589471(+)-15:81591730(-)__15_81585001_81610001D;SPAN=2259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:0 DR:10 LR:-17.84 LO:22.11);ALT=C[chr15:81591730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83419602	+	chr15	83423379	+	.	14	13	6004856_1	57.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6004856_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_83398001_83423001_161C;SPAN=3777;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:33 GQ:20.9 PL:[57.2, 0.0, 20.9] SR:13 DR:14 LR:-57.87 LO:57.87);ALT=T[chr15:83423379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83423539	+	chr15	83425652	+	GGGAGGCCACAGCTTATGTGAATGACTTTCTCAGGAGTTATAAAGTGAT	0	13	6004660_1	30.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACAG;INSERTION=GGGAGGCCACAGCTTATGTGAATGACTTTCTCAGGAGTTATAAAGTGAT;MAPQ=60;MATEID=6004660_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_83422501_83447501_232C;SPAN=2113;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:46 GQ:30.5 PL:[30.5, 0.0, 80.0] SR:13 DR:0 LR:-30.45 LO:31.73);ALT=G[chr15:83425652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83551631	+	chr15	83557671	+	.	72	41	6005337_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACCAGCCACT;MAPQ=60;MATEID=6005337_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_15_83545001_83570001_155C;SPAN=6040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:33 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:41 DR:72 LR:-267.4 LO:267.4);ALT=T[chr15:83557671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83677430	+	chr15	83678989	+	.	0	12	6005077_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6005077_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_83667501_83692501_283C;SPAN=1559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:12 DR:0 LR:-27.42 LO:28.93);ALT=G[chr15:83678989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	83679117	+	chr15	83680248	+	.	27	13	6005084_1	86.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6005084_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_83667501_83692501_295C;SPAN=1131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:61 GQ:59.6 PL:[86.0, 0.0, 59.6] SR:13 DR:27 LR:-86.0 LO:86.0);ALT=T[chr15:83680248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85144366	+	chr15	85147049	+	.	17	2	6009234_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6009234_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_85137501_85162501_389C;SPAN=2683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:105 GQ:27.8 PL:[27.8, 0.0, 225.8] SR:2 DR:17 LR:-27.67 LO:36.79);ALT=G[chr15:85147049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85198643	+	chr15	85201225	+	GATTTGGGGTGCGGGGCGGCTGAGGCTCACGCCCAGAGCCTTCTTTAGCAGGAGGATTCCGAGCAGATCATGACTCAGCTGCAGTCGCTGGTCCCTCAGGGAGGTGTGGGGAGCTGTCCCCAATGGGGATGGGCTGGAAGGCTCCAGACTCTTCTTGCCCATGAAGTG	0	20	6008710_1	32.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=GATTTGGGGTGCGGGGCGGCTGAGGCTCACGCCCAGAGCCTTCTTTAGCAGGAGGATTCCGAGCAGATCATGACTCAGCTGCAGTCGCTGGTCCCTCAGGGAGGTGTGGGGAGCTGTCCCCAATGGGGATGGGCTGGAAGGCTCCAGACTCTTCTTGCCCATGAAGTG;MAPQ=60;MATEID=6008710_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_85186501_85211501_223C;SPAN=2582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:123 GQ:32.9 PL:[32.9, 0.0, 263.9] SR:20 DR:0 LR:-32.7 LO:43.32);ALT=G[chr15:85201225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85231035	+	chr15	85259255	+	.	77	0	6008921_1	99.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6008921_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:85231035(+)-15:85259255(-)__15_85235501_85260501D;SPAN=28220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:54 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:0 DR:77 LR:-227.8 LO:227.8);ALT=A[chr15:85259255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85234879	+	chr15	85259256	+	.	92	30	6008899_1	99.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=CTGC;MAPQ=60;MATEID=6008899_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_85211001_85236001_210C;SPAN=24377;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:64 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:30 DR:92 LR:-287.2 LO:287.2);ALT=C[chr15:85259256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	85291897	+	chr15	85307936	+	.	2	2	6009436_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6009436_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_85284501_85309501_271C;SPAN=16039;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:58 GQ:2.4 PL:[0.0, 2.4, 145.2] SR:2 DR:2 LR:2.51 LO:7.082);ALT=T[chr15:85307936[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	86057011	+	chr15	86059199	+	.	0	29	6012474_1	76.0	.	EVDNC=ASSMB;HOMSEQ=TTTT;MAPQ=60;MATEID=6012474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_86044001_86069001_291C;SPAN=2188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:70 GQ:76.7 PL:[76.7, 0.0, 93.2] SR:29 DR:0 LR:-76.76 LO:76.85);ALT=T[chr15:86059199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89009007	+	chr15	89010381	+	.	0	8	6022243_1	0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6022243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_89008501_89033501_83C;SPAN=1374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:8 DR:0 LR:6.374 LO:14.01);ALT=G[chr15:89010381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89011027	+	chr15	89015854	+	.	18	0	6022249_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6022249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:89011027(+)-15:89015854(-)__15_89008501_89033501D;SPAN=4827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:128 GQ:24.8 PL:[24.8, 0.0, 285.5] SR:0 DR:18 LR:-24.74 LO:37.75);ALT=G[chr15:89015854[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89011255	+	chr15	89015855	+	.	0	20	6022251_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6022251_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_89008501_89033501_163C;SPAN=4600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:131 GQ:30.8 PL:[30.8, 0.0, 284.9] SR:20 DR:0 LR:-30.53 LO:42.72);ALT=G[chr15:89015855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89015956	+	chr15	89018341	+	.	0	12	6022266_1	10.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6022266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_89008501_89033501_61C;SPAN=2385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:109 GQ:10.1 PL:[10.1, 0.0, 254.3] SR:12 DR:0 LR:-10.08 LO:23.8);ALT=A[chr15:89018341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89631800	+	chr15	89636861	+	.	10	0	6024444_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6024444_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:89631800(+)-15:89636861(-)__15_89621001_89646001D;SPAN=5061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:113 GQ:2.6 PL:[2.6, 0.0, 269.9] SR:0 DR:10 LR:-2.396 LO:18.83);ALT=G[chr15:89636861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89631824	+	chr15	89659551	+	.	8	0	6024510_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6024510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:89631824(+)-15:89659551(-)__15_89645501_89670501D;SPAN=27727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=A[chr15:89659551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	89745014	+	chr18	9914144	-	.	11	0	6538664_1	26.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=6538664_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:89745014(+)-18:9914144(+)__18_9898001_9923001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:35 GQ:26.9 PL:[26.9, 0.0, 56.6] SR:0 DR:11 LR:-26.83 LO:27.46);ALT=G]chr18:9914144];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr15	90628620	+	chr15	90630343	+	.	6	3	6028505_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6028505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90625501_90650501_399C;SPAN=1723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:3 DR:6 LR:2.902 LO:12.57);ALT=C[chr15:90630343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90631981	+	chr15	90633711	+	.	5	4	6028519_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6028519_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90625501_90650501_341C;SPAN=1730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:98 GQ:0 PL:[0.0, 0.0, 237.6] SR:4 DR:5 LR:0.1426 LO:14.77);ALT=T[chr15:90633711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90633923	+	chr15	90645507	+	.	24	0	6028530_1	50.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6028530_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:90633923(+)-15:90645507(-)__15_90625501_90650501D;SPAN=11584;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:106 GQ:50.6 PL:[50.6, 0.0, 205.7] SR:0 DR:24 LR:-50.51 LO:55.87);ALT=A[chr15:90645507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90634876	+	chr15	90645508	+	.	0	77	6028535_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6028535_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90625501_90650501_209C;SPAN=10632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:113 GQ:48.8 PL:[223.7, 0.0, 48.8] SR:77 DR:0 LR:-229.7 LO:229.7);ALT=T[chr15:90645508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90774928	+	chr15	90777080	+	.	71	0	6029401_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6029401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:90774928(+)-15:90777080(-)__15_90772501_90797501D;SPAN=2152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:117 GQ:80.6 PL:[202.7, 0.0, 80.6] SR:0 DR:71 LR:-205.5 LO:205.5);ALT=G[chr15:90777080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90775618	+	chr15	90777093	+	.	101	0	6029407_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6029407_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:90775618(+)-15:90777093(-)__15_90772501_90797501D;SPAN=1475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:101 DP:143 GQ:50.6 PL:[294.8, 0.0, 50.6] SR:0 DR:101 LR:-304.3 LO:304.3);ALT=T[chr15:90777093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	90931628	+	chr15	90934006	+	.	47	32	6030140_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6030140_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_90919501_90944501_281C;SPAN=2378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:115 GQ:94.4 PL:[183.5, 0.0, 94.4] SR:32 DR:47 LR:-184.9 LO:184.9);ALT=T[chr15:90934006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91383130	+	chr15	91384381	+	.	0	17	6031949_1	22.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6031949_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91360501_91385501_249C;SPAN=1251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:124 GQ:22.7 PL:[22.7, 0.0, 276.8] SR:17 DR:0 LR:-22.52 LO:35.45);ALT=G[chr15:91384381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91437289	+	chr15	91438645	+	.	0	6	6032052_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6032052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91434001_91459001_243C;SPAN=1356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:103 GQ:7.8 PL:[0.0, 7.8, 264.0] SR:6 DR:0 LR:8.099 LO:10.17);ALT=G[chr15:91438645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91459488	+	chr15	91461422	+	.	9	9	6032348_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6032348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91458501_91483501_83C;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:105 GQ:14.6 PL:[14.6, 0.0, 239.0] SR:9 DR:9 LR:-14.47 LO:26.49);ALT=T[chr15:91461422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91981580	+	chr15	91989266	+	.	49	34	6034063_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AAA;MAPQ=60;MATEID=6034063_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91973001_91998001_93C;SPAN=7686;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:94 GQ:27.5 PL:[199.1, 0.0, 27.5] SR:34 DR:49 LR:-206.3 LO:206.3);ALT=A[chr15:91989266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	91989617	+	chr15	91983461	+	A	35	27	6034067_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=6034067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_91973001_91998001_397C;SPAN=6156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:64 GQ:0.6 PL:[155.1, 0.6, 0.0] SR:27 DR:35 LR:-163.7 LO:163.7);ALT=]chr15:91989617]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	92674576	+	chr15	92677071	+	.	109	87	6036556_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6036556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_92659001_92684001_237C;SPAN=2495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:44 GQ:46 PL:[505.0, 46.0, 0.0] SR:87 DR:109 LR:-505.0 LO:505.0);ALT=T[chr15:92677071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93429484	+	chr15	93435234	+	.	2	3	6039476_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6039476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_93418501_93443501_152C;SPAN=5750;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:115 GQ:14.4 PL:[0.0, 14.4, 306.9] SR:3 DR:2 LR:14.65 LO:7.827);ALT=A[chr15:93435234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93431544	+	chr15	93435234	+	.	3	5	6039487_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6039487_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_93418501_93443501_178C;SPAN=3690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:120 GQ:12.6 PL:[0.0, 12.6, 316.8] SR:5 DR:3 LR:12.71 LO:9.763);ALT=T[chr15:93435234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93435332	+	chr15	93440986	+	.	9	0	6039499_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6039499_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:93435332(+)-15:93440986(-)__15_93418501_93443501D;SPAN=5654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:108 GQ:0.5 PL:[0.5, 0.0, 261.2] SR:0 DR:9 LR:-0.4492 LO:16.7);ALT=C[chr15:93440986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93470561	+	chr15	93480748	+	CAAGTAGCGGGTCTGAGAGTGGGAGCCCAAAAAGAAGAGGCCAGAGGCAGCTGAAAAAACA	0	13	6039558_1	11.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CAAGTAGCGGGTCTGAGAGTGGGAGCCCAAAAAGAAGAGGCCAGAGGCAGCTGAAAAAACA;MAPQ=60;MATEID=6039558_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_15_93467501_93492501_276C;SPAN=10187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:116 GQ:11.6 PL:[11.6, 0.0, 269.0] SR:13 DR:0 LR:-11.49 LO:25.89);ALT=G[chr15:93480748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	93480855	+	chr15	93482806	+	.	2	3	6039593_1	0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6039593_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_93467501_93492501_339C;SPAN=1951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:110 GQ:16.5 PL:[0.0, 16.5, 300.3] SR:3 DR:2 LR:16.6 LO:5.948);ALT=G[chr15:93482806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	94774894	+	chr15	94841428	+	.	11	2	6044324_1	20.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6044324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_94839501_94864501_18C;SPAN=66534;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:2 DR:11 LR:-20.87 LO:24.74);ALT=G[chr15:94841428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	94774894	+	chr15	94780957	+	.	27	7	6044155_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6044155_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_94766001_94791001_106C;SPAN=6063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:104 GQ:71 PL:[71.0, 0.0, 179.9] SR:7 DR:27 LR:-70.85 LO:73.54);ALT=G[chr15:94780957[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	99379574	-	chr15	99380633	+	.	8	0	6059188_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6059188_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:99379574(-)-15:99380633(-)__15_99372001_99397001D;SPAN=1059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:0 DR:8 LR:-0.9411 LO:14.92);ALT=[chr15:99380633[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	99587325	-	chr15	99588687	+	.	8	0	6060173_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6060173_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:99587325(-)-15:99588687(-)__15_99568001_99593001D;SPAN=1362;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:120 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.103 LO:14.04);ALT=[chr15:99588687[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	99791772	+	chr15	99796100	+	.	14	0	6060790_1	19.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6060790_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:99791772(+)-15:99796100(-)__15_99788501_99813501D;SPAN=4328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:98 GQ:19.7 PL:[19.7, 0.0, 217.7] SR:0 DR:14 LR:-19.66 LO:29.47);ALT=G[chr15:99796100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	100106294	+	chr15	100138633	+	.	8	0	6062123_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6062123_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100106294(+)-15:100138633(-)__15_100131501_100156501D;SPAN=32339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=C[chr15:100138633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	100106315	+	chr15	100173180	+	.	9	0	6062039_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6062039_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100106315(+)-15:100173180(-)__15_100156001_100181001D;SPAN=66865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=G[chr15:100173180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	100416715	+	chr15	100423235	+	.	40	0	6062961_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6062961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100416715(+)-15:100423235(-)__15_100401001_100426001D;SPAN=6520;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:63 GQ:35.9 PL:[115.1, 0.0, 35.9] SR:0 DR:40 LR:-117.1 LO:117.1);ALT=T[chr15:100423235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	101616225	+	chr15	100983925	+	.	13	0	6065013_1	31.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=6065013_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:100983925(-)-15:101616225(+)__15_100964501_100989501D;SPAN=632300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:43 GQ:31.4 PL:[31.4, 0.0, 71.0] SR:0 DR:13 LR:-31.26 LO:32.19);ALT=]chr15:101616225]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr15	101459683	+	chr15	101464734	+	.	11	0	6066601_1	17.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6066601_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:101459683(+)-15:101464734(-)__15_101454501_101479501D;SPAN=5051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:72 GQ:17 PL:[17.0, 0.0, 155.6] SR:0 DR:11 LR:-16.8 LO:23.5);ALT=C[chr15:101464734[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	101815567	+	chr15	101816746	+	.	0	10	6067833_1	3.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6067833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_101797501_101822501_237C;SPAN=1179;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:111 GQ:3.2 PL:[3.2, 0.0, 263.9] SR:10 DR:0 LR:-2.937 LO:18.91);ALT=C[chr15:101816746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	102187102	+	chr15	102190206	+	.	0	10	6069316_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6069316_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_102165001_102190001_219C;SPAN=3104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:10 DR:0 LR:-13.77 LO:20.98);ALT=C[chr15:102190206[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	102190355	+	chr15	102192473	+	.	9	0	6069098_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6069098_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:102190355(+)-15:102192473(-)__15_102189501_102214501D;SPAN=2118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:0 DR:9 LR:-0.7201 LO:16.74);ALT=T[chr15:102192473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	97560	+	chr16	101558	+	.	0	9	6071182_1	18.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6071182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_98001_123001_298C;SPAN=3998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:43 GQ:18.2 PL:[18.2, 0.0, 84.2] SR:9 DR:0 LR:-18.06 LO:20.6);ALT=G[chr16:101558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	97624	+	chr16	103501	+	.	11	0	6071183_1	21.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6071183_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:97624(+)-16:103501(-)__16_98001_123001D;SPAN=5877;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=G[chr16:103501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	101647	+	chr16	103474	+	.	0	8	6071201_1	4.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6071201_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_98001_123001_385C;SPAN=1827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:8 DR:0 LR:-4.192 LO:15.42);ALT=T[chr16:103474[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	104060	+	chr16	105457	+	.	31	31	6071216_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6071216_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_98001_123001_130C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:115 GQ:99 PL:[120.8, 0.0, 157.1] SR:31 DR:31 LR:-120.7 LO:121.0);ALT=T[chr16:105457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	128332	+	chr16	129421	+	.	135	13	6071097_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6071097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_122501_147501_174C;SPAN=1089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:69 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:13 DR:135 LR:-409.3 LO:409.3);ALT=G[chr16:129421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	129701	+	chr16	133047	+	.	0	7	6071101_1	3.0	.	EVDNC=ASSMB;HOMSEQ=ACAGGT;MAPQ=60;MATEID=6071101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_122501_147501_74C;SPAN=3346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:72 GQ:3.8 PL:[3.8, 0.0, 168.8] SR:7 DR:0 LR:-3.6 LO:13.48);ALT=T[chr16:133047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	243015	+	chr16	249061	+	.	3	5	6072036_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6072036_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_220501_245501_45C;SPAN=6046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:38 GQ:16.1 PL:[16.1, 0.0, 75.5] SR:5 DR:3 LR:-16.11 LO:18.33);ALT=C[chr16:249061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	284906	+	chr16	304376	+	.	9	0	6072835_1	18.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6072835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:284906(+)-16:304376(-)__16_269501_294501D;SPAN=19470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=C[chr16:304376[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	447314	+	chr16	448989	+	.	0	11	6072318_1	22.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6072318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_441001_466001_384C;SPAN=1675;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:11 DR:0 LR:-22.49 LO:25.34);ALT=G[chr16:448989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	620064	+	chr16	624063	+	.	11	0	6073042_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6073042_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:620064(+)-16:624063(-)__16_612501_637501D;SPAN=3999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:0 DR:11 LR:-19.51 LO:24.29);ALT=C[chr16:624063[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	684800	+	chr16	686093	+	.	0	13	6073516_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=6073516_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_661501_686501_313C;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:110 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:13 DR:0 LR:-13.11 LO:26.21);ALT=G[chr16:686093[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	789741	+	chr16	790930	+	.	11	0	6073745_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6073745_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:789741(+)-16:790930(-)__16_784001_809001D;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:0 DR:11 LR:-13.55 LO:22.7);ALT=A[chr16:790930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1359775	+	chr16	1364019	+	.	45	27	6075526_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6075526_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1347501_1372501_55C;SPAN=4244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:59 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:27 DR:45 LR:-174.9 LO:174.9);ALT=G[chr16:1364019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1359780	+	chr16	1364293	+	.	47	0	6075527_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6075527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1359780(+)-16:1364293(-)__16_1347501_1372501D;SPAN=4513;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:61 GQ:6.8 PL:[138.8, 0.0, 6.8] SR:0 DR:47 LR:-145.3 LO:145.3);ALT=C[chr16:1364293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1359783	+	chr16	1365653	+	.	17	0	6075528_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6075528_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1359783(+)-16:1365653(-)__16_1347501_1372501D;SPAN=5870;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.57 LO:43.16);ALT=G[chr16:1365653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1364098	+	chr16	1370175	+	GTTTCGTGGCTGTCCCAACAAAAAATCCCGATGGCACGATGAACCTCATGAACTGGGAGTGCGCCATTCCAGGAAAGAAAGGGACTCCGTGGGAAGGAGGCTTGTTTAAACTACGGATGCTTTTCAAAGATGATTATCCATCTTCGCCACCAAAAT	0	77	6075541_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GTAA;INSERTION=GTTTCGTGGCTGTCCCAACAAAAAATCCCGATGGCACGATGAACCTCATGAACTGGGAGTGCGCCATTCCAGGAAAGAAAGGGACTCCGTGGGAAGGAGGCTTGTTTAAACTACGGATGCTTTTCAAAGATGATTATCCATCTTCGCCACCAAAAT;MAPQ=60;MATEID=6075541_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_16_1347501_1372501_292C;SPAN=6077;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:79 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:77 DR:0 LR:-234.4 LO:234.4);ALT=G[chr16:1370175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1402047	+	chr16	1411742	+	.	40	0	6075659_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6075659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1402047(+)-16:1411742(-)__16_1396501_1421501D;SPAN=9695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:73 GQ:62.9 PL:[112.4, 0.0, 62.9] SR:0 DR:40 LR:-112.9 LO:112.9);ALT=G[chr16:1411742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1422869	+	chr16	1424141	+	.	35	0	6075579_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6075579_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1422869(+)-16:1424141(-)__16_1421001_1446001D;SPAN=1272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:58 GQ:40.4 PL:[99.8, 0.0, 40.4] SR:0 DR:35 LR:-101.2 LO:101.2);ALT=T[chr16:1424141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1790220	+	chr16	1788564	+	.	23	0	6076732_1	51.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=6076732_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1788564(-)-16:1790220(+)__16_1788501_1813501D;SPAN=1656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:92 GQ:51.2 PL:[51.2, 0.0, 170.0] SR:0 DR:23 LR:-51.0 LO:54.69);ALT=]chr16:1790220]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	1828616	+	chr16	1831359	+	.	10	38	6076853_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6076853_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1813001_1838001_253C;SPAN=2743;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:93 GQ:93.8 PL:[130.1, 0.0, 93.8] SR:38 DR:10 LR:-130.2 LO:130.2);ALT=G[chr16:1831359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1828661	+	chr16	1832500	+	.	53	0	6076854_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6076854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1828661(+)-16:1832500(-)__16_1813001_1838001D;SPAN=3839;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:75 GQ:26 PL:[154.7, 0.0, 26.0] SR:0 DR:53 LR:-159.7 LO:159.7);ALT=C[chr16:1832500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1831498	+	chr16	1832503	+	.	21	16	6076859_1	84.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6076859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1813001_1838001_234C;SPAN=1005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:89 GQ:84.8 PL:[84.8, 0.0, 131.0] SR:16 DR:21 LR:-84.82 LO:85.37);ALT=T[chr16:1832503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1833085	+	chr16	1836560	+	.	40	0	6076861_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6076861_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1833085(+)-16:1836560(-)__16_1813001_1838001D;SPAN=3475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:0 DR:40 LR:-109.9 LO:109.9);ALT=G[chr16:1836560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1833085	+	chr16	1837675	+	.	11	0	6077093_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6077093_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:1833085(+)-16:1837675(-)__16_1837501_1862501D;SPAN=4590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:40 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:0 DR:11 LR:-25.47 LO:26.69);ALT=G[chr16:1837675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1836656	+	chr16	1837676	+	.	0	5	6077094_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6077094_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1837501_1862501_23C;SPAN=1020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:40 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:5 DR:0 LR:-5.668 LO:10.21);ALT=G[chr16:1837676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1873039	+	chr16	1876711	+	.	17	4	6077037_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6077037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1862001_1887001_160C;SPAN=3672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:45 GQ:44 PL:[44.0, 0.0, 63.8] SR:4 DR:17 LR:-43.93 LO:44.15);ALT=C[chr16:1876711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1873040	+	chr16	1876506	+	.	3	2	6077038_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6077038_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1862001_1887001_350C;SPAN=3466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:52 GQ:2.6 PL:[2.6, 0.0, 121.4] SR:2 DR:3 LR:-2.417 LO:9.606);ALT=T[chr16:1876506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	1991407	+	chr16	1993102	+	.	10	3	6077323_1	18.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6077323_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_1984501_2009501_153C;SPAN=1695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:78 GQ:18.5 PL:[18.5, 0.0, 170.3] SR:3 DR:10 LR:-18.48 LO:25.68);ALT=C[chr16:1993102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2009755	+	chr16	2011152	+	.	74	122	6077699_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6077699_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2009001_2034001_286C;SPAN=1397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:168 DP:155 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:122 DR:74 LR:-498.4 LO:498.4);ALT=G[chr16:2011152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2083604	+	chr16	2086321	+	.	13	0	6077980_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6077980_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:2083604(+)-16:2086321(-)__16_2082501_2107501D;SPAN=2717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:67 GQ:24.8 PL:[24.8, 0.0, 137.0] SR:0 DR:13 LR:-24.76 LO:29.27);ALT=G[chr16:2086321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2090240	+	chr16	2093568	+	.	0	9	6078006_1	7.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6078006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2082501_2107501_65C;SPAN=3328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:9 DR:0 LR:-6.951 LO:17.74);ALT=C[chr16:2093568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2096371	+	chr16	2097710	+	.	23	5	6078027_1	58.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTGC;MAPQ=60;MATEID=6078027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_2082501_2107501_34C;SPAN=1339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:77 GQ:58.4 PL:[58.4, 0.0, 127.7] SR:5 DR:23 LR:-58.36 LO:59.81);ALT=C[chr16:2097710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2205860	+	chr16	2213883	+	.	7	4	6078222_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6078222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2205001_2230001_241C;SPAN=8023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:60 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:4 DR:7 LR:-13.45 LO:19.15);ALT=G[chr16:2213883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2205888	+	chr16	2215878	+	.	19	0	6078224_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6078224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:2205888(+)-16:2215878(-)__16_2205001_2230001D;SPAN=9990;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:109 GQ:33.2 PL:[33.2, 0.0, 231.2] SR:0 DR:19 LR:-33.19 LO:41.79);ALT=G[chr16:2215878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2214002	+	chr16	2218076	+	ACCAGAATGGAAACGACCTTCGGACCCGCCTTTTCAGCCGTCACCACCATCACAAA	0	25	6078247_1	66.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACCAGAATGGAAACGACCTTCGGACCCGCCTTTTCAGCCGTCACCACCATCACAAA;MAPQ=60;MATEID=6078247_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_2205001_2230001_323C;SPAN=4074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:59 GQ:66.5 PL:[66.5, 0.0, 76.4] SR:25 DR:0 LR:-66.54 LO:66.58);ALT=G[chr16:2218076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2290148	+	chr16	2293047	+	.	0	11	6078605_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6078605_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2278501_2303501_346C;SPAN=2899;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:11 DR:0 LR:-8.677 LO:21.71);ALT=T[chr16:2293047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2296989	+	chr16	2301316	+	.	0	11	6078629_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6078629_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2278501_2303501_69C;SPAN=4327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:11 DR:0 LR:-15.72 LO:23.22);ALT=T[chr16:2301316[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2564183	+	chr16	2569218	+	.	84	185	6080032_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6080032_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2548001_2573001_120C;SPAN=5035;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:233 DP:187 GQ:62.8 PL:[689.8, 62.8, 0.0] SR:185 DR:84 LR:-689.9 LO:689.9);ALT=G[chr16:2569218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2802849	+	chr16	2807472	+	.	0	19	6080817_1	35.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=6080817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2793001_2818001_158C;SPAN=4623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:103 GQ:35 PL:[35.0, 0.0, 213.2] SR:19 DR:0 LR:-34.81 LO:42.31);ALT=T[chr16:2807472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2802856	+	chr16	2806334	+	.	51	21	6080818_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6080818_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2793001_2818001_240C;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:127 GQ:99 PL:[153.8, 0.0, 153.8] SR:21 DR:51 LR:-153.8 LO:153.8);ALT=G[chr16:2806334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2822105	+	chr16	2826994	+	.	16	14	6080716_1	50.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6080716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2817501_2842501_363C;SPAN=4889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:169 GQ:50 PL:[50.0, 0.0, 360.2] SR:14 DR:16 LR:-49.94 LO:63.57);ALT=T[chr16:2826994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2825559	+	chr16	2826993	+	.	0	117	6080731_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6080731_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2817501_2842501_357C;SPAN=1434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:117 DP:168 GQ:66.8 PL:[340.7, 0.0, 66.8] SR:117 DR:0 LR:-351.1 LO:351.1);ALT=T[chr16:2826993[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2933368	+	chr16	2945220	+	.	13	6	6081385_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6081385_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_2940001_2965001_263C;SPAN=11852;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:49 GQ:39.5 PL:[39.5, 0.0, 79.1] SR:6 DR:13 LR:-39.54 LO:40.27);ALT=G[chr16:2945220[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2933387	+	chr16	2946350	+	.	18	0	6081386_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6081386_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:2933387(+)-16:2946350(-)__16_2940001_2965001D;SPAN=12963;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:36 GQ:36.5 PL:[49.7, 0.0, 36.5] SR:0 DR:18 LR:-49.75 LO:49.75);ALT=G[chr16:2946350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	2945322	+	chr16	2946351	+	.	0	14	6081411_1	24.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6081411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_2940001_2965001_147C;SPAN=1029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:81 GQ:24.5 PL:[24.5, 0.0, 169.7] SR:14 DR:0 LR:-24.27 LO:30.74);ALT=G[chr16:2946351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	3074366	+	chr16	3075706	+	.	0	6	6081643_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6081643_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_3062501_3087501_337C;SPAN=1340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:115 GQ:11.1 PL:[0.0, 11.1, 300.3] SR:6 DR:0 LR:11.35 LO:9.877);ALT=G[chr16:3075706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	3089322	+	chr20	62261478	+	.	5	22	7094979_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTTTGAGATGGAGTCTCG;MAPQ=60;MATEID=7094979_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62254501_62279501_392C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:50 GQ:59 PL:[62.3, 0.0, 59.0] SR:22 DR:5 LR:-62.38 LO:62.38);ALT=G[chr20:62261478[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr16	3554831	+	chr16	3556329	+	.	0	4	6083300_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6083300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_3552501_3577501_161C;SPAN=1498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:95 GQ:12.3 PL:[0.0, 12.3, 254.1] SR:4 DR:0 LR:12.53 LO:6.205);ALT=G[chr16:3556329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	3714462	+	chr16	3715971	+	.	2	3	6083900_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6083900_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_3699501_3724501_314C;SPAN=1509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:102 GQ:14.1 PL:[0.0, 14.1, 273.9] SR:3 DR:2 LR:14.43 LO:6.08);ALT=T[chr16:3715971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	3739139	+	chr16	3740826	+	.	0	9	6084006_1	5.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=6084006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_3724001_3749001_386C;SPAN=1687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:9 DR:0 LR:-5.326 LO:17.45);ALT=C[chr16:3740826[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	3740988	+	chr16	3767421	+	.	15	2	6084361_1	45.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6084361_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_3748501_3773501_288C;SPAN=26433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:28 GQ:22.1 PL:[45.2, 0.0, 22.1] SR:2 DR:15 LR:-45.63 LO:45.63);ALT=T[chr16:3767421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4209090	+	chr16	4210458	-	.	8	0	6086071_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6086071_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4209090(+)-16:4210458(+)__16_4189501_4214501D;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=G]chr16:4210458];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	4391643	+	chr16	4401230	+	.	48	0	6086527_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6086527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4391643(+)-16:4401230(-)__16_4385501_4410501D;SPAN=9587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:79 GQ:54.5 PL:[137.0, 0.0, 54.5] SR:0 DR:48 LR:-139.0 LO:139.0);ALT=C[chr16:4401230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4393338	+	chr16	4401231	+	.	13	0	6086531_1	18.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6086531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4393338(+)-16:4401231(-)__16_4385501_4410501D;SPAN=7893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:90 GQ:18.5 PL:[18.5, 0.0, 200.0] SR:0 DR:13 LR:-18.53 LO:27.43);ALT=C[chr16:4401231[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4463454	+	chr16	4466526	+	.	14	0	6086646_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6086646_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4463454(+)-16:4466526(-)__16_4459001_4484001D;SPAN=3072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:79 GQ:24.8 PL:[24.8, 0.0, 166.7] SR:0 DR:14 LR:-24.81 LO:30.91);ALT=T[chr16:4466526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4486744	-	chr16	4487906	+	.	8	0	6086748_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6086748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4486744(-)-16:4487906(-)__16_4483501_4508501D;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:102 GQ:0.9 PL:[0.0, 0.9, 247.5] SR:0 DR:8 LR:1.226 LO:14.63);ALT=[chr16:4487906[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	4511962	+	chr16	4513661	+	.	0	10	6087132_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6087132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_4508001_4533001_14C;SPAN=1699;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:10 DR:0 LR:-8.627 LO:19.88);ALT=T[chr16:4513661[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4519468	+	chr16	4524091	+	.	0	20	6087158_1	40.0	.	EVDNC=ASSMB;HOMSEQ=CACCT;MAPQ=60;MATEID=6087158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_4508001_4533001_309C;SPAN=4623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:96 GQ:40.1 PL:[40.1, 0.0, 191.9] SR:20 DR:0 LR:-40.01 LO:45.73);ALT=T[chr16:4524091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4519729	+	chr16	4524475	+	.	23	0	6087159_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6087159_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4519729(+)-16:4524475(-)__16_4508001_4533001D;SPAN=4746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:100 GQ:48.8 PL:[48.8, 0.0, 194.0] SR:0 DR:23 LR:-48.83 LO:53.72);ALT=G[chr16:4524475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4526527	+	chr16	4556893	+	.	9	0	6087193_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6087193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4526527(+)-16:4556893(-)__16_4508001_4533001D;SPAN=30366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:29 GQ:21.8 PL:[21.8, 0.0, 48.2] SR:0 DR:9 LR:-21.85 LO:22.41);ALT=C[chr16:4556893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4526532	+	chr16	4555480	+	.	18	0	6087194_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6087194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4526532(+)-16:4555480(-)__16_4508001_4533001D;SPAN=28948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:29 GQ:18.5 PL:[51.5, 0.0, 18.5] SR:0 DR:18 LR:-52.4 LO:52.4);ALT=T[chr16:4555480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4555611	+	chr16	4556894	+	.	0	18	6087015_1	32.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6087015_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_4532501_4557501_246C;SPAN=1283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:18 DR:0 LR:-32.87 LO:40.05);ALT=G[chr16:4556894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4564194	+	chr16	4588709	+	.	16	0	6087027_1	44.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6087027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4564194(+)-16:4588709(-)__16_4581501_4606501D;SPAN=24515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:29 GQ:25.1 PL:[44.9, 0.0, 25.1] SR:0 DR:16 LR:-45.25 LO:45.25);ALT=T[chr16:4588709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4675050	+	chr16	4700365	+	.	0	16	6087703_1	43.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6087703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_4679501_4704501_234C;SPAN=25315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:34 GQ:37.1 PL:[43.7, 0.0, 37.1] SR:16 DR:0 LR:-43.62 LO:43.62);ALT=G[chr16:4700365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	4769956	+	chr16	4772365	+	.	28	0	6087962_1	76.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6087962_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:4769956(+)-16:4772365(-)__16_4753001_4778001D;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:60 GQ:69.5 PL:[76.1, 0.0, 69.5] SR:0 DR:28 LR:-76.19 LO:76.19);ALT=A[chr16:4772365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	8715643	+	chr16	8719351	+	.	10	0	6100427_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6100427_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:8715643(+)-16:8719351(-)__16_8697501_8722501D;SPAN=3708;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:84 GQ:10.4 PL:[10.4, 0.0, 191.9] SR:0 DR:10 LR:-10.25 LO:20.2);ALT=G[chr16:8719351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	8953216	+	chr16	8962820	+	.	8	0	6101683_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6101683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:8953216(+)-16:8962820(-)__16_8942501_8967501D;SPAN=9604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=G[chr16:8962820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18797660	+	chr16	18799383	+	.	0	11	6138783_1	8.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6138783_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_109C;SPAN=1723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:104 GQ:8.3 PL:[8.3, 0.0, 242.6] SR:11 DR:0 LR:-8.135 LO:21.61);ALT=T[chr16:18799383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18800442	+	chr16	18801566	+	.	38	19	6138794_1	99.0	.	DISC_MAPQ=26;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=54;MATEID=6138794_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_144C;SPAN=1124;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:146 GQ:99 PL:[112.4, 0.0, 241.1] SR:19 DR:38 LR:-112.3 LO:114.9);ALT=T[chr16:18801566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18804694	+	chr16	18805921	+	.	2	30	6138809_1	83.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=28;MATEID=6138809_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_94C;SPAN=1227;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:83 GQ:83.3 PL:[83.3, 0.0, 116.3] SR:30 DR:2 LR:-83.15 LO:83.48);ALT=T[chr16:18805921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18809410	+	chr16	18812805	+	.	33	0	6138826_1	73.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6138826_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:18809410(+)-16:18812805(-)__16_18791501_18816501D;SPAN=3395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:132 GQ:73.4 PL:[73.4, 0.0, 245.0] SR:0 DR:33 LR:-73.17 LO:78.46);ALT=T[chr16:18812805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18810157	+	chr16	18812752	+	.	79	25	6138829_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6138829_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18791501_18816501_205C;SPAN=2595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:112 GQ:16.8 PL:[303.6, 16.8, 0.0] SR:25 DR:79 LR:-308.5 LO:308.5);ALT=C[chr16:18812752[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	18908280	+	chr16	18937272	+	.	2	2	6139742_1	4.0	.	DISC_MAPQ=13;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=48;MATEID=6139742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_18889501_18914501_456C;SPAN=28992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:33 GQ:4.4 PL:[4.4, 0.0, 73.7] SR:2 DR:2 LR:-4.264 LO:8.111);ALT=T[chr16:18937272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	19576274	+	chr16	19580746	+	.	6	3	6141770_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=6141770_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_19575501_19600501_194C;SPAN=4472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:3 DR:6 LR:-2.296 LO:15.12);ALT=T[chr16:19580746[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	19726348	+	chr16	19729478	+	.	13	0	6142199_1	18.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6142199_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:19726348(+)-16:19729478(-)__16_19722501_19747501D;SPAN=3130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:89 GQ:18.8 PL:[18.8, 0.0, 197.0] SR:0 DR:13 LR:-18.8 LO:27.5);ALT=T[chr16:19729478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	42458191	+	chr16	20202872	+	.	5	18	7183592_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAAAGAAAGAAAGAAAGAAAGAAAGAAA;MAPQ=60;MATEID=7183592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_42434001_42459001_8C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:22 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:18 DR:5 LR:-62.72 LO:62.72);ALT=]chr21:42458191]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	20911857	+	chr16	20926878	+	.	14	6	6146340_1	37.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=6146340_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_20923001_20948001_283C;SPAN=15021;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:56 GQ:37.7 PL:[37.7, 0.0, 97.1] SR:6 DR:14 LR:-37.64 LO:39.14);ALT=A[chr16:20926878[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	20912227	+	chr16	20926875	+	.	28	0	6146048_1	76.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6146048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:20912227(+)-16:20926875(-)__16_20898501_20923501D;SPAN=14648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:60 GQ:69.5 PL:[76.1, 0.0, 69.5] SR:0 DR:28 LR:-76.19 LO:76.19);ALT=G[chr16:20926875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	20927036	+	chr16	20931444	+	.	0	16	6146362_1	29.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6146362_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_20923001_20948001_132C;SPAN=4408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:87 GQ:29.3 PL:[29.3, 0.0, 181.1] SR:16 DR:0 LR:-29.25 LO:35.61);ALT=T[chr16:20931444[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	20931536	+	chr16	20935322	+	.	3	10	6146374_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6146374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_20923001_20948001_84C;SPAN=3786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:81 GQ:17.9 PL:[17.9, 0.0, 176.3] SR:10 DR:3 LR:-17.67 LO:25.46);ALT=A[chr16:20935322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21170099	+	chr16	21172295	+	.	38	0	6147051_1	98.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6147051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:21170099(+)-16:21172295(-)__16_21168001_21193001D;SPAN=2196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:101 GQ:98.3 PL:[98.3, 0.0, 144.5] SR:0 DR:38 LR:-98.08 LO:98.61);ALT=G[chr16:21172295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21594442	+	chr16	22710751	-	ATG	48	34	6154760_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;INSERTION=ATG;MAPQ=60;MATEID=6154760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_22687001_22712001_390C;SPAN=1116309;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:50 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:34 DR:48 LR:-204.7 LO:204.7);ALT=C]chr16:22710751];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	21611219	+	chr16	21623964	+	.	20	32	6149572_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6149572_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21609001_21634001_34C;SPAN=12745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:92 GQ:99 PL:[104.0, 0.0, 117.2] SR:32 DR:20 LR:-103.8 LO:103.9);ALT=G[chr16:21623964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21611221	+	chr16	21629183	+	.	2	2	6149573_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=6149573_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21609001_21634001_240C;SPAN=17962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:96 GQ:12.6 PL:[0.0, 12.6, 257.4] SR:2 DR:2 LR:12.8 LO:6.187);ALT=T[chr16:21629183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21624158	+	chr16	21629185	+	.	5	4	6149619_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6149619_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21609001_21634001_324C;SPAN=5027;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:4 DR:5 LR:2.581 LO:14.46);ALT=T[chr16:21629185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21629395	+	chr16	21636250	+	.	11	6	6149632_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6149632_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21609001_21634001_363C;SPAN=6855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:39 GQ:42.2 PL:[42.2, 0.0, 52.1] SR:6 DR:11 LR:-42.25 LO:42.31);ALT=G[chr16:21636250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21636438	+	chr16	21666550	+	.	6	6	6149684_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6149684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21658001_21683001_8C;SPAN=30112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:6 DR:6 LR:-20.01 LO:22.86);ALT=T[chr16:21666550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21658848	+	chr16	21663865	+	.	23	0	6149685_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6149685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:21658848(+)-16:21663865(-)__16_21658001_21683001D;SPAN=5017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:92 GQ:51.2 PL:[51.2, 0.0, 170.0] SR:0 DR:23 LR:-51.0 LO:54.69);ALT=C[chr16:21663865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29119271	+	chr16	21946770	+	GATCGCCTGTGTGCA	2	17	6177146_1	50.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=GATCGCCTGTGTGCA;MAPQ=60;MATEID=6177146_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_29106001_29131001_325C;SPAN=7172501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:47 GQ:50 PL:[50.0, 0.0, 63.2] SR:17 DR:2 LR:-49.99 LO:50.08);ALT=]chr16:29119271]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	21964777	+	chr16	21968555	+	.	63	15	6150819_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6150819_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21952001_21977001_384C;SPAN=3778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:77 DP:98 GQ:9.8 PL:[227.6, 0.0, 9.8] SR:15 DR:63 LR:-239.6 LO:239.6);ALT=G[chr16:21968555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21968887	+	chr16	21973779	+	ACGACAAAAGGAGCTTCATCTTTCAAGATAACCCGTGGAATTGAAGCAGTTGGTGGCAAATTA	4	25	6150842_1	57.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACGACAAAAGGAGCTTCATCTTTCAAGATAACCCGTGGAATTGAAGCAGTTGGTGGCAAATTA;MAPQ=60;MATEID=6150842_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_16_21952001_21977001_32C;SPAN=4892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:92 GQ:57.8 PL:[57.8, 0.0, 163.4] SR:25 DR:4 LR:-57.6 LO:60.51);ALT=G[chr16:21973779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21974206	+	chr16	21979947	+	ATGTCATTGAAAATTTGCATGCAGCAGCTTACCGGAATGCCTTGGCTAATCCCTTGTATTGTCCTGACTATAGGATTGGAAAAGTGACATCAGAGG	0	13	6150890_1	32.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATGTCATTGAAAATTTGCATGCAGCAGCTTACCGGAATGCCTTGGCTAATCCCTTGTATTGTCCTGACTATAGGATTGGAAAAGTGACATCAGAGG;MAPQ=60;MATEID=6150890_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_21976501_22001501_155C;SPAN=5741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:37 GQ:32.9 PL:[32.9, 0.0, 56.0] SR:13 DR:0 LR:-32.89 LO:33.24);ALT=C[chr16:21979947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	21992022	+	chr16	21994412	+	CA	0	31	6150942_1	68.0	.	EVDNC=ASSMB;INSERTION=CA;MAPQ=60;MATEID=6150942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_21976501_22001501_306C;SPAN=2390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:126 GQ:68.3 PL:[68.3, 0.0, 236.6] SR:31 DR:0 LR:-68.2 LO:73.45);ALT=G[chr16:21994412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23047775	+	chr16	23049532	+	GATTCT	50	32	6155842_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GATTCT;MAPQ=60;MATEID=6155842_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23030001_23055001_306C;SPAN=1757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:74 GQ:16.5 PL:[211.2, 16.5, 0.0] SR:32 DR:50 LR:-211.3 LO:211.3);ALT=A[chr16:23049532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23505700	+	chr16	23521644	+	CATTGGGGTCAGTGTTCACCTGCTCACAGAAATTCTGGATAGCTGACCAATCCTGTTCCGACATGCTTGGGTCTGTGGCTTTGTTC	0	8	6157381_1	13.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATTGGGGTCAGTGTTCACCTGCTCACAGAAATTCTGGATAGCTGACCAATCCTGTTCCGACATGCTTGGGTCTGTGGCTTTGTTC;MAPQ=60;MATEID=6157381_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_16_23495501_23520501_179C;SPAN=15944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:8 DR:0 LR:-13.67 LO:17.51);ALT=C[chr16:23521644[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23592497	+	chr16	23593597	+	.	0	53	6157980_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6157980_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23593501_23618501_319C;SPAN=1100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:48 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:53 DR:0 LR:-155.1 LO:155.1);ALT=G[chr16:23593597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23593697	+	chr16	23596656	+	.	3	24	6157981_1	66.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6157981_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23593501_23618501_260C;SPAN=2959;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:83 GQ:66.8 PL:[66.8, 0.0, 132.8] SR:24 DR:3 LR:-66.64 LO:67.91);ALT=C[chr16:23596656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23596746	+	chr16	23598518	+	.	0	20	6157990_1	39.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6157990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23593501_23618501_291C;SPAN=1772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:99 GQ:39.2 PL:[39.2, 0.0, 200.9] SR:20 DR:0 LR:-39.2 LO:45.43);ALT=T[chr16:23598518[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23596793	+	chr16	23607500	+	.	10	0	6157991_1	1.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6157991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:23596793(+)-16:23607500(-)__16_23593501_23618501D;SPAN=10707;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:118 GQ:1.1 PL:[1.1, 0.0, 284.9] SR:0 DR:10 LR:-1.041 LO:18.64);ALT=G[chr16:23607500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	23598642	+	chr16	23607442	+	.	69	90	6157996_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6157996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_23593501_23618501_192C;SPAN=8800;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:134 GQ:19.5 PL:[363.0, 19.5, 0.0] SR:90 DR:69 LR:-369.8 LO:369.8);ALT=T[chr16:23607442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66002029	+	chr16	24423750	+	.	14	0	6477044_1	35.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6477044_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:24423750(-)-17:66002029(+)__17_65978501_66003501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:40 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:0 DR:14 LR:-35.38 LO:35.77);ALT=]chr17:66002029]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr16	24517998	+	chr16	24519033	-	.	8	0	6161037_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6161037_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:24517998(+)-16:24519033(+)__16_24500001_24525001D;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-2.025 LO:15.08);ALT=G]chr16:24519033];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	24988686	+	chr16	25026591	+	.	9	0	6162924_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6162924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:24988686(+)-16:25026591(-)__16_25014501_25039501D;SPAN=37905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=T[chr16:25026591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	25137760	+	chr16	25066604	+	.	23	0	6163318_1	66.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6163318_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:25066604(-)-16:25137760(+)__16_25112501_25137501D;SPAN=71156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:0 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:23 LR:-66.02 LO:66.02);ALT=]chr16:25137760]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	25123319	+	chr16	25139794	+	.	0	14	6163336_1	36.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=6163336_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_25112501_25137501_277C;SPAN=16475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:35 GQ:36.8 PL:[36.8, 0.0, 46.7] SR:14 DR:0 LR:-36.73 LO:36.82);ALT=T[chr16:25139794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	25186356	+	chr16	25189321	+	.	2	15	6163592_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6163592_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_25186001_25211001_204C;SPAN=2965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:113 GQ:22.4 PL:[22.4, 0.0, 250.1] SR:15 DR:2 LR:-22.2 LO:33.61);ALT=G[chr16:25189321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	25340111	+	chr16	25343128	+	.	0	87	6164173_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6164173_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_25333001_25358001_263C;SPAN=3017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:39 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:87 DR:0 LR:-257.5 LO:257.5);ALT=G[chr16:25343128[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	28500708	+	chr16	28503034	+	AGAAGCCCACCGCGTTCTTCCAATGCGCGCCCTGATGGTCCAACAGAGGGAGCCGGGGCTCCGGGACGGTCTCCTCC	3	11	6174048_1	11.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=AGAAGCCCACCGCGTTCTTCCAATGCGCGCCCTGATGGTCCAACAGAGGGAGCCGGGGCTCCGGGACGGTCTCCTCC;MAPQ=60;MATEID=6174048_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_28493501_28518501_236C;SPAN=2326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:105 GQ:11.3 PL:[11.3, 0.0, 242.3] SR:11 DR:3 LR:-11.17 LO:24.01);ALT=C[chr16:28503034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	28565384	+	chr16	28596230	+	.	9	0	6174994_1	16.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6174994_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:28565384(+)-16:28596230(-)__16_28542501_28567501D;SPAN=30846;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=T[chr16:28596230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	28565420	+	chr16	28592375	+	.	8	10	6174995_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6174995_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_28542501_28567501_33C;SPAN=26955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:10 DR:8 LR:-25.25 LO:27.93);ALT=T[chr16:28592375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	28875273	+	chr16	28877328	+	.	9	0	6176557_1	1.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6176557_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:28875273(+)-16:28877328(-)__16_28861001_28886001D;SPAN=2055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:0 DR:9 LR:-1.262 LO:16.82);ALT=C[chr16:28877328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29309436	+	chr16	88305441	+	.	0	33	6273595_1	97.0	.	EVDNC=ASSMB;HOMSEQ=TGGGTAGATGGATGAATT;MAPQ=60;MATEID=6273595_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_16_88298001_88323001_87C;SPAN=58996005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:44 GQ:8 PL:[97.1, 0.0, 8.0] SR:33 DR:0 LR:-101.2 LO:101.2);ALT=T[chr16:88305441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29690584	+	chr16	29705982	+	.	14	0	6180496_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6180496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:29690584(+)-16:29705982(-)__16_29694001_29719001D;SPAN=15398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:57 GQ:30.8 PL:[30.8, 0.0, 106.7] SR:0 DR:14 LR:-30.77 LO:33.16);ALT=C[chr16:29705982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29802155	+	chr16	29808218	+	.	15	0	6180753_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6180753_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:29802155(+)-16:29808218(-)__16_29792001_29817001D;SPAN=6063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:102 GQ:22.1 PL:[22.1, 0.0, 223.4] SR:0 DR:15 LR:-21.88 LO:31.78);ALT=T[chr16:29808218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29814929	+	chr16	29816133	+	TTCAGGAGCAGGCAGCATCCCCAAATGCCGAGATCCACATCCTGAAGAATAAAGGCCGGAAGAGAA	0	7	6180785_1	0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTCAGGAGCAGGCAGCATCCCCAAATGCCGAGATCCACATCCTGAAGAATAAAGGCCGGAAGAGAA;MAPQ=60;MATEID=6180785_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_29792001_29817001_245C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:90 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.276 LO:12.77);ALT=A[chr16:29816133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29831874	+	chr16	29842196	+	.	13	0	6181076_1	30.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6181076_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:29831874(+)-16:29842196(-)__16_29841001_29866001D;SPAN=10322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:0 DR:13 LR:-30.18 LO:31.58);ALT=A[chr16:29842196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29831877	+	chr16	29841848	+	.	14	0	6181077_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6181077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:29831877(+)-16:29841848(-)__16_29841001_29866001D;SPAN=9971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:56 GQ:31.1 PL:[31.1, 0.0, 103.7] SR:0 DR:14 LR:-31.04 LO:33.29);ALT=T[chr16:29841848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29979576	+	chr16	29982728	+	.	7	36	6181766_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6181766_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_29963501_29988501_321C;SPAN=3152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:105 GQ:99 PL:[110.3, 0.0, 143.3] SR:36 DR:7 LR:-110.2 LO:110.5);ALT=G[chr16:29982728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	29982902	+	chr16	29984268	+	.	4	49	6181778_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGTG;MAPQ=60;MATEID=6181778_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_29963501_29988501_283C;SPAN=1366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:119 GQ:99 PL:[142.7, 0.0, 146.0] SR:49 DR:4 LR:-142.7 LO:142.7);ALT=G[chr16:29984268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30007713	+	chr16	30012078	+	AGCACGAGTGCTTCCAGGAGGAGCTGAGGAAAGCGCAAAGGAAATTACTGAAGGTGTCCCGGGACAAGAGTTTCCTCCTAGACCGACTTCTGCAGTACGAGAACGTGGATGAAGACTCTTCG	0	36	6181580_1	93.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AGCACGAGTGCTTCCAGGAGGAGCTGAGGAAAGCGCAAAGGAAATTACTGAAGGTGTCCCGGGACAAGAGTTTCCTCCTAGACCGACTTCTGCAGTACGAGAACGTGGATGAAGACTCTTCG;MAPQ=60;MATEID=6181580_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_16_29988001_30013001_103C;SPAN=4365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:94 GQ:93.5 PL:[93.5, 0.0, 133.1] SR:36 DR:0 LR:-93.37 LO:93.78);ALT=G[chr16:30012078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30008181	+	chr16	30012078	+	.	8	14	6181584_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6181584_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_16_29988001_30013001_103C;SPAN=3897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:91 GQ:35 PL:[35.0, 0.0, 183.5] SR:14 DR:8 LR:-34.76 LO:40.7);ALT=G[chr16:30012078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30012851	+	chr16	30016540	+	.	6	4	6181619_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6181619_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30012501_30037501_122C;SPAN=3689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:85 GQ:6.8 PL:[6.8, 0.0, 198.2] SR:4 DR:6 LR:-6.68 LO:17.69);ALT=G[chr16:30016540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30075855	+	chr16	30078767	+	.	40	0	6182052_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6182052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30075855(+)-16:30078767(-)__16_30061501_30086501D;SPAN=2912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:103 GQ:99 PL:[104.3, 0.0, 143.9] SR:0 DR:40 LR:-104.1 LO:104.5);ALT=A[chr16:30078767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30075855	+	chr16	30078550	+	.	100	0	6182051_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6182051_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30075855(+)-16:30078550(-)__16_30061501_30086501D;SPAN=2695;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:158 GQ:95.9 PL:[287.3, 0.0, 95.9] SR:0 DR:100 LR:-292.5 LO:292.5);ALT=A[chr16:30078550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30077166	+	chr16	30078769	+	.	44	0	6182055_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6182055_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30077166(+)-16:30078769(-)__16_30061501_30086501D;SPAN=1603;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:252 GQ:77.2 PL:[77.2, 0.0, 532.7] SR:0 DR:44 LR:-76.97 LO:96.82);ALT=C[chr16:30078769[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30077249	+	chr16	30078551	+	.	100	74	6182056_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAGG;MAPQ=60;MATEID=6182056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30061501_30086501_297C;SPAN=1302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:211 GQ:99 PL:[405.2, 0.0, 104.8] SR:74 DR:100 LR:-414.6 LO:414.6);ALT=G[chr16:30078551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30079036	+	chr16	30080135	+	.	21	0	6182065_1	45.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6182065_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30079036(+)-16:30080135(-)__16_30061501_30086501D;SPAN=1099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:88 GQ:45.5 PL:[45.5, 0.0, 167.6] SR:0 DR:21 LR:-45.48 LO:49.44);ALT=T[chr16:30080135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30087452	+	chr16	30093800	+	.	11	0	6181908_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6181908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30087452(+)-16:30093800(-)__16_30086001_30111001D;SPAN=6348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:80 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:0 DR:11 LR:-14.64 LO:22.95);ALT=G[chr16:30093800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30087463	+	chr16	30092518	+	.	28	0	6181909_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6181909_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30087463(+)-16:30092518(-)__16_30086001_30111001D;SPAN=5055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:85 GQ:69.5 PL:[69.5, 0.0, 135.5] SR:0 DR:28 LR:-69.4 LO:70.61);ALT=C[chr16:30092518[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30087796	+	chr16	30094067	+	AGAGATCTTGGTAGAGGAGAGCAACGTGCAGAGGGTGGACTCGCCAGTCACAGTGTGCGGCGACATCCATGGACAATTCTATGACCTCAAAGAGCTGTTCAGA	0	79	6181912_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GTA;INSERTION=AGAGATCTTGGTAGAGGAGAGCAACGTGCAGAGGGTGGACTCGCCAGTCACAGTGTGCGGCGACATCCATGGACAATTCTATGACCTCAAAGAGCTGTTCAGA;MAPQ=60;MATEID=6181912_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_16_30086001_30111001_3C;SPAN=6271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:132 GQ:93.2 PL:[225.2, 0.0, 93.2] SR:79 DR:0 LR:-227.9 LO:227.9);ALT=G[chr16:30094067[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30195046	+	chr16	30197917	+	AATGAGCCGGCAGGTGGTCCGCTCCAGCAAGTTCCGCCACGTGTTTGGACAGCCGGCCAAGGCCGACCAGTGCTATGAAGATGTGCGCGTCTCACAGACCACCTGGGACAGTGGCTTCTGTGCTGTCAACCCTAAGTTTGTGGCCCTGATCTGTGAGGCCAGCGGGGGAGGGGCCTTCCTGGTGCTGCCCCTGGGCA	41	109	6182552_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AATGAGCCGGCAGGTGGTCCGCTCCAGCAAGTTCCGCCACGTGTTTGGACAGCCGGCCAAGGCCGACCAGTGCTATGAAGATGTGCGCGTCTCACAGACCACCTGGGACAGTGGCTTCTGTGCTGTCAACCCTAAGTTTGTGGCCCTGATCTGTGAGGCCAGCGGGGGAGGGGCCTTCCTGGTGCTGCCCCTGGGCA;MAPQ=60;MATEID=6182552_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_30184001_30209001_269C;SPAN=2871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:125 DP:110 GQ:33.6 PL:[369.6, 33.6, 0.0] SR:109 DR:41 LR:-369.7 LO:369.7);ALT=G[chr16:30197917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30195046	+	chr16	30196527	+	.	163	22	6182551_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=6182551_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GACGAC;SCTG=c_16_30184001_30209001_269C;SPAN=1481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:171 DP:137 GQ:45.8 PL:[397.9, 45.8, 0.0] SR:22 DR:163 LR:-397.9 LO:397.9);ALT=G[chr16:30196527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30196728	+	chr16	30197917	+	.	3	81	6182556_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6182556_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_30184001_30209001_269C;SPAN=1189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:148 GQ:99 PL:[230.6, 0.0, 128.3] SR:81 DR:3 LR:-232.1 LO:232.1);ALT=G[chr16:30197917[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30435854	+	chr16	30440378	+	.	4	43	6183823_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6183823_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30429001_30454001_168C;SPAN=4524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:119 GQ:99 PL:[116.3, 0.0, 172.4] SR:43 DR:4 LR:-116.3 LO:116.9);ALT=A[chr16:30440378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30435905	+	chr16	30441102	+	.	31	0	6183824_1	75.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6183824_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30435905(+)-16:30441102(-)__16_30429001_30454001D;SPAN=5197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:100 GQ:75.2 PL:[75.2, 0.0, 167.6] SR:0 DR:31 LR:-75.24 LO:77.17);ALT=G[chr16:30441102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30484219	+	chr16	30485516	+	.	0	5	6184034_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6184034_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30478001_30503001_139C;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:108 GQ:12.6 PL:[0.0, 12.6, 287.1] SR:5 DR:0 LR:12.75 LO:7.966);ALT=G[chr16:30485516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30759848	+	chr16	30762422	+	.	24	0	6185777_1	48.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6185777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:30759848(+)-16:30762422(-)__16_30747501_30772501D;SPAN=2574;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:115 GQ:48.2 PL:[48.2, 0.0, 229.7] SR:0 DR:24 LR:-48.07 LO:54.89);ALT=C[chr16:30762422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30760236	+	chr16	30762423	+	.	0	21	6185780_1	39.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=6185780_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30747501_30772501_441C;SPAN=2187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:109 GQ:39.8 PL:[39.8, 0.0, 224.6] SR:21 DR:0 LR:-39.79 LO:47.21);ALT=G[chr16:30762423[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30768976	+	chr16	30770498	+	.	0	7	6185815_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6185815_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30747501_30772501_16C;SPAN=1522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:105 GQ:5.1 PL:[0.0, 5.1, 264.0] SR:7 DR:0 LR:5.34 LO:12.29);ALT=C[chr16:30770498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30900268	+	chr16	30903907	+	.	0	10	6185547_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6185547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30894501_30919501_173C;SPAN=3639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:98 GQ:6.5 PL:[6.5, 0.0, 230.9] SR:10 DR:0 LR:-6.459 LO:19.48);ALT=T[chr16:30903907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	30960841	+	chr16	30964505	+	.	6	2	6185953_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6185953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_30943501_30968501_144C;SPAN=3664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:79 GQ:1.5 PL:[0.0, 1.5, 194.7] SR:2 DR:6 LR:1.597 LO:10.88);ALT=G[chr16:30964505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31102665	+	chr16	31104631	+	.	4	31	6186469_1	81.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6186469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_31090501_31115501_236C;SPAN=1966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:115 GQ:81.2 PL:[81.2, 0.0, 196.7] SR:31 DR:4 LR:-81.08 LO:83.78);ALT=T[chr16:31104631[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31102666	+	chr16	31105876	+	.	32	20	6186471_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=6186471_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_31090501_31115501_120C;SPAN=3210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:119 GQ:99 PL:[103.1, 0.0, 185.6] SR:20 DR:32 LR:-103.1 LO:104.4);ALT=G[chr16:31105876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31104787	+	chr16	31105872	+	.	51	0	6186478_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6186478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:31104787(+)-16:31105872(-)__16_31090501_31115501D;SPAN=1085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:105 GQ:99 PL:[140.0, 0.0, 113.6] SR:0 DR:51 LR:-140.0 LO:140.0);ALT=A[chr16:31105872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31129213	+	chr16	31131507	+	.	0	18	6186651_1	34.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6186651_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_31115001_31140001_255C;SPAN=2294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:93 GQ:34.4 PL:[34.4, 0.0, 189.5] SR:18 DR:0 LR:-34.22 LO:40.51);ALT=C[chr16:31131507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31191545	+	chr16	31195178	+	.	9	0	6186844_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6186844_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:31191545(+)-16:31195178(-)__16_31188501_31213501D;SPAN=3633;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:116 GQ:1.5 PL:[0.0, 1.5, 283.8] SR:0 DR:9 LR:1.718 LO:16.41);ALT=A[chr16:31195178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31191548	+	chr16	31193832	+	ATTATACCCAACAAGCAACCCAA	86	25	6186845_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=ATTATACCCAACAAGCAACCCAA;MAPQ=60;MATEID=6186845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_31188501_31213501_357C;SPAN=2284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:121 GQ:13.7 PL:[277.7, 0.0, 13.7] SR:25 DR:86 LR:-291.4 LO:291.4);ALT=G[chr16:31193832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31193986	+	chr16	31195182	+	.	0	24	6186856_1	41.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6186856_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_31188501_31213501_29C;SPAN=1196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:142 GQ:41 PL:[41.0, 0.0, 301.7] SR:24 DR:0 LR:-40.75 LO:52.43);ALT=G[chr16:31195182[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31196550	+	chr16	31200442	+	.	9	0	6186870_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6186870_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:31196550(+)-16:31200442(-)__16_31188501_31213501D;SPAN=3892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:120 GQ:2.7 PL:[0.0, 2.7, 297.0] SR:0 DR:9 LR:2.802 LO:16.28);ALT=T[chr16:31200442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31885235	+	chr16	31895817	+	.	10	0	6189088_1	9.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6189088_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:31885235(+)-16:31895817(-)__16_31874501_31899501D;SPAN=10582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:0 DR:10 LR:-9.44 LO:20.03);ALT=C[chr16:31895817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	31885291	+	chr16	31896481	+	GACTGTTGACATTCAGGGATGTGGCCGTAGAATTCTCTTTGGAGGAGTGGGAACACCTGGAACCAGCTCAGAAGAATTTGTATCAGGATGTGATGTTAGAAAACTACAGAAACCTGGTCTCTCTG	0	14	6189090_1	20.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=GACTGTTGACATTCAGGGATGTGGCCGTAGAATTCTCTTTGGAGGAGTGGGAACACCTGGAACCAGCTCAGAAGAATTTGTATCAGGATGTGATGTTAGAAAACTACAGAAACCTGGTCTCTCTG;MAPQ=60;MATEID=6189090_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_31874501_31899501_19C;SPAN=11190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:95 GQ:20.6 PL:[20.6, 0.0, 208.7] SR:14 DR:0 LR:-20.48 LO:29.67);ALT=G[chr16:31896481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	32296411	+	chr16	32294446	+	.	11	0	6191350_1	21.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=6191350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:32294446(-)-16:32296411(+)__16_32291001_32316001D;SPAN=1965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=]chr16:32296411]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	32495601	+	chr16	32497776	+	.	24	6	6192421_1	66.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=TTAAACCTTTCTTTTCATTCATCAGTTTGGAAACACTGTTTTTGT;MAPQ=60;MATEID=6192421_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_32487001_32512001_413C;SPAN=2175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:95 GQ:66.8 PL:[66.8, 0.0, 162.5] SR:6 DR:24 LR:-66.69 LO:68.95);ALT=T[chr16:32497776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	32600335	+	chr16	32601844	+	.	40	17	6192885_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAGGCCTATGGTGACAAACTGAATATCCCCAGATAA;MAPQ=60;MATEID=6192885_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_32585001_32610001_34C;SPAN=1509;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:83 GQ:43.7 PL:[155.9, 0.0, 43.7] SR:17 DR:40 LR:-159.1 LO:159.1);ALT=A[chr16:32601844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	33075735	+	chr16	33074021	+	.	11	0	6196740_1	26.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6196740_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:33074021(-)-16:33075735(+)__16_33050501_33075501D;SPAN=1714;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:0 DR:11 LR:-26.02 LO:26.98);ALT=]chr16:33075735]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	33238416	+	chr16	33237191	+	.	32	0	6197586_1	34.0	.	DISC_MAPQ=13;EVDNC=DSCRD;IMPRECISE;MAPQ=13;MATEID=6197586_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:33237191(-)-16:33238416(+)__16_33222001_33247001D;SPAN=1225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:263 GQ:34.6 PL:[34.6, 0.0, 602.3] SR:0 DR:32 LR:-34.38 LO:64.95);ALT=]chr16:33238416]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	33374049	+	chr16	33379406	+	TTTAGGT	46	28	6198019_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;INSERTION=TTTAGGT;MAPQ=60;MATEID=6198019_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_16_33369001_33394001_144C;SPAN=5357;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:149 GQ:99 PL:[184.1, 0.0, 177.5] SR:28 DR:46 LR:-184.1 LO:184.1);ALT=C[chr16:33379406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	33891555	+	chr16	33888137	+	.	28	1	6203098_1	59.0	.	DISC_MAPQ=46;EVDNC=TSI_L;HOMSEQ=GATGATTCC;MAPQ=22;MATEID=6203098_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_16_33883501_33908501_239C;SPAN=3418;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:121 GQ:59.9 PL:[59.9, 0.0, 231.5] SR:1 DR:28 LR:-59.65 LO:65.48);ALT=]chr16:33891555]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	54953121	+	chr16	54959013	+	ATTTTTCATTTCAACATTTCCAGTGGCATCCTCCTTATCTTCAGAATCTCCTCCTTCCAATAGCCAGTACAGTAGCTCCATTATGAATTGCAGACT	0	10	6216515_1	26.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=ATTTTTCATTTCAACATTTCCAGTGGCATCCTCCTTATCTTCAGAATCTCCTCCTTCCAATAGCCAGTACAGTAGCTCCATTATGAATTGCAGACT;MAPQ=60;MATEID=6216515_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_54953501_54978501_190C;SPAN=5892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:10 DR:0 LR:-26.24 LO:26.3);ALT=T[chr16:54959013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	55543264	+	chr16	55559417	+	.	8	8	6217324_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6217324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_55541501_55566501_143C;SPAN=16153;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:57 GQ:27.5 PL:[27.5, 0.0, 110.0] SR:8 DR:8 LR:-27.47 LO:30.31);ALT=G[chr16:55559417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56466648	+	chr16	56468241	+	.	0	8	6218797_1	15.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=6218797_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_56448001_56473001_242C;SPAN=1593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:8 DR:0 LR:-15.3 LO:18.03);ALT=G[chr16:56468241[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56481901	+	chr16	56484996	+	.	0	34	6218862_1	90.0	.	EVDNC=ASSMB;HOMSEQ=TAC;MAPQ=60;MATEID=6218862_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_56472501_56497501_147C;SPAN=3095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:80 GQ:90.5 PL:[90.5, 0.0, 103.7] SR:34 DR:0 LR:-90.56 LO:90.61);ALT=C[chr16:56484996[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56716468	+	chr16	56717869	+	.	12	0	6219366_1	32.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6219366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:56716468(+)-16:56717869(-)__16_56717501_56742501D;SPAN=1401;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:28 GQ:32 PL:[32.0, 0.0, 35.3] SR:0 DR:12 LR:-32.03 LO:32.04);ALT=T[chr16:56717869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56764172	+	chr16	56782209	+	.	9	0	6219694_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6219694_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:56764172(+)-16:56782209(-)__16_56766501_56791501D;SPAN=18037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:0 DR:9 LR:-22.12 LO:22.58);ALT=A[chr16:56782209[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	56966303	+	chr16	56969146	+	.	0	19	6219991_1	49.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6219991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_56962501_56987501_115C;SPAN=2843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:51 GQ:49.1 PL:[49.1, 0.0, 72.2] SR:19 DR:0 LR:-48.9 LO:49.2);ALT=G[chr16:56969146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57105772	+	chr16	57104515	+	.	29	1	6220197_1	80.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=TGCT;MAPQ=60;MATEID=6220197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57085001_57110001_13C;SPAN=1257;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:68 GQ:80.6 PL:[80.6, 0.0, 83.9] SR:1 DR:29 LR:-80.61 LO:80.61);ALT=]chr16:57105772]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	57207785	+	chr16	57219733	+	.	19	8	6220383_1	57.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=CTAC;MAPQ=60;MATEID=6220383_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57207501_57232501_49C;SPAN=11948;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:82 GQ:57.2 PL:[57.2, 0.0, 139.7] SR:8 DR:19 LR:-57.01 LO:59.01);ALT=C[chr16:57219733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57279317	+	chr16	57282448	+	CTCCTCCGCCTCTGATGCAGAATTTGATGCTGTGGTTGGATATTTAGAGGACATTATCATG	3	18	6220486_1	62.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=TGTGGTTGGATATTTAGAGGACATTATCATGG;INSERTION=CTCCTCCGCCTCTGATGCAGAATTTGATGCTGTGGTTGGATATTTAGAGGACATTATCATG;MAPQ=60;MATEID=6220486_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_57281001_57306001_233C;SECONDARY;SPAN=3131;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:21 DP:26 GQ:0.3 PL:[62.7, 0.3, 0.0] SR:18 DR:3 LR:-65.96 LO:65.96);ALT=T[chr16:57282448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57481490	+	chr16	57484951	+	.	13	3	6220945_1	27.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6220945_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57477001_57502001_254C;SPAN=3461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:3 DR:13 LR:-27.52 LO:31.83);ALT=G[chr16:57484951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57496690	+	chr16	57499861	+	.	9	0	6220963_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6220963_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:57496690(+)-16:57499861(-)__16_57477001_57502001D;SPAN=3171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:68 GQ:11.3 PL:[11.3, 0.0, 153.2] SR:0 DR:9 LR:-11.29 LO:18.62);ALT=T[chr16:57499861[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57496723	+	chr16	57503076	+	GTGGCCAATTCGATTCGGAGGGTCTTCATCGCTGAGGTTCCCATAATAGCCATTGACTGGGTTCAGATTGATGCCAATTCCTCAGTTCTTCATGATGAATTCATTGCTCACAGGCTTGGATTAATTCCCCTCATTAGTGATGACATTGTGGACAAGCTGCAGTACTCTCG	0	17	6220966_1	48.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=GTGGCCAATTCGATTCGGAGGGTCTTCATCGCTGAGGTTCCCATAATAGCCATTGACTGGGTTCAGATTGATGCCAATTCCTCAGTTCTTCATGATGAATTCATTGCTCACAGGCTTGGATTAATTCCCCTCATTAGTGATGACATTGTGGACAAGCTGCAGTACTCTCG;MAPQ=60;MATEID=6220966_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_16_57477001_57502001_161C;SPAN=6353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:27 GQ:15.8 PL:[48.8, 0.0, 15.8] SR:17 DR:0 LR:-49.67 LO:49.67);ALT=G[chr16:57503076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	57725300	-	chr16	57727956	+	.	3	2	6221379_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGGGTGCA;MAPQ=60;MATEID=6221379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57722001_57747001_159C;SPAN=2656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:61 GQ:3 PL:[0.0, 3.0, 151.8] SR:2 DR:3 LR:3.322 LO:6.992);ALT=[chr16:57727956[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	57725395	+	chr16	57727847	+	.	83	50	6221380_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6221380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_57722001_57747001_146C;SPAN=2452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:22 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:50 DR:83 LR:-340.0 LO:340.0);ALT=G[chr16:57727847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58555223	+	chr16	58557274	+	.	3	3	6222927_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6222927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_58555001_58580001_28C;SPAN=2051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:46 GQ:0.8 PL:[0.8, 0.0, 109.7] SR:3 DR:3 LR:-0.7415 LO:7.501);ALT=T[chr16:58557274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58624545	+	chr16	58663331	+	CCAG	69	33	6223031_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;INSERTION=CCAG;MAPQ=60;MATEID=6223031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_58653001_58678001_43C;SPAN=38786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:11 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:33 DR:69 LR:-254.2 LO:254.2);ALT=T[chr16:58663331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58657315	+	chr16	58663628	+	.	7	5	6223035_1	29.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TCACCT;MAPQ=60;MATEID=6223035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_58653001_58678001_116C;SPAN=6313;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:36 GQ:29.9 PL:[29.9, 0.0, 56.3] SR:5 DR:7 LR:-29.86 LO:30.34);ALT=T[chr16:58663628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58658700	+	chr16	58663632	+	.	13	4	6223036_1	36.0	.	DISC_MAPQ=45;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6223036_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_58653001_58678001_144C;SPAN=4932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:36 GQ:36.5 PL:[36.5, 0.0, 49.7] SR:4 DR:13 LR:-36.46 LO:36.59);ALT=T[chr16:58663632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	58757809	+	chr16	58768044	+	.	0	24	6223317_1	60.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6223317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_58751001_58776001_156C;SPAN=10235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:68 GQ:60.8 PL:[60.8, 0.0, 103.7] SR:24 DR:0 LR:-60.8 LO:61.43);ALT=G[chr16:58768044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66586696	+	chr16	66596974	+	.	32	3	6234080_1	92.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6234080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66566501_66591501_200C;SPAN=10278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:59 GQ:50 PL:[92.9, 0.0, 50.0] SR:3 DR:32 LR:-93.63 LO:93.63);ALT=G[chr16:66596974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66586697	+	chr16	66592092	+	.	55	61	6234081_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6234081_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66566501_66591501_80C;SPAN=5395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:56 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:61 DR:55 LR:-283.9 LO:283.9);ALT=G[chr16:66592092[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66586699	+	chr16	66599788	+	.	13	10	6234083_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6234083_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66566501_66591501_46C;SPAN=13089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:51 GQ:59 PL:[59.0, 0.0, 62.3] SR:10 DR:13 LR:-58.81 LO:58.82);ALT=G[chr16:66599788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66592252	+	chr16	66597025	+	.	0	16	6233960_1	26.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6233960_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66591001_66616001_107C;SPAN=4773;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:97 GQ:26.6 PL:[26.6, 0.0, 208.1] SR:16 DR:0 LR:-26.54 LO:34.77);ALT=G[chr16:66597025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66592253	+	chr16	66599789	+	.	2	22	6233961_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=6233961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66591001_66616001_67C;SPAN=7536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:92 GQ:47.9 PL:[47.9, 0.0, 173.3] SR:22 DR:2 LR:-47.7 LO:51.81);ALT=T[chr16:66599789[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66597122	+	chr16	66599788	+	.	0	83	6233968_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=6233968_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66591001_66616001_110C;SPAN=2666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:95 GQ:18.9 PL:[267.3, 18.9, 0.0] SR:83 DR:0 LR:-269.1 LO:269.1);ALT=T[chr16:66599788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66638856	+	chr16	66642211	+	.	0	26	6234294_1	75.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6234294_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66615501_66640501_93C;SPAN=3355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:26 DP:24 GQ:6.9 PL:[75.9, 6.9, 0.0] SR:26 DR:0 LR:-75.92 LO:75.92);ALT=G[chr16:66642211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66860685	+	chr16	66864748	+	.	15	2	6234600_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6234600_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_66836001_66861001_259C;SPAN=4063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:20 GQ:4.4 PL:[44.0, 0.0, 4.4] SR:2 DR:15 LR:-45.99 LO:45.99);ALT=T[chr16:66864748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	66966205	+	chr16	66967517	+	GCATGCTCTGAGGCATGGGTCCCCGGAGTAATGTGCACGTCCAT	0	59	6234867_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GCATGCTCTGAGGCATGGGTCCCCGGAGTAATGTGCACGTCCAT;MAPQ=60;MATEID=6234867_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_66958501_66983501_129C;SPAN=1312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:81 GQ:21.2 PL:[173.0, 0.0, 21.2] SR:59 DR:0 LR:-179.3 LO:179.3);ALT=T[chr16:66967517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67144143	+	chr16	67154014	+	.	3	3	6235291_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6235291_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_67130001_67155001_269C;SPAN=9871;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:65 GQ:4.2 PL:[0.0, 4.2, 165.0] SR:3 DR:3 LR:4.406 LO:6.878);ALT=G[chr16:67154014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67190581	+	chr16	67193739	+	.	15	0	6235186_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6235186_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67190581(+)-16:67193739(-)__16_67179001_67204001D;SPAN=3158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:47 GQ:36.8 PL:[36.8, 0.0, 76.4] SR:0 DR:15 LR:-36.78 LO:37.57);ALT=C[chr16:67193739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67261164	+	chr16	67262255	+	.	54	0	6235464_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6235464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67261164(+)-16:67262255(-)__16_67252501_67277501D;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:58 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:0 DR:54 LR:-171.6 LO:171.6);ALT=A[chr16:67262255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67487619	+	chr16	67514860	+	.	29	28	6235890_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6235890_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_67497501_67522501_242C;SPAN=27241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:31 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:28 DR:29 LR:-138.6 LO:138.6);ALT=C[chr16:67514860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67515411	+	chr16	67518010	+	.	11	0	6235922_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6235922_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67515411(+)-16:67518010(-)__16_67497501_67522501D;SPAN=2599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:58 GQ:20.6 PL:[20.6, 0.0, 119.6] SR:0 DR:11 LR:-20.6 LO:24.64);ALT=G[chr16:67518010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67596627	+	chr16	67605049	+	.	5	4	6236237_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6236237_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_67595501_67620501_45C;SPAN=8422;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:44 GQ:11.3 PL:[11.3, 0.0, 93.8] SR:4 DR:5 LR:-11.19 LO:15.09);ALT=G[chr16:67605049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67866449	+	chr16	67867653	+	.	18	10	6236831_1	43.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6236831_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_67865001_67890001_80C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:73 GQ:43.1 PL:[43.1, 0.0, 132.2] SR:10 DR:18 LR:-42.94 LO:45.56);ALT=C[chr16:67867653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67880931	+	chr16	67902397	+	.	18	0	6236864_1	52.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=6236864_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67880931(+)-16:67902397(-)__16_67865001_67890001D;SPAN=21466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:16 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:0 DR:18 LR:-52.81 LO:52.81);ALT=A[chr16:67902397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	67880931	+	chr16	67899003	+	.	15	0	6236863_1	46.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=6236863_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:67880931(+)-16:67899003(-)__16_67865001_67890001D;SPAN=18072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:16 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:0 DR:15 LR:-46.21 LO:46.21);ALT=A[chr16:67899003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	68300625	+	chr16	68308591	+	.	3	8	6237939_1	23.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6237939_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_68306001_68331001_155C;SPAN=7966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:34 GQ:23.9 PL:[23.9, 0.0, 56.9] SR:8 DR:3 LR:-23.8 LO:24.62);ALT=G[chr16:68308591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69154588	+	chr16	69166413	+	.	10	0	6239612_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6239612_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:69154588(+)-16:69166413(-)__16_69163501_69188501D;SPAN=11825;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:24 GQ:26.6 PL:[26.6, 0.0, 29.9] SR:0 DR:10 LR:-26.51 LO:26.53);ALT=G[chr16:69166413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69345435	+	chr16	69349906	+	.	26	17	6239905_1	96.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=TCCAG;MAPQ=60;MATEID=6239905_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_16_69335001_69360001_123C;SPAN=4471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:47 GQ:17 PL:[96.2, 0.0, 17.0] SR:17 DR:26 LR:-99.25 LO:99.25);ALT=G[chr16:69349906[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69458760	+	chr16	69481051	+	.	0	21	6240182_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6240182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69457501_69482501_159C;SPAN=22291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:71 GQ:50.3 PL:[50.3, 0.0, 119.6] SR:21 DR:0 LR:-50.09 LO:51.75);ALT=G[chr16:69481051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	69761829	-	chr16	69762896	+	.	41	41	6241149_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TCAAG;MAPQ=60;MATEID=6241149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69751501_69776501_123C;SPAN=1067;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:56 GQ:18 PL:[198.0, 18.0, 0.0] SR:41 DR:41 LR:-198.0 LO:198.0);ALT=[chr16:69762896[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr16	69791912	+	chrX	70503589	-	.	12	0	7445429_1	34.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=7445429_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:69791912(+)-23:70503589(+)__23_70486501_70511501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:18 GQ:8.3 PL:[34.7, 0.0, 8.3] SR:0 DR:12 LR:-35.58 LO:35.58);ALT=A]chrX:70503589];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr16	69820983	+	chr16	69832583	+	.	0	8	6240880_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6240880_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_69800501_69825501_101C;SPAN=11600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:20 GQ:20.9 PL:[20.9, 0.0, 27.5] SR:8 DR:0 LR:-20.99 LO:21.04);ALT=G[chr16:69832583[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	74587100	+	chr16	70112512	+	.	0	10	6250379_1	26.0	.	EVDNC=ASSMB;HOMSEQ=TGGGCAACA;MAPQ=49;MATEID=6250379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_74578001_74603001_138C;SPAN=4474588;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:25 GQ:26.3 PL:[26.3, 0.0, 32.9] SR:10 DR:0 LR:-26.24 LO:26.3);ALT=]chr16:74587100]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	70333257	+	chr16	70349870	+	TTGAGCAACTTGCATCTTAAGGAAGAGAAAATCAAACCAGATACCAATGGTGCTGTTGTCAAGACCAATGCCAATGCAGAGAAGACAGATGAAGAAGAGAA	5	17	6242694_1	51.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTGAGCAACTTGCATCTTAAGGAAGAGAAAATCAAACCAGATACCAATGGTGCTGTTGTCAAGACCAATGCCAATGCAGAGAAGACAGATGAAGAAGAGAA;MAPQ=60;MATEID=6242694_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_16_70339501_70364501_38C;SPAN=16613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:28 GQ:15.5 PL:[51.8, 0.0, 15.5] SR:17 DR:5 LR:-52.87 LO:52.87);ALT=G[chr16:70349870[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	70553636	+	chr16	70557276	+	.	6	4	6243220_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6243220_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_70535501_70560501_251C;SPAN=3640;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:4 DR:6 LR:-11.24 LO:16.84);ALT=T[chr16:70557276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	70599427	+	chr16	70601312	+	.	3	2	6243149_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6243149_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_70584501_70609501_165C;SPAN=1885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:56 GQ:1.4 PL:[1.4, 0.0, 133.4] SR:2 DR:3 LR:-1.333 LO:9.437);ALT=G[chr16:70601312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	74330817	+	chr16	74334009	+	.	31	0	6249585_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6249585_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:74330817(+)-16:74334009(-)__16_74333001_74358001D;SPAN=3192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:38 GQ:0.3 PL:[92.4, 0.3, 0.0] SR:0 DR:31 LR:-97.71 LO:97.71);ALT=C[chr16:74334009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	74330849	+	chr17	64193917	+	.	17	0	6470527_1	42.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6470527_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:74330849(+)-17:64193917(-)__17_64190001_64215001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.57 LO:43.16);ALT=C[chr17:64193917[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr16	75339081	+	chr16	75428986	+	.	3	5	6252171_1	15.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=6252171_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_16_75411001_75436001_133C;SPAN=89905;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:29 GQ:15.2 PL:[15.2, 0.0, 54.8] SR:5 DR:3 LR:-15.25 LO:16.52);ALT=C[chr16:75428986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75446653	+	chr16	75467186	+	.	8	2	6252242_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6252242_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75435501_75460501_126C;SPAN=20533;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:2 DR:8 LR:-19.14 LO:21.04);ALT=C[chr16:75467186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75446654	+	chr16	75448475	+	.	8	14	6252243_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=6252243_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_75435501_75460501_264C;SPAN=1821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:73 GQ:43.1 PL:[43.1, 0.0, 132.2] SR:14 DR:8 LR:-42.94 LO:45.56);ALT=T[chr16:75448475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75448594	+	chr16	75467184	+	.	29	25	6252350_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=6252350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75460001_75485001_75C;SPAN=18590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:39 DP:35 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:25 DR:29 LR:-115.5 LO:115.5);ALT=C[chr16:75467184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75485739	+	chr16	75498366	+	.	0	13	6252465_1	28.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6252465_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75484501_75509501_292C;SPAN=12627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:53 GQ:28.7 PL:[28.7, 0.0, 98.0] SR:13 DR:0 LR:-28.55 LO:30.78);ALT=T[chr16:75498366[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75600418	+	chr16	75601934	+	AACACAGATGCGTGGAGTCCGCGAAGATTCGAGCGAAATATCCCGACAGGGTTCC	71	99	6252445_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GGTGA;INSERTION=AACACAGATGCGTGGAGTCCGCGAAGATTCGAGCGAAATATCCCGACAGGGTTCC;MAPQ=60;MATEID=6252445_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_75582501_75607501_157C;SPAN=1516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:62 GQ:37.3 PL:[409.3, 37.3, 0.0] SR:99 DR:71 LR:-409.3 LO:409.3);ALT=G[chr16:75601934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75602107	+	chr16	75611175	+	.	7	14	6252558_1	62.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6252558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75607001_75632001_167C;SPAN=9068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:22 GQ:5.7 PL:[62.7, 5.7, 0.0] SR:14 DR:7 LR:-61.26 LO:61.26);ALT=G[chr16:75611175[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75661893	+	chr16	75663312	+	TGATGTTGTTGGAGTCCGTGAGAAACATGGCGACTCGATCAATGCCCATGCCCCAGCCAGCTGTGGGGGGCAGCCCATATTCCAGGGCAGTACAGAAGTTTTCATCTATGAACATGGCCTCATCATCACCTGCAGCCTTGG	0	32	6252709_1	89.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TGATGTTGTTGGAGTCCGTGAGAAACATGGCGACTCGATCAATGCCCATGCCCCAGCCAGCTGTGGGGGGCAGCCCATATTCCAGGGCAGTACAGAAGTTTTCATCTATGAACATGGCCTCATCATCACCTGCAGCCTTGG;MAPQ=60;MATEID=6252709_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_75656001_75681001_172C;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:62 GQ:59.3 PL:[89.0, 0.0, 59.3] SR:32 DR:0 LR:-89.1 LO:89.1);ALT=T[chr16:75663312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75674247	+	chr16	75675462	+	.	5	14	6252732_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6252732_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_75656001_75681001_30C;SPAN=1215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:50 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:14 DR:5 LR:-42.57 LO:43.16);ALT=G[chr16:75675462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	75675664	+	chr16	75681490	+	.	18	0	6252737_1	52.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6252737_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:75675664(+)-16:75681490(-)__16_75656001_75681001D;SPAN=5826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:27 GQ:12.5 PL:[52.1, 0.0, 12.5] SR:0 DR:18 LR:-53.38 LO:53.38);ALT=G[chr16:75681490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	76539133	+	chr16	76544026	+	C	0	60	6253873_1	99.0	.	EVDNC=ASSMB;INSERTION=C;MAPQ=60;MATEID=6253873_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_76538001_76563001_111C;SPAN=4893;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:29 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:60 DR:0 LR:-178.2 LO:178.2);ALT=G[chr16:76544026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	83841726	+	chr16	83845022	+	.	14	0	6265374_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6265374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:83841726(+)-16:83845022(-)__16_83839001_83864001D;SPAN=3296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:85 GQ:23.3 PL:[23.3, 0.0, 181.7] SR:0 DR:14 LR:-23.19 LO:30.41);ALT=G[chr16:83845022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	83841728	+	chr16	83842910	+	GCAGACACTCCTGCAGCAGATGCAAGATAAATTTCAGACCATGTCTGACCAGATCATTGGGAGAA	73	137	6265376_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=GGT;INSERTION=GCAGACACTCCTGCAGCAGATGCAAGATAAATTTCAGACCATGTCTGACCAGATCATTGGGAGAA;MAPQ=60;MATEID=6265376_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_83839001_83864001_27C;SPAN=1182;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:192 DP:83 GQ:51.7 PL:[567.7, 51.7, 0.0] SR:137 DR:73 LR:-567.7 LO:567.7);ALT=T[chr16:83842910[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	83843032	+	chr16	83845024	+	.	0	77	6265378_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=6265378_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_83839001_83864001_161C;SPAN=1992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:89 GQ:14.1 PL:[244.2, 14.1, 0.0] SR:77 DR:0 LR:-248.5 LO:248.5);ALT=T[chr16:83845024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	84600564	+	chr16	84651107	+	TACGACCTCCTTCACCAGGGTCTTGTCCGTCCCGGTTTTGGCGCGCTGCAGCCCGCTGACGTTCTCACCGATCCACGTGATGAGGGCAAACTTGGACCTCTTGCTCATGGCATCCCCGGTGGTGAAGCGCACGAAGGCAAACAACCGGACGTCAT	2	100	6266907_1	99.0	.	DISC_MAPQ=18;EVDNC=TSI_G;HOMSEQ=CTGTG;INSERTION=TACGACCTCCTTCACCAGGGTCTTGTCCGTCCCGGTTTTGGCGCGCTGCAGCCCGCTGACGTTCTCACCGATCCACGTGATGAGGGCAAACTTGGACCTCTTGCTCATGGCATCCCCGGTGGTGAAGCGCACGAAGGCAAACAACCGGACGTCAT;MAPQ=60;MATEID=6266907_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_84647501_84672501_75C;SPAN=50543;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:48 GQ:27 PL:[297.0, 27.0, 0.0] SR:100 DR:2 LR:-297.1 LO:297.1);ALT=G[chr16:84651107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	84600564	+	chr16	84623711	+	.	6	45	6266855_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6266855_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_84623001_84648001_230C;SPAN=23147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:29 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:45 DR:6 LR:-148.5 LO:148.5);ALT=G[chr16:84623711[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	84623821	+	chr16	84651104	+	.	17	0	6266908_1	45.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6266908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:84623821(+)-16:84651104(-)__16_84647501_84672501D;SPAN=27283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:40 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:0 DR:17 LR:-45.28 LO:45.31);ALT=T[chr16:84651104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	84623920	+	chr16	84651442	+	.	37	0	6266910_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6266910_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:84623920(+)-16:84651442(-)__16_84647501_84672501D;SPAN=27522;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:70 GQ:66.8 PL:[103.1, 0.0, 66.8] SR:0 DR:37 LR:-103.6 LO:103.6);ALT=G[chr16:84651442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85302493	+	chr16	85304391	+	.	52	33	6267974_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6267974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85284501_85309501_134C;SPAN=1898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:17 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:33 DR:52 LR:-224.5 LO:224.5);ALT=G[chr16:85304391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85699954	+	chr16	85701744	+	.	4	3	6268832_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6268832_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85701001_85726001_260C;SPAN=1790;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:26 GQ:9.5 PL:[9.5, 0.0, 52.4] SR:3 DR:4 LR:-9.461 LO:11.24);ALT=G[chr16:85701744[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85712272	+	chr16	85721066	+	TGATTTAACAGGAGCTTCGTAAGTTCCATGTAGTAAGGGCTGGGCATTGGGGTAAAAGTTTCTTCCTTTCGTTCATGATCCCTCATCTTCTCCAACTTTT	0	18	6268853_1	44.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGATTTAACAGGAGCTTCGTAAGTTCCATGTAGTAAGGGCTGGGCATTGGGGTAAAAGTTTCTTCCTTTCGTTCATGATCCCTCATCTTCTCCAACTTTT;MAPQ=60;MATEID=6268853_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_85701001_85726001_16C;SPAN=8794;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:57 GQ:44 PL:[44.0, 0.0, 93.5] SR:18 DR:0 LR:-43.98 LO:44.99);ALT=A[chr16:85721066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85715289	+	chr16	85721066	+	.	0	9	6268856_1	2.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6268856_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CATCCATC;SCTG=c_16_85701001_85726001_16C;SPAN=5777;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:59 GQ:2.2 PL:[2.2, 0.0, 72.0] SR:9 DR:0 LR:-2.015 LO:7.655);ALT=T[chr16:85721066[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85721220	+	chr16	85722479	+	.	15	0	6268869_1	33.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=6268869_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85721220(+)-16:85722479(-)__16_85701001_85726001D;SPAN=1259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:0 DR:15 LR:-33.8 LO:35.92);ALT=A[chr16:85722479[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85741674	+	chr16	85768796	+	.	2	5	6269008_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6269008_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_85725501_85750501_182C;SPAN=27122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:31 GQ:14.9 PL:[14.9, 0.0, 57.8] SR:5 DR:2 LR:-14.71 LO:16.28);ALT=T[chr16:85768796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85744084	+	chr16	85784586	+	.	13	0	6269247_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6269247_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85744084(+)-16:85784586(-)__16_85774501_85799501D;SPAN=40502;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:18 GQ:5 PL:[38.0, 0.0, 5.0] SR:0 DR:13 LR:-39.41 LO:39.41);ALT=G[chr16:85784586[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85833358	+	chr16	85834808	+	.	37	29	6269443_1	75.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6269443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85823501_85848501_176C;SPAN=1450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:333 GQ:75 PL:[75.0, 0.0, 731.9] SR:29 DR:37 LR:-74.83 LO:106.4);ALT=G[chr16:85834808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85833390	+	chr16	85839338	+	.	8	0	6269446_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6269446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85833390(+)-16:85839338(-)__16_85823501_85848501D;SPAN=5948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:0 DR:8 LR:-0.6702 LO:14.89);ALT=C[chr16:85839338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85833409	+	chr16	85838538	+	.	186	0	6269447_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6269447_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85833409(+)-16:85838538(-)__16_85823501_85848501D;SPAN=5129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:186 DP:114 GQ:50.2 PL:[551.2, 50.2, 0.0] SR:0 DR:186 LR:-551.2 LO:551.2);ALT=G[chr16:85838538[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85834884	+	chr16	85838542	+	.	19	97	6269451_1	99.0	.	DISC_MAPQ=15;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6269451_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_16_85823501_85848501_94C;SPAN=3658;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:115 DP:204 GQ:99 PL:[324.5, 0.0, 169.4] SR:97 DR:19 LR:-326.9 LO:326.9);ALT=G[chr16:85838542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85834884	+	chr16	85839339	+	AAAGTGTTGTGAAGAGCGAAGACTTTTCGCTCCCAGCTTATATGGATCGGCGTGACCACCCCTTGCCGGAGGTGGCCCATGTCAAGCACCTGTCTGCCAGCCAGAAGGCACTGAAGGAGAAGGAGAAGGCCTCCTGGAGCAGCCTCTCCATGGATGAGAAAGTCGAGT	4	199	6269452_1	99.0	.	DISC_MAPQ=31;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AAAGTGTTGTGAAGAGCGAAGACTTTTCGCTCCCAGCTTATATGGATCGGCGTGACCACCCCTTGCCGGAGGTGGCCCATGTCAAGCACCTGTCTGCCAGCCAGAAGGCACTGAAGGAGAAGGAGAAGGCCTCCTGGAGCAGCCTCTCCATGGATGAGAAAGTCGAGT;MAPQ=60;MATEID=6269452_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_85823501_85848501_94C;SPAN=4455;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:202 DP:149 GQ:54.4 PL:[597.4, 54.4, 0.0] SR:199 DR:4 LR:-597.4 LO:597.4);ALT=G[chr16:85839339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85932830	+	chr16	85936619	+	.	31	3	6269352_1	88.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6269352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_85921501_85946501_15C;SPAN=3789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:63 GQ:62.3 PL:[88.7, 0.0, 62.3] SR:3 DR:31 LR:-88.77 LO:88.77);ALT=G[chr16:85936619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85932853	+	chr16	85942593	+	.	17	0	6269353_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6269353_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:85932853(+)-16:85942593(-)__16_85921501_85946501D;SPAN=9740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:55 GQ:41.3 PL:[41.3, 0.0, 90.8] SR:0 DR:17 LR:-41.22 LO:42.29);ALT=C[chr16:85942593[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	85936796	+	chr16	85943090	+	CCTGGGCAGTTTTTAAAGGGAAGTTTAAAGAAGGGGACAAAGCTGAACCAGCCACTTGGAAGACGAGGTTACGCTGTGCTTTGAATAAGAGCCCAGATTTTGAGGAAGTGACGGACCGGTCCCAACTGGACATTTCCGAGCCATACAAAGTTTACCGAATTGTTCCTGAGGAAGAGCAAAAAT	0	29	6269360_1	79.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CCTGGGCAGTTTTTAAAGGGAAGTTTAAAGAAGGGGACAAAGCTGAACCAGCCACTTGGAAGACGAGGTTACGCTGTGCTTTGAATAAGAGCCCAGATTTTGAGGAAGTGACGGACCGGTCCCAACTGGACATTTCCGAGCCATACAAAGTTTACCGAATTGTTCCTGAGGAAGAGCAAAAAT;MAPQ=60;MATEID=6269360_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_85921501_85946501_26C;SPAN=6294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:59 GQ:63.2 PL:[79.7, 0.0, 63.2] SR:29 DR:0 LR:-79.84 LO:79.84);ALT=G[chr16:85943090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	86379126	+	chr16	86385686	-	.	14	0	6270061_1	32.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6270061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:86379126(+)-16:86385686(+)__16_86362501_86387501D;SPAN=6560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:49 GQ:32.9 PL:[32.9, 0.0, 85.7] SR:0 DR:14 LR:-32.94 LO:34.25);ALT=C]chr16:86385686];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr16	86622031	+	chr16	86621014	+	.	50	0	6270611_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6270611_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:86621014(-)-16:86622031(+)__16_86607501_86632501D;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:72 GQ:26.9 PL:[145.7, 0.0, 26.9] SR:0 DR:50 LR:-149.9 LO:149.9);ALT=]chr16:86622031]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	87773402	+	chr16	87771949	+	.	59	0	6272747_1	99.0	.	DISC_MAPQ=14;EVDNC=DSCRD;IMPRECISE;MAPQ=14;MATEID=6272747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:87771949(-)-16:87773402(+)__16_87759001_87784001D;SPAN=1453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:67 GQ:14.7 PL:[191.4, 14.7, 0.0] SR:0 DR:59 LR:-192.0 LO:192.0);ALT=]chr16:87773402]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr16	87795686	+	chr16	87799496	+	.	9	0	6272684_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6272684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:87795686(+)-16:87799496(-)__16_87783501_87808501D;SPAN=3810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:52 GQ:15.8 PL:[15.8, 0.0, 108.2] SR:0 DR:9 LR:-15.62 LO:19.77);ALT=G[chr16:87799496[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88311285	+	chr16	88312817	+	.	8	0	6273616_1	17.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6273616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88311285(+)-16:88312817(-)__16_88298001_88323001D;SPAN=1532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:32 GQ:17.9 PL:[17.9, 0.0, 57.5] SR:0 DR:8 LR:-17.74 LO:19.02);ALT=A[chr16:88312817[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88636974	+	chr16	88643516	+	.	17	8	6274208_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6274208_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_88641001_88666001_263C;SPAN=6542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:21 DP:26 GQ:0.3 PL:[62.7, 0.3, 0.0] SR:8 DR:17 LR:-65.96 LO:65.96);ALT=G[chr16:88643516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88709980	+	chr16	88712523	+	.	0	85	6274383_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6274383_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_88690001_88715001_34C;SPAN=2543;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:247 GQ:99 PL:[213.7, 0.0, 385.4] SR:85 DR:0 LR:-213.7 LO:216.4);ALT=C[chr16:88712523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88710010	+	chr16	88713161	+	.	8	0	6274384_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6274384_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88710010(+)-16:88713161(-)__16_88690001_88715001D;SPAN=3151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:136 GQ:10.2 PL:[0.0, 10.2, 349.8] SR:0 DR:8 LR:10.44 LO:13.6);ALT=C[chr16:88713161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88714522	+	chr16	88717364	+	.	0	54	6274412_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6274412_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_88714501_88739501_115C;SPAN=2842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:132 GQ:99 PL:[142.7, 0.0, 175.7] SR:54 DR:0 LR:-142.5 LO:142.7);ALT=A[chr16:88717364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88724440	+	chr16	88729418	+	GTCCTGGTGCAGAGTGACGCTCAGGGAGGAGTTGATGGGCAGAACCAGCTCTTCATCGCGCTTGCCC	5	11	6274430_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTCCTGGTGCAGAGTGACGCTCAGGGAGGAGTTGATGGGCAGAACCAGCTCTTCATCGCGCTTGCCC;MAPQ=60;MATEID=6274430_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_16_88714501_88739501_16C;SPAN=4978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:11 DR:5 LR:-25.25 LO:27.93);ALT=G[chr16:88729418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88725128	+	chr16	88729418	+	.	6	5	6274433_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6274433_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCCC;SCTG=c_16_88714501_88739501_16C;SPAN=4290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:65 GQ:5.6 PL:[5.6, 0.0, 150.8] SR:5 DR:6 LR:-5.497 LO:13.81);ALT=C[chr16:88729418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88748302	+	chr16	88752738	+	.	8	0	6274314_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6274314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88748302(+)-16:88752738(-)__16_88739001_88764001D;SPAN=4436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=T[chr16:88752738[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88767826	+	chr16	88772577	+	.	0	17	6274252_1	45.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=6274252_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_16_88763501_88788501_24C;SPAN=4751;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:40 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:17 DR:0 LR:-45.28 LO:45.31);ALT=C[chr16:88772577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88876593	+	chr16	88878256	+	.	17	0	6275054_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6275054_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88876593(+)-16:88878256(-)__16_88861501_88886501D;SPAN=1663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:88 GQ:32.3 PL:[32.3, 0.0, 180.8] SR:0 DR:17 LR:-32.28 LO:38.24);ALT=G[chr16:88878256[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88876967	+	chr16	88878227	+	CGATGTAGTCGATGCGGCCCCCGTGGGTCGCCTTCAGGTGTCGCGCCAGGAGGCCGATGGCGGCGCGGAAGGAGGCGGGGTCCTTCAGGACGGGCGAGATGTC	120	166	6275057_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=CGATGTAGTCGATGCGGCCCCCGTGGGTCGCCTTCAGGTGTCGCGCCAGGAGGCCGATGGCGGCGCGGAAGGAGGCGGGGTCCTTCAGGACGGGCGAGATGTC;MAPQ=60;MATEID=6275057_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_88861501_88886501_194C;SPAN=1260;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:222 DP:91 GQ:59.8 PL:[656.8, 59.8, 0.0] SR:166 DR:120 LR:-656.9 LO:656.9);ALT=G[chr16:88878227[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88923634	+	chr16	88925024	+	.	40	0	6274707_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6274707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88923634(+)-16:88925024(-)__16_88910501_88935501D;SPAN=1390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:40 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:40 LR:-118.8 LO:118.8);ALT=C[chr16:88925024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88923634	+	chr16	88926070	+	.	34	0	6274708_1	96.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6274708_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:88923634(+)-16:88926070(-)__16_88910501_88935501D;SPAN=2436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:59 GQ:46.7 PL:[96.2, 0.0, 46.7] SR:0 DR:34 LR:-97.17 LO:97.17);ALT=C[chr16:88926070[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	88925199	+	chr16	88926301	+	ATACGGCTACGTCACCAACTCCAAGGTGAAGTTTGTCATGGTGGTAGATTCCTCCAACACAGCCCTTCGAGACAACGAAATTCGCAGC	0	84	6274712_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=ATACGGCTACGTCACCAACTCCAAGGTGAAGTTTGTCATGGTGGTAGATTCCTCCAACACAGCCCTTCGAGACAACGAAATTCGCAGC;MAPQ=60;MATEID=6274712_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_16_88910501_88935501_228C;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:63 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:84 DR:0 LR:-247.6 LO:247.6);ALT=T[chr16:88926301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89160405	+	chr16	89165007	+	.	8	0	6275203_1	15.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6275203_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:89160405(+)-16:89165007(-)__16_89155501_89180501D;SPAN=4602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:0 DR:8 LR:-15.03 LO:17.94);ALT=G[chr16:89165007[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89160413	+	chr16	89167068	+	.	8	0	6275204_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6275204_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:89160413(+)-16:89167068(-)__16_89155501_89180501D;SPAN=6655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=G[chr16:89167068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89574902	+	chr16	89576894	+	.	8	0	6275892_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6275892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:89574902(+)-16:89576894(-)__16_89572001_89597001D;SPAN=1992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=G[chr16:89576894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89628750	-	chr17	17286897	+	.	21	0	6332548_1	0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6332548_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:89628750(-)-17:17286897(-)__17_17272501_17297501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:21 DP:1213 GQ:99 PL:[0.0, 258.8, 3462.0] SR:0 DR:21 LR:259.3 LO:24.48);ALT=[chr17:17286897[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr16	89715907	+	chr16	89717976	+	.	2	18	6276290_1	52.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6276290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_89694501_89719501_54C;SPAN=2069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:18 DR:2 LR:-52.2 LO:52.37);ALT=T[chr16:89717976[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89715957	+	chr16	89724022	+	.	17	0	6276459_1	47.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6276459_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:89715957(+)-16:89724022(-)__16_89719001_89744001D;SPAN=8065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:32 GQ:27.8 PL:[47.6, 0.0, 27.8] SR:0 DR:17 LR:-47.65 LO:47.65);ALT=C[chr16:89724022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89718056	+	chr16	89723990	+	TCAACTGGAACAGGGTAT	0	12	6276460_1	31.0	.	EVDNC=ASSMB;INSERTION=TCAACTGGAACAGGGTAT;MAPQ=60;MATEID=6276460_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_89719001_89744001_17C;SPAN=5934;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:31 GQ:31.4 PL:[31.4, 0.0, 41.3] SR:12 DR:0 LR:-31.21 LO:31.33);ALT=T[chr16:89723990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89940267	+	chr16	89949758	+	.	26	81	6276958_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6276958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_89939501_89964501_35C;SPAN=9491;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:83 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:81 DR:26 LR:-267.4 LO:267.4);ALT=G[chr16:89949758[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89949920	+	chr16	89950988	+	.	0	8	6276987_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6276987_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_89939501_89964501_158C;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:8 DR:0 LR:-9.882 LO:16.52);ALT=G[chr16:89950988[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89951065	+	chr16	89952255	+	.	0	10	6276993_1	13.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6276993_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_89939501_89964501_114C;SPAN=1190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:73 GQ:13.4 PL:[13.4, 0.0, 161.9] SR:10 DR:0 LR:-13.23 LO:20.85);ALT=G[chr16:89952255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	89967871	+	chr16	89969134	+	.	55	19	6277041_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GAGGGGCTGTGAGGGGTGAGGGTGAAATCCCTCCTTAAGACGGGCCTCC;MAPQ=60;MATEID=6277041_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_16_89964001_89989001_53C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:13 GQ:18 PL:[198.0, 18.0, 0.0] SR:19 DR:55 LR:-198.0 LO:198.0);ALT=C[chr16:89969134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	20626	+	chr17	21729	+	.	56	0	6277629_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6277629_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:20626(+)-17:21729(-)__17_1_25001D;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:42 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:56 LR:-165.0 LO:165.0);ALT=G[chr17:21729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	193767	+	chr17	197058	+	AAATGGTTATTATT	21	17	6278713_1	89.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAATGGTTATTATT;MAPQ=60;MATEID=6278713_2;MATENM=0;NM=6;NUMPARTS=2;SCTG=c_17_196001_221001_191C;SPAN=3291;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:27 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:17 DR:21 LR:-89.12 LO:89.12);ALT=A[chr17:197058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	680259	+	chr17	685442	+	.	20	0	6279949_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6279949_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:680259(+)-17:685442(-)__17_661501_686501D;SPAN=5183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:76 GQ:45.5 PL:[45.5, 0.0, 137.9] SR:0 DR:20 LR:-45.43 LO:48.08);ALT=C[chr17:685442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	681986	+	chr17	685404	+	.	11	11	6279954_1	17.0	.	DISC_MAPQ=35;EVDNC=TSI_L;HOMSEQ=ACCT;MAPQ=60;MATEID=6279954_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_661501_686501_337C;SPAN=3418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:11 DR:11 LR:-17.4 LO:25.39);ALT=T[chr17:685404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	799035	+	chr19	6630325	+	.	2	43	6280396_1	99.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GTGAGCCGAGATCGCACCACTGCACTCCAGCCTGGG;MAPQ=60;MATEID=6280396_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_784001_809001_295C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:17 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:43 DR:2 LR:-128.7 LO:128.7);ALT=G[chr19:6630325[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr17	862402	-	chr19	5680466	+	.	35	0	6708496_1	97.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6708496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:862402(-)-19:5680466(-)__19_5659501_5684501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:67 GQ:64.4 PL:[97.4, 0.0, 64.4] SR:0 DR:35 LR:-97.72 LO:97.72);ALT=[chr19:5680466[G;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr17	900621	+	chr17	902017	+	.	0	6	6280837_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6280837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_882001_907001_2C;SPAN=1396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:73 GQ:0.2 PL:[0.2, 0.0, 175.1] SR:6 DR:0 LR:-0.02851 LO:11.1);ALT=G[chr17:902017[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1248794	+	chr17	1257503	+	.	6	4	6282185_1	15.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6282185_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_1225001_1250001_3C;SPAN=8709;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:4 DR:6 LR:-15.67 LO:21.47);ALT=C[chr17:1257503[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1257652	+	chr17	1264384	+	.	10	0	6281801_1	8.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=6281801_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1257652(+)-17:1264384(-)__17_1249501_1274501D;SPAN=6732;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:91 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:0 DR:10 LR:-8.356 LO:19.82);ALT=T[chr17:1264384[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1268383	+	chr17	1303387	+	.	97	0	6282326_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6282326_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1268383(+)-17:1303387(-)__17_1298501_1323501D;SPAN=35004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:97 DP:45 GQ:26.1 PL:[287.1, 26.1, 0.0] SR:0 DR:97 LR:-287.2 LO:287.2);ALT=C[chr17:1303387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1417319	+	chr17	1419838	+	.	11	0	6282545_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6282545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1417319(+)-17:1419838(-)__17_1396501_1421501D;SPAN=2519;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:0 DR:11 LR:-12.74 LO:22.52);ALT=A[chr17:1419838[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1585588	+	chr17	1586827	+	.	0	6	6283404_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6283404_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_1568001_1593001_179C;SPAN=1239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:82 GQ:2.1 PL:[0.0, 2.1, 201.3] SR:6 DR:0 LR:2.41 LO:10.78);ALT=C[chr17:1586827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1731301	+	chr17	1733020	+	.	7	3	6283745_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6283745_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_1715001_1740001_262C;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:3 DR:7 LR:-9.119 LO:18.15);ALT=C[chr17:1733020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1733421	+	chr17	1746096	+	.	2	3	6284044_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6284044_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_1739501_1764501_278C;SPAN=12675;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:42 GQ:5.3 PL:[5.3, 0.0, 94.4] SR:3 DR:2 LR:-5.126 LO:10.1);ALT=G[chr17:1746096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	1733462	+	chr17	1747212	+	.	14	0	6284046_1	35.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6284046_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:1733462(+)-17:1747212(-)__17_1739501_1764501D;SPAN=13750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:41 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:0 DR:14 LR:-35.11 LO:35.58);ALT=T[chr17:1747212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	2719930	+	chr17	2721218	+	.	58	42	6287557_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6287557_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_2719501_2744501_109C;SPAN=1288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:42 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:42 DR:58 LR:-237.7 LO:237.7);ALT=T[chr17:2721218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3568093	+	chr17	3571782	+	.	34	4	6289413_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6289413_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=CC;SCTG=c_17_3552501_3577501_138C;SPAN=3689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:61 GQ:46.4 PL:[99.2, 0.0, 46.4] SR:4 DR:34 LR:-99.92 LO:99.92);ALT=C[chr17:3571782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3618238	+	chr17	3619982	+	.	7	33	6290101_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6290101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_3601501_3626501_78C;SPAN=1744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:94 GQ:99 PL:[100.1, 0.0, 126.5] SR:33 DR:7 LR:-99.97 LO:100.2);ALT=T[chr17:3619982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3618278	+	chr17	3627011	+	.	13	0	6290311_1	29.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6290311_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:3618278(+)-17:3627011(-)__17_3626001_3651001D;SPAN=8733;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:49 GQ:29.6 PL:[29.6, 0.0, 89.0] SR:0 DR:13 LR:-29.64 LO:31.3);ALT=A[chr17:3627011[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3620094	+	chr17	3623601	+	.	0	68	6290108_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6290108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_3601501_3626501_344C;SPAN=3507;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:68 DP:113 GQ:78.5 PL:[194.0, 0.0, 78.5] SR:68 DR:0 LR:-196.4 LO:196.4);ALT=T[chr17:3623601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3620138	+	chr17	3627014	+	.	41	0	6290312_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6290312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:3620138(+)-17:3627014(-)__17_3626001_3651001D;SPAN=6876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:49 GQ:3.3 PL:[125.4, 3.3, 0.0] SR:0 DR:41 LR:-130.5 LO:130.5);ALT=A[chr17:3627014[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3623698	+	chr17	3626982	+	.	58	24	6290314_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6290314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_3626001_3651001_6C;SPAN=3284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:66 DP:41 GQ:17.7 PL:[194.7, 17.7, 0.0] SR:24 DR:58 LR:-194.7 LO:194.7);ALT=T[chr17:3626982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3665278	+	chr17	3667163	+	.	0	10	6290266_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6290266_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_3650501_3675501_207C;SPAN=1885;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:10 DR:0 LR:-12.69 LO:20.72);ALT=T[chr17:3667163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3667301	+	chr17	3704403	+	.	9	0	6290273_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6290273_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:3667301(+)-17:3704403(-)__17_3650501_3675501D;SPAN=37102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=G[chr17:3704403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	3743501	+	chr17	3749334	+	TGGAGGTGACATCAATTCCAGTGATGAAGCTGCCAGCCTTGTTTTCATATCTTCTGCTCGTGT	0	13	6290497_1	31.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGGAGGTGACATCAATTCCAGTGATGAAGCTGCCAGCCTTGTTTTCATATCTTCTGCTCGTGT;MAPQ=60;MATEID=6290497_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_3748501_3773501_155C;SPAN=5833;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:43 GQ:31.4 PL:[31.4, 0.0, 71.0] SR:13 DR:0 LR:-31.26 LO:32.19);ALT=T[chr17:3749334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4210421	+	chr17	4269566	+	.	0	7	6292869_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6292869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4263001_4288001_359C;SPAN=59145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:22 GQ:17.3 PL:[17.3, 0.0, 33.8] SR:7 DR:0 LR:-17.15 LO:17.52);ALT=G[chr17:4269566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4337453	+	chr17	4348239	+	.	13	0	6292534_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6292534_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:4337453(+)-17:4348239(-)__17_4336501_4361501D;SPAN=10786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:142 GQ:4.7 PL:[4.7, 0.0, 338.0] SR:0 DR:13 LR:-4.442 LO:24.68);ALT=T[chr17:4348239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4337462	+	chr17	4342948	+	.	52	102	6292535_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TGCAGG;MAPQ=60;MATEID=6292535_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_4336501_4361501_356C;SPAN=5486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:119 DP:140 GQ:14.7 PL:[369.6, 14.7, 0.0] SR:102 DR:52 LR:-381.1 LO:381.1);ALT=G[chr17:4342948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4337503	+	chr17	4349341	+	.	8	0	6292536_1	2.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6292536_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:4337503(+)-17:4349341(-)__17_4336501_4361501D;SPAN=11838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=G[chr17:4349341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4343018	+	chr17	4348326	+	.	0	39	6292557_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6292557_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4336501_4361501_164C;SPAN=5308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:109 GQ:99 PL:[99.2, 0.0, 165.2] SR:39 DR:0 LR:-99.21 LO:100.1);ALT=G[chr17:4348326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4343018	+	chr17	4349342	+	.	0	8	6292558_1	2.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6292558_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4336501_4361501_364C;SPAN=6324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:8 DR:0 LR:-1.754 LO:15.04);ALT=G[chr17:4349342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4349537	+	chr17	4351449	+	.	11	0	6292578_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6292578_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:4349537(+)-17:4351449(-)__17_4336501_4361501D;SPAN=1912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:73 GQ:16.7 PL:[16.7, 0.0, 158.6] SR:0 DR:11 LR:-16.53 LO:23.43);ALT=A[chr17:4351449[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4350259	+	chr17	4351450	+	.	3	2	6292582_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=6292582_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_4336501_4361501_152C;SPAN=1191;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:80 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:2 DR:3 LR:5.169 LO:8.632);ALT=T[chr17:4351450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4352682	+	chr17	4356308	+	.	8	6	6292591_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6292591_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4336501_4361501_110C;SPAN=3626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:95 GQ:17.3 PL:[17.3, 0.0, 212.0] SR:6 DR:8 LR:-17.18 LO:27.1);ALT=G[chr17:4356308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4389879	+	chr17	4391098	+	.	0	14	6292697_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6292697_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4385501_4410501_226C;SPAN=1219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:93 GQ:21.2 PL:[21.2, 0.0, 202.7] SR:14 DR:0 LR:-21.02 LO:29.81);ALT=G[chr17:4391098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4614040	+	chr17	4619266	+	GTCTTCAAGAAGTCGAGCCCTAACTGCA	28	18	6293606_1	83.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GTCTTCAAGAAGTCGAGCCCTAACTGCA;MAPQ=60;MATEID=6293606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4606001_4631001_30C;SPAN=5226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:82 GQ:83.6 PL:[83.6, 0.0, 113.3] SR:18 DR:28 LR:-83.42 LO:83.7);ALT=G[chr17:4619266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4614078	+	chr17	4619704	+	.	54	0	6293607_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6293607_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:4614078(+)-17:4619704(-)__17_4606001_4631001D;SPAN=5626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:96 GQ:79.7 PL:[152.3, 0.0, 79.7] SR:0 DR:54 LR:-153.4 LO:153.4);ALT=G[chr17:4619704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4844453	+	chr17	4845633	+	.	6	7	6294186_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6294186_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4826501_4851501_114C;SPAN=1180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:86 GQ:6.5 PL:[6.5, 0.0, 201.2] SR:7 DR:6 LR:-6.41 LO:17.64);ALT=G[chr17:4845633[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4850116	+	chr17	4851558	+	.	0	99	6294528_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6294528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4851001_4876001_18C;SPAN=1442;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:99 DP:223 GQ:99 PL:[266.6, 0.0, 273.2] SR:99 DR:0 LR:-266.4 LO:266.4);ALT=C[chr17:4851558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4863843	+	chr17	4871015	+	CTTTTACGAAACTCCACTTTCTGTTGTTTCTCTTGCTCTTGTAGTTTCTTCAGGCGGGCGGCCTGTT	49	23	6294571_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CTTTTACGAAACTCCACTTTCTGTTGTTTCTCTTGCTCTTGTAGTTTCTTCAGGCGGGCGGCCTGTT;MAPQ=60;MATEID=6294571_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_4851001_4876001_106C;SPAN=7172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:103 GQ:68 PL:[180.2, 0.0, 68.0] SR:23 DR:49 LR:-182.7 LO:182.7);ALT=C[chr17:4871015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	4864150	+	chr17	4871015	+	.	12	5	6294572_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6294572_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_17_4851001_4876001_106C;SPAN=6865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:81 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:5 DR:12 LR:-20.97 LO:28.08);ALT=T[chr17:4871015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5015383	+	chr17	5017452	+	.	14	0	6294835_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6294835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5015383(+)-17:5017452(-)__17_4998001_5023001D;SPAN=2069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:0 DR:14 LR:-23.73 LO:30.57);ALT=C[chr17:5017452[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5015413	+	chr17	5016681	+	.	10	9	6294837_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6294837_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_4998001_5023001_94C;SPAN=1268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:9 DR:10 LR:-19.29 LO:25.9);ALT=T[chr17:5016681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5136451	-	chr17	5137486	+	.	10	0	6295406_1	9.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6295406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5136451(-)-17:5137486(-)__17_5120501_5145501D;SPAN=1035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:0 DR:10 LR:-9.44 LO:20.03);ALT=[chr17:5137486[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	5323605	+	chr17	5324612	+	.	43	0	6296485_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6296485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5323605(+)-17:5324612(-)__17_5316501_5341501D;SPAN=1007;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:81 GQ:74 PL:[120.2, 0.0, 74.0] SR:0 DR:43 LR:-120.5 LO:120.5);ALT=C[chr17:5324612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5324786	+	chr17	5335860	+	CTGGAGGAGCTGATAGACATGGCTGTGCTGGAGGAAATTCAACAGGAGCTGATCAACCA	0	24	6296492_1	55.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CTGGAGGAGCTGATAGACATGGCTGTGCTGGAGGAAATTCAACAGGAGCTGATCAACCA;MAPQ=60;MATEID=6296492_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_5316501_5341501_72C;SPAN=11074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:87 GQ:55.7 PL:[55.7, 0.0, 154.7] SR:24 DR:0 LR:-55.65 LO:58.27);ALT=G[chr17:5335860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5384709	+	chr17	5388471	+	AGAAAAATCATGTTAAATAAAAAATTGAATCCAACTGGCCCAAAAAATAAGAAGTTGGTGATTAATCTCCATAT	0	19	6296266_1	42.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=AGAAAAATCATGTTAAATAAAAAATTGAATCCAACTGGCCCAAAAAATAAGAAGTTGGTGATTAATCTCCATAT;MAPQ=60;MATEID=6296266_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_5365501_5390501_251C;SPAN=3762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:74 GQ:42.8 PL:[42.8, 0.0, 135.2] SR:19 DR:0 LR:-42.67 LO:45.43);ALT=T[chr17:5388471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	5386244	+	chr17	5389428	+	.	8	0	6296274_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6296274_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:5386244(+)-17:5389428(-)__17_5365501_5390501D;SPAN=3184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=A[chr17:5389428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	6465014	+	chr17	6463699	+	.	30	0	6299748_1	88.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=6299748_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:6463699(-)-17:6465014(+)__17_6443501_6468501D;SPAN=1315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:40 GQ:8.9 PL:[88.1, 0.0, 8.9] SR:0 DR:30 LR:-91.98 LO:91.98);ALT=]chr17:6465014]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	6905940	+	chr17	6913115	+	.	0	9	6301151_1	16.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6301151_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_6909001_6934001_5C;SPAN=7175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:9 DR:0 LR:-16.7 LO:20.11);ALT=C[chr17:6913115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	6905974	+	chr17	6915578	+	.	13	0	6301152_1	32.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6301152_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:6905974(+)-17:6915578(-)__17_6909001_6934001D;SPAN=9604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:38 GQ:32.6 PL:[32.6, 0.0, 59.0] SR:0 DR:13 LR:-32.62 LO:33.05);ALT=A[chr17:6915578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	6918215	+	chr17	6919812	+	.	14	0	6301188_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6301188_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:6918215(+)-17:6919812(-)__17_6909001_6934001D;SPAN=1597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:0 DR:14 LR:-27.52 LO:31.83);ALT=G[chr17:6919812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7144278	+	chr17	7145471	+	.	49	0	6301878_1	99.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6301878_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7144278(+)-17:7145471(-)__17_7129501_7154501D;SPAN=1193;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:98 GQ:99 PL:[135.2, 0.0, 102.2] SR:0 DR:49 LR:-135.4 LO:135.4);ALT=A[chr17:7145471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7155915	+	chr17	7157901	+	ATTCCGTGGAGTGGGAGGGGCGCAGTCTCTTGAAGGCGCTTGTCAAGAAATCTGCACTGTGTGGGGAGCAAGTGCATATCCTGGGCTGTGAAGTGAGCGAGGAAGAGTTTCGTGAAGGTTTTGACTCTGATATCAACAATC	0	32	6301922_1	77.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=ATTCCGTGGAGTGGGAGGGGCGCAGTCTCTTGAAGGCGCTTGTCAAGAAATCTGCACTGTGTGGGGAGCAAGTGCATATCCTGGGCTGTGAAGTGAGCGAGGAAGAGTTTCGTGAAGGTTTTGACTCTGATATCAACAATC;MAPQ=60;MATEID=6301922_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_7154001_7179001_82C;SPAN=1986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:105 GQ:77.3 PL:[77.3, 0.0, 176.3] SR:32 DR:0 LR:-77.19 LO:79.37);ALT=G[chr17:7157901[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7156196	+	chr17	7157900	+	.	23	0	6301923_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6301923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7156196(+)-17:7157900(-)__17_7154001_7179001D;SPAN=1704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:85 GQ:53 PL:[53.0, 0.0, 152.0] SR:0 DR:23 LR:-52.89 LO:55.62);ALT=T[chr17:7157900[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7210470	+	chr17	7212933	+	.	17	0	6302545_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6302545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7210470(+)-17:7212933(-)__17_7203001_7228001D;SPAN=2463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:101 GQ:29 PL:[29.0, 0.0, 213.8] SR:0 DR:17 LR:-28.75 LO:37.11);ALT=G[chr17:7212933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7211075	+	chr17	7212929	+	.	111	0	6302549_1	99.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6302549_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7211075(+)-17:7212929(-)__17_7203001_7228001D;SPAN=1854;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:107 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:0 DR:111 LR:-326.8 LO:326.8);ALT=A[chr17:7212929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7211432	+	chr17	7212932	+	.	51	7	6302550_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6302550_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_7203001_7228001_234C;SPAN=1500;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:108 GQ:99 PL:[149.0, 0.0, 112.7] SR:7 DR:51 LR:-149.3 LO:149.3);ALT=G[chr17:7212932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7240106	+	chr17	7245265	+	AGCCTCTATTGAGCTGGTGGAAGCCGAAGTGTCAGAATTGGAGACCCGTCTGGAAA	12	40	6302035_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGCCTCTATTGAGCTGGTGGAAGCCGAAGTGTCAGAATTGGAGACCCGTCTGGAAA;MAPQ=60;MATEID=6302035_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_7227501_7252501_94C;SPAN=5159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:96 GQ:99 PL:[125.9, 0.0, 106.1] SR:40 DR:12 LR:-125.9 LO:125.9);ALT=G[chr17:7245265[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7253557	+	chr17	7254611	+	CTACGACTGGCAAAGATGAGGGAGGCTGAAGCGGCCCAGGGGCAGG	0	47	6302187_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CTACGACTGGCAAAGATGAGGGAGGCTGAAGCGGCCCAGGGGCAGG;MAPQ=60;MATEID=6302187_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_7252001_7277001_290C;SPAN=1054;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:84 GQ:69.8 PL:[132.5, 0.0, 69.8] SR:47 DR:0 LR:-133.4 LO:133.4);ALT=G[chr17:7254611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7264613	+	chr17	7265990	+	.	14	7	6302223_1	47.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=TGCCTGCAGTCCCAGCTACTCAGGAGGCTGAGGTG;MAPQ=39;MATEID=6302223_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_7252001_7277001_218C;SPAN=1377;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:68 GQ:47.6 PL:[47.6, 0.0, 116.9] SR:7 DR:14 LR:-47.6 LO:49.23);ALT=G[chr17:7265990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7336437	+	chr17	7337683	+	.	44	0	6302286_1	99.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6302286_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7336437(+)-17:7337683(-)__17_7325501_7350501D;SPAN=1246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:30 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:0 DR:44 LR:-128.7 LO:128.7);ALT=C[chr17:7337683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7487261	+	chr17	7489258	+	.	23	0	6303021_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6303021_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7487261(+)-17:7489258(-)__17_7472501_7497501D;SPAN=1997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:86 GQ:52.7 PL:[52.7, 0.0, 155.0] SR:0 DR:23 LR:-52.62 LO:55.48);ALT=C[chr17:7489258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7487261	+	chr17	7489013	+	.	8	0	6303020_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6303020_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7487261(+)-17:7489013(-)__17_7472501_7497501D;SPAN=1752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:0 DR:8 LR:-0.6702 LO:14.89);ALT=C[chr17:7489013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7579941	+	chr17	7590695	+	.	7	4	6303595_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6303595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_7570501_7595501_155C;SPAN=10754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:87 GQ:12.8 PL:[12.8, 0.0, 197.6] SR:4 DR:7 LR:-12.74 LO:22.52);ALT=C[chr17:7590695[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7788401	+	chr17	7792980	+	.	6	12	6304260_1	30.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6304260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_7791001_7816001_12C;SPAN=4579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:12 DR:6 LR:-30.18 LO:31.58);ALT=G[chr17:7792980[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	7798847	+	chr17	7800398	+	.	8	0	6304276_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6304276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:7798847(+)-17:7800398(-)__17_7791001_7816001D;SPAN=1551;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=C[chr17:7800398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8065086	+	chr17	8066194	+	CATCCACCTGGGCCTGGGTCTGCTGCAGTCTCCTGTTACTGGTGAGGTTTGGAGGGGGTGCAGGGGGACCACCCTCCCCAGCCGGGGCAGCAGGGGGGGCCGTGGCAGCGGTAGCAG	81	92	6305596_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=CATCCACCTGGGCCTGGGTCTGCTGCAGTCTCCTGTTACTGGTGAGGTTTGGAGGGGGTGCAGGGGGACCACCCTCCCCAGCCGGGGCAGCAGGGGGGGCCGTGGCAGCGGTAGCAG;MAPQ=60;MATEID=6305596_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_8060501_8085501_71C;SPAN=1108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:132 DP:107 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:92 DR:81 LR:-389.5 LO:389.5);ALT=T[chr17:8066194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8111210	+	chr17	8113847	+	.	11	0	6305214_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6305214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:8111210(+)-17:8113847(-)__17_8109501_8134501D;SPAN=2637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:112 GQ:6.2 PL:[6.2, 0.0, 263.6] SR:0 DR:11 LR:-5.968 LO:21.24);ALT=G[chr17:8113847[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8246645	+	chr17	8247969	+	.	63	11	6306144_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=GCTAATTTTTGTATTTTTAGTAGAGACGGGGTTT;MAPQ=60;MATEID=6306144_2;MATENM=0;NM=4;NUMPARTS=2;SCTG=c_17_8232001_8257001_352C;SPAN=1324;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:37 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:11 DR:63 LR:-208.0 LO:208.0);ALT=T[chr17:8247969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	8631471	+	chr19	35976906	-	.	12	20	6307100_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TGGGTGGGTGGATGG;MAPQ=60;MATEID=6307100_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_8624001_8649001_224C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:28 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:20 DR:12 LR:-82.01 LO:82.01);ALT=A]chr19:35976906];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr17	8814829	+	chr17	8868912	+	.	4	2	6307850_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTGCA;MAPQ=60;MATEID=6307850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_8869001_8894001_277C;SPAN=54083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:4 DP:1 GQ:0.9 PL:[9.9, 0.9, 0.0] SR:2 DR:4 LR:-9.903 LO:9.903);ALT=A[chr17:8868912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	9448599	+	chr17	9460751	+	.	0	28	6309649_1	79.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6309649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_9457001_9482001_187C;SPAN=12152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:47 GQ:33.5 PL:[79.7, 0.0, 33.5] SR:28 DR:0 LR:-80.67 LO:80.67);ALT=T[chr17:9460751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	9448649	+	chr17	9471687	+	.	11	0	6309650_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6309650_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:9448649(+)-17:9471687(-)__17_9457001_9482001D;SPAN=23038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:40 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:0 DR:11 LR:-25.47 LO:26.69);ALT=A[chr17:9471687[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	9460847	+	chr17	9471688	+	.	31	24	6309664_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6309664_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_9457001_9482001_247C;SPAN=10841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:90 GQ:99 PL:[110.9, 0.0, 107.6] SR:24 DR:31 LR:-111.0 LO:111.0);ALT=T[chr17:9471688[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	9460887	+	chr17	9479106	+	.	11	0	6309665_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6309665_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:9460887(+)-17:9479106(-)__17_9457001_9482001D;SPAN=18219;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:0 DR:11 LR:-10.84 LO:22.13);ALT=T[chr17:9479106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	20541255	+	chr17	15723274	+	.	16	0	6327132_1	33.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6327132_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:15723274(-)-17:20541255(+)__17_15704501_15729501D;SPAN=4817981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:73 GQ:33.2 PL:[33.2, 0.0, 142.1] SR:0 DR:16 LR:-33.04 LO:36.98);ALT=]chr17:20541255]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	15723555	+	chr17	20541424	+	.	16	0	6327134_1	36.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6327134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:15723555(+)-17:20541424(-)__17_15704501_15729501D;SPAN=4817869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:61 GQ:36.5 PL:[36.5, 0.0, 109.1] SR:0 DR:16 LR:-36.29 LO:38.43);ALT=A[chr17:20541424[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	15881478	+	chr17	15884354	+	.	0	9	6327710_1	7.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6327710_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_15876001_15901001_130C;SPAN=2876;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:82 GQ:7.7 PL:[7.7, 0.0, 189.2] SR:9 DR:0 LR:-7.493 LO:17.84);ALT=C[chr17:15884354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	15884507	+	chr17	15902863	+	.	9	0	6327724_1	20.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6327724_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:15884507(+)-17:15902863(-)__17_15876001_15901001D;SPAN=18356;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=C[chr17:15902863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	15890682	+	chr17	15902833	+	GATAACAGATATTCATCAGGAA	0	38	6327750_1	99.0	.	EVDNC=ASSMB;INSERTION=GATAACAGATATTCATCAGGAA;MAPQ=60;MATEID=6327750_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_15876001_15901001_82C;SPAN=12151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:45 GQ:5.4 PL:[118.8, 5.4, 0.0] SR:38 DR:0 LR:-121.4 LO:121.4);ALT=C[chr17:15902833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	15905339	+	chr17	15907512	+	ATGGCCAACTTAGCATTTATACGGGGTCAGCTTGAAAATGCTGAACAACTTTTTAAAGCAACAATGAGTTACCTCCTTGGAGGGGGCATGAAG	0	12	6327426_1	15.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=ATGGCCAACTTAGCATTTATACGGGGTCAGCTTGAAAATGCTGAACAACTTTTTAAAGCAACAATGAGTTACCTCCTTGGAGGGGGCATGAAG;MAPQ=60;MATEID=6327426_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_15900501_15925501_245C;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:12 DR:0 LR:-15.23 LO:24.87);ALT=G[chr17:15907512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16042502	+	chr17	16046920	+	.	5	2	6327934_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6327934_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_16023001_16048001_363C;SPAN=4418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:76 GQ:0.6 PL:[0.0, 0.6, 184.8] SR:2 DR:5 LR:0.7843 LO:10.99);ALT=T[chr17:16046920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16097996	+	chr17	16118783	+	.	26	0	6328601_1	66.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6328601_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:16097996(+)-17:16118783(-)__17_16096501_16121501D;SPAN=20787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:73 GQ:66.2 PL:[66.2, 0.0, 109.1] SR:0 DR:26 LR:-66.05 LO:66.68);ALT=C[chr17:16118783[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16102061	+	chr17	16118787	+	.	9	0	6328620_1	8.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6328620_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:16102061(+)-17:16118787(-)__17_16096501_16121501D;SPAN=16726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:0 DR:9 LR:-8.306 LO:17.99);ALT=T[chr17:16118787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16319190	+	chr17	16320874	+	.	17	0	6329040_1	35.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6329040_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:16319190(+)-17:16320874(-)__17_16317001_16342001D;SPAN=1684;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:75 GQ:35.9 PL:[35.9, 0.0, 144.8] SR:0 DR:17 LR:-35.8 LO:39.58);ALT=T[chr17:16320874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16342722	+	chr17	16344679	+	.	25	0	6329155_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6329155_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:16342722(+)-17:16344679(-)__17_16341501_16366501D;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:25 DP:336 GQ:8.3 PL:[0.0, 8.3, 831.8] SR:0 DR:25 LR:8.506 LO:45.12);ALT=G[chr17:16344679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	16343569	+	chr17	16344680	+	.	15	11	6329169_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6329169_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_16341501_16366501_239C;SPAN=1111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:26 DP:441 GQ:33.3 PL:[0.0, 33.3, 1135.0] SR:11 DR:15 LR:33.65 LO:44.21);ALT=T[chr17:16344680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	17163790	+	chr17	17165280	+	.	5	2	6332134_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6332134_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_17150001_17175001_139C;SPAN=1490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:82 GQ:2.1 PL:[0.0, 2.1, 201.3] SR:2 DR:5 LR:2.41 LO:10.78);ALT=T[chr17:17165280[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	17174370	+	chr17	17184450	+	.	21	0	6332276_1	56.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6332276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:17174370(+)-17:17184450(-)__17_17174501_17199501D;SPAN=10080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:46 GQ:53.6 PL:[56.9, 0.0, 53.6] SR:0 DR:21 LR:-56.86 LO:56.86);ALT=A[chr17:17184450[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	17179480	+	chr17	17184445	+	.	0	15	6332297_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6332297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_17174501_17199501_388C;SPAN=4965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:95 GQ:23.9 PL:[23.9, 0.0, 205.4] SR:15 DR:0 LR:-23.78 LO:32.28);ALT=T[chr17:17184445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	17480344	+	chr17	17494844	+	.	23	12	6333135_1	80.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6333135_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_17493001_17518001_279C;SPAN=14500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:46 GQ:30.5 PL:[80.0, 0.0, 30.5] SR:12 DR:23 LR:-81.11 LO:81.11);ALT=G[chr17:17494844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	17991401	+	chr17	17997126	+	.	18	4	6334973_1	46.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6334973_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_17983001_18008001_379C;SPAN=5725;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:72 GQ:46.7 PL:[46.7, 0.0, 125.9] SR:4 DR:18 LR:-46.51 LO:48.63);ALT=G[chr17:17997126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	18007995	+	chr17	18010467	+	TGCCACCGCATCCACCGGTCACTCGCCAGCCAGTTCAAGTACGCCCTGGTGTG	0	10	6334540_1	8.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=TGCCACCGCATCCACCGGTCACTCGCCAGCCAGTTCAAGTACGCCCTGGTGTG;MAPQ=60;MATEID=6334540_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_18007501_18032501_111C;SPAN=2472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:10 DR:0 LR:-8.627 LO:19.88);ALT=G[chr17:18010467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	18160335	+	chr17	18161941	+	.	8	1	6335154_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6335154_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_18154501_18179501_307C;SPAN=1606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:1 DR:8 LR:-8.256 LO:16.17);ALT=T[chr17:18161941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	18761560	+	chr17	18769112	+	.	9	0	6337678_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6337678_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:18761560(+)-17:18769112(-)__17_18767001_18792001D;SPAN=7552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:0 DR:9 LR:-21.04 LO:21.94);ALT=T[chr17:18769112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	18761575	+	chr17	18768778	+	.	6	3	6337679_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAGG;MAPQ=60;MATEID=6337679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_18767001_18792001_101C;SPAN=7203;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:35 GQ:10.4 PL:[10.4, 0.0, 73.1] SR:3 DR:6 LR:-10.32 LO:13.15);ALT=G[chr17:18768778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	19977050	+	chr17	19999946	+	.	12	0	6342399_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6342399_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:19977050(+)-17:19999946(-)__17_19992001_20017001D;SPAN=22896;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:45 GQ:27.5 PL:[27.5, 0.0, 80.3] SR:0 DR:12 LR:-27.42 LO:28.93);ALT=T[chr17:19999946[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	20000111	+	chr17	20013739	+	.	0	10	6342428_1	6.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6342428_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_19992001_20017001_294C;SPAN=13628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:97 GQ:6.8 PL:[6.8, 0.0, 227.9] SR:10 DR:0 LR:-6.73 LO:19.53);ALT=G[chr17:20013739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	21102128	+	chr17	21117412	+	.	21	0	6345815_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6345815_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:21102128(+)-17:21117412(-)__17_21094501_21119501D;SPAN=15284;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:79 GQ:47.9 PL:[47.9, 0.0, 143.6] SR:0 DR:21 LR:-47.92 LO:50.59);ALT=A[chr17:21117412[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	22071212	+	chr17	22069912	+	.	12	0	6348713_1	21.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6348713_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:22069912(-)-17:22071212(+)__17_22050001_22075001D;SPAN=1300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:0 DR:12 LR:-21.73 LO:26.64);ALT=]chr17:22071212]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	25536553	+	chr17	25540382	+	.	38	22	6349875_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAATTCACATGGCA;MAPQ=60;MATEID=6349875_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25529001_25554001_137C;SPAN=3829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:92 GQ:71 PL:[150.2, 0.0, 71.0] SR:22 DR:38 LR:-151.5 LO:151.5);ALT=A[chr17:25540382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25621461	+	chr17	25628821	+	TGAGATC	0	10	6350423_1	20.0	.	EVDNC=ASSMB;INSERTION=TGAGATC;MAPQ=60;MATEID=6350423_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25627001_25652001_13C;SPAN=7360;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:10 DR:0 LR:-20.82 LO:23.18);ALT=G[chr17:25628821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25628982	+	chr17	25630393	+	.	2	3	6350435_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6350435_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_25627001_25652001_214C;SPAN=1411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:82 GQ:8.7 PL:[0.0, 8.7, 214.5] SR:3 DR:2 LR:9.012 LO:6.465);ALT=T[chr17:25630393[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25958358	+	chr17	25967595	+	.	89	0	6351234_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6351234_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:25958358(+)-17:25967595(-)__17_25945501_25970501D;SPAN=9237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:89 DP:75 GQ:24 PL:[264.0, 24.0, 0.0] SR:0 DR:89 LR:-264.1 LO:264.1);ALT=C[chr17:25967595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25974146	+	chr17	25975862	+	TCCACATCAACCTGTGCTCTGGGAACCACATCGCCTTCCACCTGAACCCCCGTTTTGATGAGAATGCTGTGGTCCGCAACACCCAGATCGACAACTCCTGGGGGTCTGAGGAGCGAAGTCTGCCCCGAAAAATGCCCTTCGTCCGTGGCCAGAGCTTCTCA	2	12	6351307_1	20.0	.	DISC_MAPQ=28;EVDNC=TSI_G;HOMSEQ=GT;INSERTION=TCCACATCAACCTGTGCTCTGGGAACCACATCGCCTTCCACCTGAACCCCCGTTTTGATGAGAATGCTGTGGTCCGCAACACCCAGATCGACAACTCCTGGGGGTCTGAGGAGCGAAGTCTGCCCCGAAAAATGCCCTTCGTCCGTGGCCAGAGCTTCTCA;MAPQ=28;MATEID=6351307_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_25970001_25995001_223C;SPAN=1716;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:82 GQ:20.9 PL:[20.9, 0.0, 176.0] SR:12 DR:2 LR:-20.7 LO:28.0);ALT=T[chr17:25975862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25974460	+	chr17	25975862	+	.	8	7	6351309_1	15.0	.	DISC_MAPQ=44;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=6351309_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_25970001_25995001_223C;SPAN=1402;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:7 DR:8 LR:-15.23 LO:24.87);ALT=T[chr17:25975862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	25982467	+	chr17	26087797	+	.	9	0	6351333_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6351333_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:25982467(+)-17:26087797(-)__17_25970001_25995001D;SPAN=105330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:0 DR:9 LR:-21.04 LO:21.94);ALT=G[chr17:26087797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26594299	+	chr17	26592913	+	.	8	10	6352951_1	39.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=TTCTTTGCCCTGCCTCTCGACCCTTTTTGTC;MAPQ=59;MATEID=6352951_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_26582501_26607501_192C;SPAN=1386;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:75 GQ:39.2 PL:[39.2, 0.0, 141.5] SR:10 DR:8 LR:-39.1 LO:42.43);ALT=]chr17:26594299]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	26657554	+	chr17	26658885	+	.	0	13	6353243_1	21.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6353243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_26656001_26681001_333C;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:80 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:13 DR:0 LR:-21.24 LO:28.16);ALT=T[chr17:26658885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26659037	+	chr17	26662385	+	.	15	0	6353248_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6353248_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:26659037(+)-17:26662385(-)__17_26656001_26681001D;SPAN=3348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:78 GQ:28.4 PL:[28.4, 0.0, 160.4] SR:0 DR:15 LR:-28.38 LO:33.71);ALT=C[chr17:26662385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26681614	+	chr17	26682821	+	.	0	6	6353380_1	0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6353380_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_26680501_26705501_127C;SPAN=1207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:74 GQ:0 PL:[0.0, 0.0, 178.2] SR:6 DR:0 LR:0.2424 LO:11.06);ALT=G[chr17:26682821[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26682903	+	chr17	26684314	+	.	0	14	6353385_1	27.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6353385_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_26680501_26705501_311C;SPAN=1411;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:69 GQ:27.5 PL:[27.5, 0.0, 139.7] SR:14 DR:0 LR:-27.52 LO:31.83);ALT=C[chr17:26684314[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26684904	+	chr17	26685938	+	.	0	9	6353396_1	8.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6353396_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_26680501_26705501_76C;SPAN=1034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-7.764 LO:17.89);ALT=G[chr17:26685938[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26982521	+	chr17	26988761	+	.	11	0	6354301_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6354301_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:26982521(+)-17:26988761(-)__17_26974501_26999501D;SPAN=6240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:95 GQ:10.7 PL:[10.7, 0.0, 218.6] SR:0 DR:11 LR:-10.57 LO:22.07);ALT=G[chr17:26988761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26989360	+	chr17	27000392	+	TTG	7	1	6354457_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TTG;MAPQ=60;MATEID=6354457_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_26999001_27024001_346C;SPAN=11032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:1 DR:7 LR:-9.832 LO:14.73);ALT=G[chr17:27000392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	26989372	+	chr17	26997587	+	.	15	0	6354332_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6354332_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:26989372(+)-17:26997587(-)__17_26974501_26999501D;SPAN=8215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:86 GQ:26.3 PL:[26.3, 0.0, 181.4] SR:0 DR:15 LR:-26.22 LO:33.0);ALT=A[chr17:26997587[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27044052	+	chr17	27045138	+	.	9	0	6354428_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6354428_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:27044052(+)-17:27045138(-)__17_27023501_27048501D;SPAN=1086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=C[chr17:27045138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27210252	+	chr17	27215962	+	GGCGACACCCGTCACAGTTAAAGCTACCCCCTCGGCCGTCTCTACGTCCTCGCAGCGGGGCTGCAACGTCATAATCTCTAGGGAAAT	0	39	6355101_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GGCGACACCCGTCACAGTTAAAGCTACCCCCTCGGCCGTCTCTACGTCCTCGCAGCGGGGCTGCAACGTCATAATCTCTAGGGAAAT;MAPQ=60;MATEID=6355101_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_27195001_27220001_361C;SPAN=5710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:88 GQ:99 PL:[104.9, 0.0, 108.2] SR:39 DR:0 LR:-104.9 LO:104.9);ALT=G[chr17:27215962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27211381	+	chr17	27224591	+	.	17	0	6355105_1	45.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6355105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:27211381(+)-17:27224591(-)__17_27195001_27220001D;SPAN=13210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:0 DR:17 LR:-45.01 LO:45.06);ALT=T[chr17:27224591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27216047	+	chr17	27224543	+	.	32	19	6355115_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6355115_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_27195001_27220001_204C;SPAN=8496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:19 DR:32 LR:-112.2 LO:112.2);ALT=G[chr17:27224543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27685161	-	chr17	27686697	+	.	8	0	6356757_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6356757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:27685161(-)-17:27686697(-)__17_27685001_27710001D;SPAN=1536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:97 GQ:0.2 PL:[0.2, 0.0, 234.5] SR:0 DR:8 LR:-0.1283 LO:14.81);ALT=[chr17:27686697[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	27895836	+	chr17	27898605	+	.	11	0	6357254_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6357254_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:27895836(+)-17:27898605(-)__17_27881001_27906001D;SPAN=2769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:62 GQ:19.7 PL:[19.7, 0.0, 128.6] SR:0 DR:11 LR:-19.51 LO:24.29);ALT=G[chr17:27898605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	27896106	+	chr17	27898606	+	GTCACCAAGAGTGACCTACACACGAGTGAGCCCAGGG	0	23	6357258_1	49.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=GTCACCAAGAGTGACCTACACACGAGTGAGCCCAGGG;MAPQ=60;MATEID=6357258_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_27881001_27906001_27C;SPAN=2500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:98 GQ:49.4 PL:[49.4, 0.0, 188.0] SR:23 DR:0 LR:-49.37 LO:53.95);ALT=T[chr17:27898606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	28252574	+	chr17	28256956	+	.	0	17	6358696_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6358696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_28248501_28273501_221C;SPAN=4382;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:99 GQ:29.3 PL:[29.3, 0.0, 210.8] SR:17 DR:0 LR:-29.3 LO:37.27);ALT=C[chr17:28256956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29045669	+	chr19	14307742	+	.	0	7	6741090_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCTGGC;MAPQ=60;MATEID=6741090_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14283501_14308501_430C;SPAN=-1;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:37 GQ:13.1 PL:[13.1, 0.0, 75.8] SR:7 DR:0 LR:-13.08 LO:15.67);ALT=C[chr19:14307742[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr17	29131151	+	chr17	29151589	+	.	11	0	6361920_1	29.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6361920_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:29131151(+)-17:29151589(-)__17_29106001_29131001D;SPAN=20438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:0 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:11 LR:-29.71 LO:29.71);ALT=A[chr17:29151589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29231570	+	chr17	29233185	+	.	9	0	6362080_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6362080_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:29231570(+)-17:29233185(-)__17_29228501_29253501D;SPAN=1615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:77 GQ:8.9 PL:[8.9, 0.0, 177.2] SR:0 DR:9 LR:-8.848 LO:18.1);ALT=T[chr17:29233185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29632650	+	chr17	29640997	+	.	94	5	6363310_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6363310_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_29620501_29645501_208C;SPAN=8347;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:93 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:5 DR:94 LR:-277.3 LO:277.3);ALT=T[chr17:29640997[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	29646043	+	chr17	29648513	+	.	10	2	6363547_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6363547_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_29645001_29670001_273C;SPAN=2470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:2 DR:10 LR:-13.55 LO:22.7);ALT=T[chr17:29648513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30180096	+	chr17	30186174	+	.	8	0	6365084_1	20.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6365084_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:30180096(+)-17:30186174(-)__17_30184001_30209001D;SPAN=6078;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:0 DR:8 LR:-19.91 LO:20.23);ALT=C[chr17:30186174[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30190536	+	chr17	30192385	+	.	3	2	6365102_1	0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6365102_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30184001_30209001_36C;SPAN=1849;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:68 GQ:5.1 PL:[0.0, 5.1, 174.9] SR:2 DR:3 LR:5.219 LO:6.798);ALT=C[chr17:30192385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30226749	+	chr17	30228554	+	.	8	9	6365261_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6365261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30208501_30233501_62C;SPAN=1805;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:84 GQ:20.3 PL:[20.3, 0.0, 182.0] SR:9 DR:8 LR:-20.16 LO:27.85);ALT=C[chr17:30228554[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30666959	+	chr17	30668223	+	.	0	5	6366754_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6366754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30649501_30674501_238C;SPAN=1264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:5 DR:0 LR:5.711 LO:8.577);ALT=T[chr17:30668223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30677349	+	chr17	30678804	+	.	33	44	6366796_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTAT;MAPQ=60;MATEID=6366796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30674001_30699001_163C;SECONDARY;SPAN=1455;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:92 GQ:11.6 PL:[209.6, 0.0, 11.6] SR:44 DR:33 LR:-219.6 LO:219.6);ALT=T[chr17:30678804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30771611	+	chr17	30781509	+	.	9	0	6367367_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6367367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:30771611(+)-17:30781509(-)__17_30772001_30797001D;SPAN=9898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:0 DR:9 LR:-14.54 LO:19.45);ALT=A[chr17:30781509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30771632	+	chr17	30773962	+	.	25	10	6367368_1	71.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6367368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30772001_30797001_300C;SPAN=2330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:53 GQ:55.1 PL:[71.6, 0.0, 55.1] SR:10 DR:25 LR:-71.55 LO:71.55);ALT=G[chr17:30773962[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	30774064	+	chr17	30781510	+	.	0	17	6367376_1	29.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6367376_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_30772001_30797001_314C;SPAN=7446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:100 GQ:29 PL:[29.0, 0.0, 213.8] SR:17 DR:0 LR:-29.02 LO:37.19);ALT=G[chr17:30781510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	33307679	+	chr17	33310086	+	.	8	0	6374433_1	8.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6374433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:33307679(+)-17:33310086(-)__17_33295501_33320501D;SPAN=2407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:65 GQ:8.9 PL:[8.9, 0.0, 147.5] SR:0 DR:8 LR:-8.798 LO:16.28);ALT=C[chr17:33310086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	33467088	+	chr17	33468997	+	.	0	9	6374472_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=6374472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_33467001_33492001_107C;SPAN=1909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-8.035 LO:17.94);ALT=G[chr17:33468997[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	33467129	+	chr17	33469279	+	.	12	0	6374473_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6374473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:33467129(+)-17:33469279(-)__17_33467001_33492001D;SPAN=2150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:88 GQ:15.8 PL:[15.8, 0.0, 197.3] SR:0 DR:12 LR:-15.77 LO:24.99);ALT=C[chr17:33469279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	33862367	-	chr17	33863569	+	.	12	0	6375531_1	19.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6375531_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:33862367(-)-17:33863569(-)__17_33859001_33884001D;SPAN=1202;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:75 GQ:19.4 PL:[19.4, 0.0, 161.3] SR:0 DR:12 LR:-19.29 LO:25.9);ALT=[chr17:33863569[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	33914450	+	chr17	33921026	+	.	11	4	6376198_1	18.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6376198_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_33908001_33933001_55C;SPAN=6576;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:89 GQ:18.8 PL:[18.8, 0.0, 197.0] SR:4 DR:11 LR:-18.8 LO:27.5);ALT=G[chr17:33921026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34136580	+	chr17	34144719	+	.	3	9	6376452_1	5.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6376452_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_17_34128501_34153501_237C;SPAN=8139;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:9 DR:3 LR:-5.868 LO:17.54);ALT=G[chr17:34144719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34136609	+	chr17	34147025	+	.	71	0	6376454_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6376454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34136609(+)-17:34147025(-)__17_34128501_34153501D;SPAN=10416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:89 GQ:5.6 PL:[210.2, 0.0, 5.6] SR:0 DR:71 LR:-222.0 LO:222.0);ALT=A[chr17:34147025[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34147441	+	chr17	34151080	+	CCAAGGTGGAAGAGCACCTTCCTATGACCAGCCAGACTATGGTCAACAAGATTCATATGACCAGCAGTCAGGCTATGATCAACATCAAGGCTCATATGATGAGCAGTCAAATTATGATCAGCAGCATGATTCCTATAGTCAAAACCAGCAGTCCTATCATTCACAAAGGGAAAACTACAGCCACCACACACA	3	20	6376486_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCAAGGTGGAAGAGCACCTTCCTATGACCAGCCAGACTATGGTCAACAAGATTCATATGACCAGCAGTCAGGCTATGATCAACATCAAGGCTCATATGATGAGCAGTCAAATTATGATCAGCAGCATGATTCCTATAGTCAAAACCAGCAGTCCTATCATTCACAAAGGGAAAACTACAGCCACCACACACA;MAPQ=60;MATEID=6376486_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_34128501_34153501_44C;SPAN=3639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:91 GQ:44.9 PL:[44.9, 0.0, 173.6] SR:20 DR:3 LR:-44.67 LO:49.08);ALT=G[chr17:34151080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34149837	+	chr17	34151080	+	.	11	15	6376502_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6376502_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_34128501_34153501_44C;SPAN=1243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:87 GQ:45.8 PL:[45.8, 0.0, 164.6] SR:15 DR:11 LR:-45.75 LO:49.56);ALT=G[chr17:34151080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34165558	+	chr17	34171079	+	AAAAGAATTCCATGGCAACATCATTAAAGTGTCCTTTGCCACTAGAAGACCTGAATTCATGAGAGGAGGTGGAAGTGGAGGTGGGCGGCG	0	10	6376589_1	7.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAAAGAATTCCATGGCAACATCATTAAAGTGTCCTTTGCCACTAGAAGACCTGAATTCATGAGAGGAGGTGGAAGTGGAGGTGGGCGGCG;MAPQ=60;MATEID=6376589_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_34153001_34178001_356C;SPAN=5521;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:10 DR:0 LR:-7.272 LO:19.63);ALT=G[chr17:34171079[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34165558	+	chr17	34169370	+	.	2	5	6376588_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6376588_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAA;SCTG=c_17_34153001_34178001_356C;SPAN=3812;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:75 GQ:0.3 PL:[0.0, 0.3, 181.5] SR:5 DR:2 LR:0.5133 LO:11.02);ALT=G[chr17:34169370[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34172042	+	chr17	34173908	+	.	16	17	6376613_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6376613_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_34153001_34178001_65C;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:108 GQ:53.3 PL:[53.3, 0.0, 208.4] SR:17 DR:16 LR:-53.27 LO:58.47);ALT=G[chr17:34173908[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34199468	+	chr17	34205532	+	.	7	36	6376742_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6376742_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_17_34202001_34227001_348C;SPAN=6064;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:50 GQ:3.6 PL:[128.7, 3.6, 0.0] SR:36 DR:7 LR:-133.8 LO:133.8);ALT=G[chr17:34205532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34199515	+	chr17	34207233	+	.	25	0	6376743_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6376743_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34199515(+)-17:34207233(-)__17_34202001_34227001D;SPAN=7718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:49 GQ:49.4 PL:[69.2, 0.0, 49.4] SR:0 DR:25 LR:-69.42 LO:69.42);ALT=G[chr17:34207233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34205643	+	chr17	34207234	+	.	48	22	6376754_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6376754_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_34202001_34227001_212C;SPAN=1591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:106 GQ:93.5 PL:[162.8, 0.0, 93.5] SR:22 DR:48 LR:-163.7 LO:163.7);ALT=T[chr17:34207234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34340998	+	chr17	34344894	+	.	13	0	6377160_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6377160_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34340998(+)-17:34344894(-)__17_34324501_34349501D;SPAN=3896;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:76 GQ:22.4 PL:[22.4, 0.0, 161.0] SR:0 DR:13 LR:-22.32 LO:28.48);ALT=C[chr17:34344894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34341479	+	chr17	34344932	+	.	14	0	6377162_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6377162_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34341479(+)-17:34344932(-)__17_34324501_34349501D;SPAN=3453;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:78 GQ:25.1 PL:[25.1, 0.0, 163.7] SR:0 DR:14 LR:-25.08 LO:30.99);ALT=C[chr17:34344932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34416157	+	chr17	34417331	+	.	49	0	6377628_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6377628_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:34416157(+)-17:34417331(-)__17_34398001_34423001D;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:94 GQ:90.2 PL:[136.4, 0.0, 90.2] SR:0 DR:49 LR:-136.7 LO:136.7);ALT=A[chr17:34417331[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34842629	+	chr17	34848655	+	CTGCTCGGTAGTCTGCTTCCGGAAGCACAA	15	9	6378524_1	71.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGCTCGGTAGTCTGCTTCCGGAAGCACAA;MAPQ=60;MATEID=6378524_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_34839001_34864001_176C;SPAN=6026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:104 GQ:71 PL:[71.0, 0.0, 179.9] SR:9 DR:15 LR:-70.85 LO:73.54);ALT=A[chr17:34848655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	34935849	+	chr17	34937772	+	.	4	7	6379179_1	21.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6379179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_34937001_34962001_224C;SPAN=1923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:7 DR:4 LR:-21.04 LO:21.94);ALT=G[chr17:34937772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	35307705	+	chr17	35310185	+	.	5	2	6380312_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6380312_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_35304501_35329501_61C;SPAN=2480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:71 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:2 DR:5 LR:-3.871 LO:13.53);ALT=G[chr17:35310185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	35946659	+	chr17	35956269	+	.	0	7	6382295_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6382295_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_35941501_35966501_248C;SPAN=9610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.547 LO:12.74);ALT=T[chr17:35956269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	35956448	+	chr17	35969383	+	.	8	0	6382580_1	13.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6382580_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:35956448(+)-17:35969383(-)__17_35966001_35991001D;SPAN=12935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:47 GQ:13.7 PL:[13.7, 0.0, 99.5] SR:0 DR:8 LR:-13.67 LO:17.51);ALT=A[chr17:35969383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36002339	+	chr17	36003363	+	.	0	5	6382382_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6382382_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_35990501_36015501_61C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:74 GQ:3.3 PL:[0.0, 3.3, 184.8] SR:5 DR:0 LR:3.543 LO:8.807);ALT=T[chr17:36003363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36453222	+	chr17	36455311	+	.	10	0	6384636_1	12.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=6384636_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:36453222(+)-17:36455311(-)__17_36431501_36456501D;SPAN=2089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:75 GQ:12.8 PL:[12.8, 0.0, 167.9] SR:0 DR:10 LR:-12.69 LO:20.72);ALT=A[chr17:36455311[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36886695	+	chr17	36889525	+	.	16	0	6386214_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6386214_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:36886695(+)-17:36889525(-)__17_36872501_36897501D;SPAN=2830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:69 GQ:34.1 PL:[34.1, 0.0, 133.1] SR:0 DR:16 LR:-34.12 LO:37.43);ALT=A[chr17:36889525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36887692	+	chr17	36889526	+	.	0	17	6386218_1	33.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6386218_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36872501_36897501_275C;SPAN=1834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:85 GQ:33.2 PL:[33.2, 0.0, 171.8] SR:17 DR:0 LR:-33.09 LO:38.53);ALT=G[chr17:36889526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36909128	+	chr17	36912134	+	.	20	0	6386448_1	41.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6386448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:36909128(+)-17:36912134(-)__17_36897001_36922001D;SPAN=3006;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:90 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:0 DR:20 LR:-41.64 LO:46.37);ALT=A[chr17:36912134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36909587	+	chr17	36912136	+	.	0	112	6386451_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6386451_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36897001_36922001_49C;SPAN=2549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:110 GQ:30 PL:[330.0, 30.0, 0.0] SR:112 DR:0 LR:-330.1 LO:330.1);ALT=T[chr17:36912136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36912245	+	chr17	36916683	+	.	3	28	6386464_1	79.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6386464_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36897001_36922001_176C;SPAN=4438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:85 GQ:79.4 PL:[79.4, 0.0, 125.6] SR:28 DR:3 LR:-79.3 LO:79.91);ALT=T[chr17:36916683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36916862	+	chr17	36918663	+	.	4	124	6386478_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6386478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36897001_36922001_10C;SPAN=1801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:145 GQ:25.9 PL:[402.6, 25.9, 0.0] SR:124 DR:4 LR:-407.4 LO:407.4);ALT=G[chr17:36918663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	36977327	+	chr17	36981419	+	.	0	10	6386927_1	6.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6386927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_36970501_36995501_309C;SPAN=4092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:98 GQ:6.5 PL:[6.5, 0.0, 230.9] SR:10 DR:0 LR:-6.459 LO:19.48);ALT=C[chr17:36981419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	37026511	+	chr17	37034337	+	.	0	17	6386834_1	33.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6386834_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_37019501_37044501_342C;SPAN=7826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:17 DR:0 LR:-33.63 LO:38.73);ALT=G[chr17:37034337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	37793518	+	chr17	37809730	+	.	27	0	6389676_1	74.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6389676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:37793518(+)-17:37809730(-)__17_37803501_37828501D;SPAN=16212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:53 GQ:51.8 PL:[74.9, 0.0, 51.8] SR:0 DR:27 LR:-74.95 LO:74.95);ALT=C[chr17:37809730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	38219346	+	chr17	38230443	+	.	9	6	6391375_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6391375_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_38195501_38220501_349C;SPAN=11097;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:15 GQ:5.9 PL:[29.0, 0.0, 5.9] SR:6 DR:9 LR:-29.65 LO:29.65);ALT=G[chr17:38230443[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	38474700	+	chr17	38487107	+	.	0	9	6391795_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6391795_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_38465001_38490001_1C;SPAN=12407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:9 DR:0 LR:-9.932 LO:18.32);ALT=G[chr17:38487107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	38785249	+	chr17	38786966	+	.	5	9	6393091_1	21.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTGT;MAPQ=2;MATEID=6393091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_38783501_38808501_141C;SPAN=1717;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:90 GQ:21.8 PL:[21.8, 0.0, 196.7] SR:9 DR:5 LR:-21.83 LO:30.03);ALT=T[chr17:38786966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	38798825	+	chr17	38804023	+	.	10	0	6393118_1	2.0	.	DISC_MAPQ=19;EVDNC=DSCRD;IMPRECISE;MAPQ=19;MATEID=6393118_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:38798825(+)-17:38804023(-)__17_38783501_38808501D;SPAN=5198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:113 GQ:2.6 PL:[2.6, 0.0, 269.9] SR:0 DR:10 LR:-2.396 LO:18.83);ALT=A[chr17:38804023[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	39240803	+	chr17	39296466	-	.	24	19	6394640_1	99.0	.	DISC_MAPQ=15;EVDNC=ASDIS;HOMSEQ=GCAGCAGCTGGGGTGGCAGCAGGTGGGCTGGCAGCACACAGACTGGCAGCACTGGGG;MAPQ=29;MATEID=6394640_2;MATENM=5;NM=2;NUMPARTS=2;SCTG=c_17_39273501_39298501_252C;SPAN=55663;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:19 DR:24 LR:-132.0 LO:132.0);ALT=C]chr17:39296466];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	39274434	+	chr17	39254137	+	.	11	0	6394643_1	24.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6394643_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:39254137(-)-17:39274434(+)__17_39273501_39298501D;SPAN=20297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:0 DR:11 LR:-24.12 LO:26.03);ALT=]chr17:39274434]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	39578956	+	chr17	39595309	+	.	12	0	6395379_1	30.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6395379_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:39578956(+)-17:39595309(-)__17_39567501_39592501D;SPAN=16353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:0 DR:12 LR:-30.67 LO:30.91);ALT=G[chr17:39595309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	39595512	+	chr17	39579067	+	.	18	0	6395381_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6395381_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:39579067(-)-17:39595512(+)__17_39567501_39592501D;SPAN=16445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:36 GQ:36.5 PL:[49.7, 0.0, 36.5] SR:0 DR:18 LR:-49.75 LO:49.75);ALT=]chr17:39595512]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	39845321	+	chr17	39846339	+	.	14	22	6396253_1	55.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6396253_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_39837001_39862001_57C;SPAN=1018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:196 GQ:55.9 PL:[55.9, 0.0, 419.0] SR:22 DR:14 LR:-55.83 LO:72.04);ALT=G[chr17:39846339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40118918	+	chr17	40120094	+	.	8	0	6396999_1	10.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6396999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40118918(+)-17:40120094(-)__17_40106501_40131501D;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:0 DR:8 LR:-10.42 LO:16.64);ALT=G[chr17:40120094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40134421	+	chr17	40135581	+	.	5	4	6397407_1	2.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=7;MATEID=6397407_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40131001_40156001_234C;SPAN=1160;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:4 DR:5 LR:-2.246 LO:13.27);ALT=T[chr17:40135581[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40149261	+	chr17	40169357	+	GGCTTTTGTATAATAATTATAAGCTTCATTGTAATCTTTCTTGGCATAGTATGCATTTCCTTGTTCCTTGAAAGTCTCTGCTTC	33	39	6397494_1	99.0	.	DISC_MAPQ=56;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GGCTTTTGTATAATAATTATAAGCTTCATTGTAATCTTTCTTGGCATAGTATGCATTTCCTTGTTCCTTGAAAGTCTCTGCTTC;MAPQ=60;MATEID=6397494_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_17_40155501_40180501_306C;SPAN=20096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:53 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:39 DR:33 LR:-155.1 LO:155.1);ALT=T[chr17:40169357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40152646	+	chr17	40169365	+	.	13	0	6397496_1	28.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6397496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40152646(+)-17:40169365(-)__17_40155501_40180501D;SPAN=16719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:55 GQ:28.1 PL:[28.1, 0.0, 104.0] SR:0 DR:13 LR:-28.01 LO:30.54);ALT=T[chr17:40169365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40172242	+	chr17	40174415	+	.	17	0	6397551_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6397551_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40172242(+)-17:40174415(-)__17_40155501_40180501D;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:79 GQ:34.7 PL:[34.7, 0.0, 156.8] SR:0 DR:17 LR:-34.71 LO:39.14);ALT=G[chr17:40174415[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40172252	+	chr17	40173579	+	.	10	0	6397552_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6397552_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40172252(+)-17:40173579(-)__17_40155501_40180501D;SPAN=1327;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:0 DR:10 LR:-14.86 LO:21.25);ALT=G[chr17:40173579[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40280820	+	chr17	40282355	+	.	0	14	6397812_1	19.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6397812_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40278001_40303001_157C;SPAN=1535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:101 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:14 DR:0 LR:-18.85 LO:29.27);ALT=T[chr17:40282355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40282608	+	chr17	40306911	+	.	115	8	6397962_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6397962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40302501_40327501_150C;SPAN=24303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:40 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:8 DR:115 LR:-340.0 LO:340.0);ALT=A[chr17:40306911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40289896	+	chr17	40306911	+	.	5	2	6397963_1	5.0	.	DISC_MAPQ=36;EVDNC=ASDIS;MAPQ=60;MATEID=6397963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40302501_40327501_65C;SPAN=17015;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:40 GQ:5.6 PL:[5.6, 0.0, 91.4] SR:2 DR:5 LR:-5.668 LO:10.21);ALT=T[chr17:40306911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40498732	+	chr17	40500406	+	.	0	10	6398555_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6398555_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40498501_40523501_202C;SPAN=1674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:101 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:10 DR:0 LR:-5.647 LO:19.35);ALT=C[chr17:40500406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40498779	+	chr17	40540371	+	.	8	0	6398666_1	14.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6398666_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40498779(+)-17:40540371(-)__17_40523001_40548001D;SPAN=41592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:46 GQ:14 PL:[14.0, 0.0, 96.5] SR:0 DR:8 LR:-13.95 LO:17.59);ALT=C[chr17:40540371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40500574	+	chr17	40540378	+	.	8	0	6398668_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6398668_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40500574(+)-17:40540378(-)__17_40523001_40548001D;SPAN=39804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.59 LO:17.19);ALT=G[chr17:40540378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40611025	+	chr17	40612877	+	.	12	0	6399185_1	15.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6399185_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40611025(+)-17:40612877(-)__17_40596501_40621501D;SPAN=1852;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:89 GQ:15.5 PL:[15.5, 0.0, 200.3] SR:0 DR:12 LR:-15.5 LO:24.93);ALT=G[chr17:40612877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40613029	+	chr17	40618447	+	.	0	7	6399190_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6399190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_40596501_40621501_219C;SPAN=5418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:85 GQ:0.2 PL:[0.2, 0.0, 204.8] SR:7 DR:0 LR:-0.07842 LO:12.95);ALT=C[chr17:40618447[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40925570	+	chr17	40926663	+	.	14	0	6400062_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6400062_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40925570(+)-17:40926663(-)__17_40915001_40940001D;SPAN=1093;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:100 GQ:19.1 PL:[19.1, 0.0, 223.7] SR:0 DR:14 LR:-19.12 LO:29.33);ALT=A[chr17:40926663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40925897	+	chr17	40927397	+	AAAGCTTCCTGTGGAGTCGATCCAGATTGTATTAGAGGAACTGAGGAAGAA	0	39	6400066_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AAAGCTTCCTGTGGAGTCGATCCAGATTGTATTAGAGGAACTGAGGAAGAA;MAPQ=60;MATEID=6400066_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_40915001_40940001_325C;SPAN=1500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:90 GQ:99 PL:[104.3, 0.0, 114.2] SR:39 DR:0 LR:-104.4 LO:104.4);ALT=G[chr17:40927397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	40972910	+	chr17	40976212	+	.	11	0	6400243_1	14.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6400243_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:40972910(+)-17:40976212(-)__17_40964001_40989001D;SPAN=3302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:79 GQ:14.9 PL:[14.9, 0.0, 176.6] SR:0 DR:11 LR:-14.91 LO:23.02);ALT=G[chr17:40976212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41113371	+	chr17	41116123	+	.	0	26	6400954_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6400954_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_41111001_41136001_260C;SPAN=2752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:97 GQ:59.6 PL:[59.6, 0.0, 175.1] SR:26 DR:0 LR:-59.55 LO:62.74);ALT=G[chr17:41116123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41113419	+	chr17	41116418	+	.	23	0	6400955_1	45.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6400955_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41113419(+)-17:41116418(-)__17_41111001_41136001D;SPAN=2999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:114 GQ:45.2 PL:[45.2, 0.0, 230.0] SR:0 DR:23 LR:-45.04 LO:52.22);ALT=C[chr17:41116418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41150578	+	chr17	41151947	+	.	51	0	6401112_1	99.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6401112_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41150578(+)-17:41151947(-)__17_41135501_41160501D;SPAN=1369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:121 GQ:99 PL:[135.8, 0.0, 155.6] SR:0 DR:51 LR:-135.6 LO:135.7);ALT=C[chr17:41151947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41150848	+	chr17	41151948	+	.	0	55	6401114_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6401114_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_41135501_41160501_99C;SPAN=1100;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:122 GQ:99 PL:[148.7, 0.0, 145.4] SR:55 DR:0 LR:-148.5 LO:148.5);ALT=G[chr17:41151948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41152107	+	chr17	41154889	+	.	18	0	6401117_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6401117_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41152107(+)-17:41154889(-)__17_41135501_41160501D;SPAN=2782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:18 DP:562 GQ:92.4 PL:[0.0, 92.4, 1548.0] SR:0 DR:18 LR:92.84 LO:25.77);ALT=T[chr17:41154889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41158948	+	chr17	41164956	+	.	9	0	6401147_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6401147_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41158948(+)-17:41164956(-)__17_41135501_41160501D;SPAN=6008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:0 DR:9 LR:-15.35 LO:19.68);ALT=A[chr17:41164956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41158986	+	chr17	41164196	+	.	27	23	6401148_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6401148_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_41135501_41160501_173C;SPAN=5210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:38 GQ:10.2 PL:[112.2, 10.2, 0.0] SR:23 DR:27 LR:-112.2 LO:112.2);ALT=G[chr17:41164196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41277742	+	chr17	41290671	+	.	8	0	6401480_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6401480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41277742(+)-17:41290671(-)__17_41258001_41283001D;SPAN=12929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:32 GQ:17.9 PL:[17.9, 0.0, 57.5] SR:0 DR:8 LR:-17.74 LO:19.02);ALT=T[chr17:41290671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41363992	+	chr17	41365037	+	.	9	0	6401976_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6401976_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:41363992(+)-17:41365037(-)__17_41356001_41381001D;SPAN=1045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.326 LO:17.45);ALT=G[chr17:41365037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	41852306	+	chr17	41856166	+	.	0	10	6403508_1	11.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=6403508_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_41846001_41871001_332C;SPAN=3860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:79 GQ:11.6 PL:[11.6, 0.0, 179.9] SR:10 DR:0 LR:-11.61 LO:20.48);ALT=C[chr17:41856166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42148553	+	chr17	42151527	+	.	0	8	6404520_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=6404520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42140001_42165001_126C;SPAN=2974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:8 DR:0 LR:-2.567 LO:15.16);ALT=T[chr17:42151527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42260463	+	chr17	42263933	+	.	7	4	6404878_1	12.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6404878_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42262501_42287501_14C;SPAN=3470;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:52 GQ:12.5 PL:[12.5, 0.0, 111.5] SR:4 DR:7 LR:-12.32 LO:17.12);ALT=T[chr17:42263933[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42294074	+	chr17	42295540	+	.	0	4	6404990_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6404990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42287001_42312001_172C;SPAN=1466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:78 GQ:7.8 PL:[0.0, 7.8, 204.6] SR:4 DR:0 LR:7.928 LO:6.554);ALT=T[chr17:42295540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42387480	-	chr17	42388876	+	.	3	2	6405543_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCA;MAPQ=60;MATEID=6405543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42385001_42410001_297C;SPAN=1396;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:68 GQ:5.1 PL:[0.0, 5.1, 174.9] SR:2 DR:3 LR:5.219 LO:6.798);ALT=[chr17:42388876[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	42400275	+	chr17	42402091	+	.	22	0	6405573_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6405573_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:42400275(+)-17:42402091(-)__17_42385001_42410001D;SPAN=1816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:66 GQ:54.8 PL:[54.8, 0.0, 104.3] SR:0 DR:22 LR:-54.74 LO:55.62);ALT=C[chr17:42402091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42400948	+	chr17	42402078	+	.	0	10	6405576_1	15.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=6405576_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42385001_42410001_339C;SPAN=1130;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:65 GQ:15.5 PL:[15.5, 0.0, 140.9] SR:10 DR:0 LR:-15.4 LO:21.4);ALT=G[chr17:42402078[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42422703	+	chr17	42426522	+	.	48	2	6405863_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GCAGG;MAPQ=60;MATEID=6405863_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_42409501_42434501_444C;SPAN=3819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:207 GQ:99 PL:[214.7, 0.0, 287.3] SR:2 DR:48 LR:-214.6 LO:215.2);ALT=G[chr17:42426522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	42422754	+	chr17	42426787	+	.	52	0	6405866_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6405866_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:42422754(+)-17:42426787(-)__17_42409501_42434501D;SPAN=4033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:98 GQ:92.3 PL:[145.1, 0.0, 92.3] SR:0 DR:52 LR:-145.7 LO:145.7);ALT=C[chr17:42426787[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	43112368	+	chr17	43138254	+	.	13	4	6408006_1	36.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6408006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_43120001_43145001_280C;SPAN=25886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:48 GQ:36.5 PL:[36.5, 0.0, 79.4] SR:4 DR:13 LR:-36.51 LO:37.4);ALT=C[chr17:43138254[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	43112371	+	chr17	43128726	+	.	8	0	6408007_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6408007_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:43112371(+)-17:43128726(-)__17_43120001_43145001D;SPAN=16355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:23 GQ:20.3 PL:[20.3, 0.0, 33.5] SR:0 DR:8 LR:-20.18 LO:20.41);ALT=C[chr17:43128726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45704565	+	chr17	45706499	+	.	7	18	6416488_1	41.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCTTGAGCCCAG;MAPQ=60;MATEID=6416488_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_45692501_45717501_232C;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:92 GQ:41.3 PL:[41.3, 0.0, 179.9] SR:18 DR:7 LR:-41.1 LO:46.15);ALT=G[chr17:45706499[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45752148	+	chr17	45753773	+	.	2	7	6416741_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6416741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_45741501_45766501_236C;SPAN=1625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:7 DR:2 LR:-0.9411 LO:14.92);ALT=G[chr17:45753773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45755779	+	chr17	45757386	+	.	5	4	6416750_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6416750_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_45741501_45766501_342C;SPAN=1607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:4 DR:5 LR:-0.9411 LO:14.92);ALT=C[chr17:45757386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45758049	+	chr17	45759768	+	.	14	0	6416759_1	23.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6416759_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:45758049(+)-17:45759768(-)__17_45741501_45766501D;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:85 GQ:23.3 PL:[23.3, 0.0, 181.7] SR:0 DR:14 LR:-23.19 LO:30.41);ALT=T[chr17:45759768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45904572	+	chr17	45905866	+	.	0	13	6417114_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6417114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_45888501_45913501_210C;SPAN=1294;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:80 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:13 DR:0 LR:-21.24 LO:28.16);ALT=T[chr17:45905866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	45906023	+	chr17	45908824	+	.	16	0	6417117_1	26.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6417117_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:45906023(+)-17:45908824(-)__17_45888501_45913501D;SPAN=2801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:96 GQ:26.9 PL:[26.9, 0.0, 205.1] SR:0 DR:16 LR:-26.81 LO:34.85);ALT=G[chr17:45908824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46019180	+	chr17	46020670	+	.	0	5	6417616_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6417616_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46011001_46036001_278C;SPAN=1490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:76 GQ:3.9 PL:[0.0, 3.9, 191.4] SR:5 DR:0 LR:4.085 LO:8.747);ALT=G[chr17:46020670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46125826	+	chr17	46127969	+	.	5	3	6417918_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=6417918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46109001_46134001_38C;SPAN=2143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:3 DR:5 LR:2.36 LO:12.64);ALT=T[chr17:46127969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46154425	+	chr17	46178702	+	.	10	0	6418406_1	24.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6418406_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46154425(+)-17:46178702(-)__17_46158001_46183001D;SPAN=24277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:33 GQ:24.2 PL:[24.2, 0.0, 53.9] SR:0 DR:10 LR:-24.07 LO:24.77);ALT=A[chr17:46178702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46654382	+	chr17	46667487	+	.	38	10	6419627_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;MAPQ=60;MATEID=6419627_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46648001_46673001_284C;SPAN=13105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:86 GQ:98.9 PL:[108.8, 0.0, 98.9] SR:10 DR:38 LR:-108.8 LO:108.8);ALT=A[chr17:46667487[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46667928	+	chr17	46679434	+	.	11	0	6419667_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6419667_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46667928(+)-17:46679434(-)__17_46648001_46673001D;SPAN=11506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:61 GQ:20 PL:[20.0, 0.0, 125.6] SR:0 DR:11 LR:-19.78 LO:24.38);ALT=G[chr17:46679434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46667951	+	chr17	46681288	+	.	0	17	6419668_1	42.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6419668_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46648001_46673001_104C;SPAN=13337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:49 GQ:42.8 PL:[42.8, 0.0, 75.8] SR:17 DR:0 LR:-42.84 LO:43.35);ALT=G[chr17:46681288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46667953	+	chr17	46677808	+	.	45	58	6419669_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6419669_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46648001_46673001_154C;SPAN=9855;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:46 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:58 DR:45 LR:-241.0 LO:241.0);ALT=T[chr17:46677808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46674034	+	chr17	46675096	+	.	7	7	6419700_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=6419700_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46672501_46697501_380C;SPAN=1062;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:101 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:7 DR:7 LR:-12.25 LO:24.22);ALT=C[chr17:46675096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46677910	+	chr17	46679435	+	.	0	49	6419708_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGTA;MAPQ=60;MATEID=6419708_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46672501_46697501_169C;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:98 GQ:99 PL:[135.2, 0.0, 102.2] SR:49 DR:0 LR:-135.4 LO:135.4);ALT=A[chr17:46679435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46681408	+	chr17	46683491	+	.	0	17	6419718_1	33.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6419718_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46672501_46697501_225C;SPAN=2083;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:85 GQ:33.2 PL:[33.2, 0.0, 171.8] SR:17 DR:0 LR:-33.09 LO:38.53);ALT=G[chr17:46683491[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46685460	+	chr17	46687880	+	.	8	3	6419724_1	8.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6419724_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46672501_46697501_325C;SPAN=2420;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:3 DR:8 LR:-8.035 LO:17.94);ALT=G[chr17:46687880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46904668	+	chr17	46907511	+	.	28	0	6420344_1	77.0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=6420344_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46904668(+)-17:46907511(-)__17_46893001_46918001D;SPAN=2843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:55 GQ:54.5 PL:[77.6, 0.0, 54.5] SR:0 DR:28 LR:-77.71 LO:77.71);ALT=T[chr17:46907511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46908490	+	chr17	46925425	+	.	31	0	6420392_1	88.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6420392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46908490(+)-17:46925425(-)__17_46917501_46942501D;SPAN=16935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:50 GQ:32.6 PL:[88.7, 0.0, 32.6] SR:0 DR:31 LR:-90.21 LO:90.21);ALT=T[chr17:46925425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46908493	+	chr17	46919058	+	.	54	0	6420394_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6420394_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46908493(+)-17:46919058(-)__17_46917501_46942501D;SPAN=10565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:51 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=A[chr17:46919058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46919251	+	chr17	46925426	+	.	0	59	6420400_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6420400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46917501_46942501_241C;SPAN=6175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:102 GQ:78.2 PL:[167.3, 0.0, 78.2] SR:59 DR:0 LR:-168.8 LO:168.8);ALT=T[chr17:46925426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46919308	+	chr17	46925681	+	.	8	0	6420401_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6420401_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46919308(+)-17:46925681(-)__17_46917501_46942501D;SPAN=6373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=A[chr17:46925681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46926740	+	chr17	46928921	+	AGGAGCTAGAAACCCTACAGAGCATCAATAAGAAGTTGGAACTGAAAGTGAAAGAACAGAAGGACTATTGGGAGACAGAGCTGCTTCA	4	24	6420431_1	64.0	.	DISC_MAPQ=47;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=AGGAGCTAGAAACCCTACAGAGCATCAATAAGAAGTTGGAACTGAAAGTGAAAGAACAGAAGGACTATTGGGAGACAGAGCTGCTTCA;MAPQ=60;MATEID=6420431_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_46917501_46942501_177C;SPAN=2181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:79 GQ:64.4 PL:[64.4, 0.0, 127.1] SR:24 DR:4 LR:-64.42 LO:65.56);ALT=G[chr17:46928921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46929990	+	chr17	46933453	+	AGGAAGGACCAGAAGAAGCTCGAGCAGACAGTGGAGCAAATGAAGCAGAATGAAACTACTGCAATGAAGAAACAACAGGAATTAAT	7	16	6420446_1	41.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AGGAAGGACCAGAAGAAGCTCGAGCAGACAGTGGAGCAAATGAAGCAGAATGAAACTACTGCAATGAAGAAACAACAGGAATTAAT;MAPQ=60;MATEID=6420446_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_46917501_46942501_171C;SPAN=3463;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:81 GQ:41 PL:[41.0, 0.0, 153.2] SR:16 DR:7 LR:-40.77 LO:44.56);ALT=G[chr17:46933453[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46937814	+	chr17	46940199	+	TCCAAGAAAGTTCTTCCCCCAGCCC	6	13	6420478_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCCAAGAAAGTTCTTCCCCCAGCCC;MAPQ=60;MATEID=6420478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46917501_46942501_167C;SPAN=2385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:13 DR:6 LR:-26.49 LO:33.08);ALT=A[chr17:46940199[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	46970244	+	chr17	46972515	+	.	11	0	6420832_1	5.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=6420832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:46970244(+)-17:46972515(-)__17_46966501_46991501D;SPAN=2271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:113 GQ:5.9 PL:[5.9, 0.0, 266.6] SR:0 DR:11 LR:-5.697 LO:21.19);ALT=G[chr17:46972515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47007975	+	chr17	47009004	+	.	0	42	6420675_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6420675_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_46991001_47016001_79C;SPAN=1029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:103 GQ:99 PL:[110.9, 0.0, 137.3] SR:42 DR:0 LR:-110.7 LO:110.9);ALT=C[chr17:47009004[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47009081	+	chr17	47010567	+	.	0	8	6420679_1	0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6420679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_46991001_47016001_339C;SPAN=1486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:101 GQ:0.6 PL:[0.0, 0.6, 244.2] SR:8 DR:0 LR:0.9554 LO:14.66);ALT=T[chr17:47010567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47018439	+	chr17	47022102	+	.	12	0	6420924_1	11.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6420924_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:47018439(+)-17:47022102(-)__17_47015501_47040501D;SPAN=3663;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:104 GQ:11.6 PL:[11.6, 0.0, 239.3] SR:0 DR:12 LR:-11.44 LO:24.06);ALT=G[chr17:47022102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47700241	+	chr17	47755294	+	.	9	7	6423372_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6423372_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_47750501_47775501_70C;SPAN=55053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:50 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:7 DR:9 LR:-32.67 LO:34.1);ALT=G[chr17:47755294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	47778873	+	chr17	47780218	+	.	0	10	6423204_1	10.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=6423204_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_47775001_47800001_318C;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:10 DR:0 LR:-10.52 LO:20.25);ALT=C[chr17:47780218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48445659	+	chr17	48447814	+	ATGGGCACCTGGGTGCCAGCGGAAATGGCGCTGTGTTGCAATGATGTTCCCAGCATGAACATAGTG	0	26	6425240_1	60.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=ATGGGCACCTGGGTGCCAGCGGAAATGGCGCTGTGTTGCAATGATGTTCCCAGCATGAACATAGTG;MAPQ=60;MATEID=6425240_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_48436501_48461501_220C;SPAN=2155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:94 GQ:60.5 PL:[60.5, 0.0, 166.1] SR:26 DR:0 LR:-60.36 LO:63.17);ALT=C[chr17:48447814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48445705	+	chr17	48450490	+	.	13	0	6425242_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6425242_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:48445705(+)-17:48450490(-)__17_48436501_48461501D;SPAN=4785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:94 GQ:17.6 PL:[17.6, 0.0, 209.0] SR:0 DR:13 LR:-17.45 LO:27.16);ALT=G[chr17:48450490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48447976	+	chr17	48450490	+	.	25	0	6425246_1	58.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6425246_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:48447976(+)-17:48450490(-)__17_48436501_48461501D;SPAN=2514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:90 GQ:58.1 PL:[58.1, 0.0, 160.4] SR:0 DR:25 LR:-58.14 LO:60.79);ALT=A[chr17:48450490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48797123	+	chr17	48814320	+	.	20	0	6426625_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6426625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:48797123(+)-17:48814320(-)__17_48779501_48804501D;SPAN=17197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:69 GQ:47.3 PL:[47.3, 0.0, 119.9] SR:0 DR:20 LR:-47.33 LO:49.08);ALT=G[chr17:48814320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48818608	+	chr17	48821065	+	CCGCTGGCCCAACAGGCAAAAATGAAGAAAAAATTCAGGTTCTAACAGACAAAATTGATGTACTTCTGCAAC	0	21	6426536_1	48.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCGCTGGCCCAACAGGCAAAAATGAAGAAAAAATTCAGGTTCTAACAGACAAAATTGATGTACTTCTGCAAC;MAPQ=60;MATEID=6426536_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_48804001_48829001_57C;SPAN=2457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:76 GQ:48.8 PL:[48.8, 0.0, 134.6] SR:21 DR:0 LR:-48.73 LO:51.01);ALT=G[chr17:48821065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48819092	+	chr17	48821065	+	.	4	14	6426539_1	31.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6426539_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_17_48804001_48829001_57C;SPAN=1973;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:78 GQ:31.7 PL:[31.7, 0.0, 157.1] SR:14 DR:4 LR:-31.68 LO:36.46);ALT=G[chr17:48821065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	48824063	+	chr17	48827860	+	.	14	4	6426549_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6426549_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_17_48804001_48829001_287C;SPAN=3797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:92 GQ:28.1 PL:[28.1, 0.0, 193.1] SR:4 DR:14 LR:-27.89 LO:35.18);ALT=G[chr17:48827860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49231056	+	chr17	49233010	+	.	63	0	6428431_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6428431_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49231056(+)-17:49233010(-)__17_49220501_49245501D;SPAN=1954;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:92 GQ:38 PL:[183.2, 0.0, 38.0] SR:0 DR:63 LR:-188.2 LO:188.2);ALT=G[chr17:49233010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49231060	+	chr17	49238519	+	.	11	0	6428432_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6428432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49231060(+)-17:49238519(-)__17_49220501_49245501D;SPAN=7459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:105 GQ:8 PL:[8.0, 0.0, 245.6] SR:0 DR:11 LR:-7.864 LO:21.56);ALT=G[chr17:49238519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49231067	+	chr17	49237338	+	.	60	0	6428433_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6428433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49231067(+)-17:49237338(-)__17_49220501_49245501D;SPAN=6271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:109 GQ:95.9 PL:[168.5, 0.0, 95.9] SR:0 DR:60 LR:-169.6 LO:169.6);ALT=A[chr17:49237338[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49233142	+	chr17	49237341	+	.	2	77	6428443_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6428443_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_17_49220501_49245501_47C;SPAN=4199;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:132 GQ:96.5 PL:[221.9, 0.0, 96.5] SR:77 DR:2 LR:-224.3 LO:224.3);ALT=G[chr17:49237341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49233142	+	chr17	49239086	+	CTTCCGAAGATCTTCTCAAGGAACACTACGTTGACCTGAAGGACCGTCCATTCTTTGCCGGCCTGGTGAAATACATGCACTCAGGGCCGGTAGTTGCCATGGTCTGGGAGGGGCTGAATGTGGTGAAGACGGGCCGAGTCATGCTCGGGGAGACCAACCCTGCAGACTCCAAGCCTGGGACCATCCGTGGAGACTTCTGCATACAAGTTGG	0	100	6428444_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CTTCCGAAGATCTTCTCAAGGAACACTACGTTGACCTGAAGGACCGTCCATTCTTTGCCGGCCTGGTGAAATACATGCACTCAGGGCCGGTAGTTGCCATGGTCTGGGAGGGGCTGAATGTGGTGAAGACGGGCCGAGTCATGCTCGGGGAGACCAACCCTGCAGACTCCAAGCCTGGGACCATCCGTGGAGACTTCTGCATACAAGTTGG;MAPQ=60;MATEID=6428444_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_49220501_49245501_47C;SPAN=5944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:124 GQ:2.9 PL:[296.6, 0.0, 2.9] SR:100 DR:0 LR:-313.9 LO:313.9);ALT=G[chr17:49239086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49237444	+	chr17	49238520	+	.	0	44	6428458_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=6428458_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_49220501_49245501_47C;SPAN=1076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:111 GQ:99 PL:[115.4, 0.0, 151.7] SR:44 DR:0 LR:-115.2 LO:115.5);ALT=T[chr17:49238520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49244001	+	chr17	49245599	+	.	30	0	6428485_1	89.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6428485_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49244001(+)-17:49245599(-)__17_49220501_49245501D;SPAN=1598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=T[chr17:49245599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49244290	+	chr17	49245600	+	.	16	0	6428487_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6428487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49244290(+)-17:49245600(-)__17_49220501_49245501D;SPAN=1310;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:16 DP:251 GQ:14.8 PL:[0.0, 14.8, 637.0] SR:0 DR:16 LR:15.19 LO:27.77);ALT=C[chr17:49245600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49244307	+	chr17	49247296	+	.	10	0	6428488_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6428488_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:49244307(+)-17:49247296(-)__17_49220501_49245501D;SPAN=2989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:205 GQ:22.3 PL:[0.0, 22.3, 541.3] SR:0 DR:10 LR:22.53 LO:16.16);ALT=A[chr17:49247296[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	49338289	+	chr17	49340634	+	.	3	3	6428028_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6428028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_49318501_49343501_243C;SPAN=2345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:82 GQ:2.1 PL:[0.0, 2.1, 201.3] SR:3 DR:3 LR:2.41 LO:10.78);ALT=T[chr17:49340634[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	54949916	+	chr17	54952294	+	.	9	0	6442083_1	9.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6442083_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:54949916(+)-17:54952294(-)__17_54929001_54954001D;SPAN=2378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:0 DR:9 LR:-9.661 LO:18.26);ALT=A[chr17:54952294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55055597	+	chr17	55058439	+	.	22	0	6441931_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6441931_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55055597(+)-17:55058439(-)__17_55051501_55076501D;SPAN=2842;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:98 GQ:46.1 PL:[46.1, 0.0, 191.3] SR:0 DR:22 LR:-46.07 LO:51.12);ALT=G[chr17:55058439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55058592	+	chr17	55062737	+	.	0	11	6441942_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6441942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_55051501_55076501_137C;SPAN=4145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:97 GQ:10.1 PL:[10.1, 0.0, 224.6] SR:11 DR:0 LR:-10.03 LO:21.97);ALT=G[chr17:55062737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55089757	+	chr17	55092846	+	.	54	0	6442414_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6442414_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55089757(+)-17:55092846(-)__17_55076001_55101001D;SPAN=3089;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:5 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=T[chr17:55092846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55255418	+	chr22	22249852	-	.	9	0	6442616_1	20.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6442616_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55255418(+)-22:22249852(+)__17_55247501_55272501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=G]chr22:22249852];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr17	55338128	-	chr17	55340296	+	.	2	2	6442946_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6442946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_55321001_55346001_259C;SPAN=2168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:86 GQ:9.9 PL:[0.0, 9.9, 227.7] SR:2 DR:2 LR:10.1 LO:6.381);ALT=[chr17:55340296[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	55687811	+	chr17	55689915	+	.	70	45	6444031_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6444031_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_55688501_55713501_320C;SPAN=2104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:33 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:45 DR:70 LR:-254.2 LO:254.2);ALT=T[chr17:55689915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55918414	+	chr17	55926600	+	GTTGACAGGTAGACTTGAAGTTTGGATTGAATAGATCAAAAGCTCTTTGACCAGACCCATACACTGAATAAAACTT	0	37	6444708_1	97.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTGACAGGTAGACTTGAAGTTTGGATTGAATAGATCAAAAGCTCTTTGACCAGACCCATACACTGAATAAAACTT;MAPQ=60;MATEID=6444708_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_55909001_55934001_1C;SPAN=8186;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:90 GQ:97.7 PL:[97.7, 0.0, 120.8] SR:37 DR:0 LR:-97.75 LO:97.89);ALT=C[chr17:55926600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55918621	+	chr17	55926600	+	.	7	24	6444710_1	74.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6444710_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTCT;SCTG=c_17_55909001_55934001_1C;SPAN=7979;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:93 GQ:74 PL:[74.0, 0.0, 149.9] SR:24 DR:7 LR:-73.83 LO:75.32);ALT=C[chr17:55926600[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	55918669	+	chr17	55927326	+	.	20	0	6444711_1	47.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6444711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:55918669(+)-17:55927326(-)__17_55909001_55934001D;SPAN=8657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:69 GQ:47.3 PL:[47.3, 0.0, 119.9] SR:0 DR:20 LR:-47.33 LO:49.08);ALT=G[chr17:55927326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	56353065	+	chr17	56355187	+	.	6	3	6445962_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=6445962_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_17_56350001_56375001_171C;SPAN=2122;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:104 GQ:8.1 PL:[0.0, 8.1, 267.3] SR:3 DR:6 LR:8.37 LO:10.14);ALT=T[chr17:56355187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	56770149	+	chr17	56772290	+	.	11	1	6447324_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6447324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_56766501_56791501_247C;SPAN=2141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:81 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:1 DR:11 LR:-14.37 LO:22.89);ALT=G[chr17:56772290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57177238	-	chr17	57178271	+	.	9	0	6448476_1	6.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6448476_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:57177238(-)-17:57178271(-)__17_57158501_57183501D;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:87 GQ:6.2 PL:[6.2, 0.0, 204.2] SR:0 DR:9 LR:-6.139 LO:17.59);ALT=[chr17:57178271[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	57189745	+	chr17	57232484	+	.	8	0	6448658_1	14.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6448658_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:57189745(+)-17:57232484(-)__17_57207501_57232501D;SPAN=42739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=T[chr17:57232484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57196909	+	chr17	57232485	+	.	8	0	6448659_1	14.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6448659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:57196909(+)-17:57232485(-)__17_57207501_57232501D;SPAN=35576;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=T[chr17:57232485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57409186	+	chr17	57430575	+	.	23	7	6449150_1	59.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6449150_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_57428001_57453001_321C;SPAN=21389;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:59 GQ:59.9 PL:[59.9, 0.0, 83.0] SR:7 DR:23 LR:-59.94 LO:60.15);ALT=G[chr17:57430575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57697534	+	chr17	57721635	+	.	0	9	6450212_1	8.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6450212_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_57697501_57722501_224C;SPAN=24101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:9 DR:0 LR:-7.764 LO:17.89);ALT=G[chr17:57721635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57785109	+	chr17	57808781	+	.	13	7	6450663_1	44.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6450663_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_17_57771001_57796001_40C;SPAN=23672;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:44 GQ:44.3 PL:[44.3, 0.0, 60.8] SR:7 DR:13 LR:-44.2 LO:44.37);ALT=G[chr17:57808781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57785109	+	chr17	57812696	+	CTCCTCAAGAGTTACTGATCTATGAAATGGCAGAGAATGGAAAAAATTGTGACCAGAGACGTGTAGCAATGAACAAGGAACATCATAATGGAAATTTCA	24	26	6450664_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=CTCCTCAAGAGTTACTGATCTATGAAATGGCAGAGAATGGAAAAAATTGTGACCAGAGACGTGTAGCAATGAACAAGGAACATCATAATGGAAATTTCA;MAPQ=60;MATEID=6450664_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_57771001_57796001_40C;SPAN=27587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:44 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:26 DR:24 LR:-128.7 LO:128.7);ALT=G[chr17:57812696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57808883	+	chr17	57812696	+	.	0	18	6450697_1	52.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=6450697_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCCC;SCTG=c_17_57771001_57796001_40C;SPAN=3813;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:18 DP:0 GQ:4.8 PL:[52.8, 4.8, 0.0] SR:18 DR:0 LR:-52.81 LO:52.81);ALT=G[chr17:57812696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	57814303	+	chr17	57815391	-	.	10	0	6450605_1	5.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6450605_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:57814303(+)-17:57815391(+)__17_57795501_57820501D;SPAN=1088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=G]chr17:57815391];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr17	57915759	+	chr17	57917125	+	.	7	6	6451084_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACAGG;MAPQ=60;MATEID=6451084_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_57893501_57918501_154C;SPAN=1366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:158 GQ:3.1 PL:[0.0, 3.1, 389.4] SR:6 DR:7 LR:3.194 LO:21.77);ALT=G[chr17:57917125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	58040672	+	chr17	58042008	+	.	27	0	6451584_1	64.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6451584_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:58040672(+)-17:58042008(-)__17_58040501_58065501D;SPAN=1336;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:90 GQ:64.7 PL:[64.7, 0.0, 153.8] SR:0 DR:27 LR:-64.74 LO:66.74);ALT=A[chr17:58042008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	58180028	+	chrX	15872810	+	.	20	0	7370825_1	59.0	.	DISC_MAPQ=37;EVDNC=DSCRD;IMPRECISE;MAPQ=37;MATEID=7370825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:58180028(+)-23:15872810(-)__23_15851501_15876501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:19 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:20 LR:-59.41 LO:59.41);ALT=G[chrX:15872810[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr17	59118770	+	chr17	59128793	+	TGTAATATATATATATATATATATAT	6	6	6454888_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTAATATATATATATATATATATAT;MAPQ=60;MATEID=6454888_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_59118501_59143501_74C;SPAN=10023;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:6 DR:6 LR:-17.03 LO:21.86);ALT=G[chr17:59128793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	65214940	+	chr17	65235548	+	.	0	9	6473554_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6473554_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_65219001_65244001_9C;SPAN=20608;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:9 DR:0 LR:-17.25 LO:20.3);ALT=T[chr17:65235548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	65214960	+	chr17	65241262	+	.	15	0	6473555_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6473555_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:65214960(+)-17:65241262(-)__17_65219001_65244001D;SPAN=26302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:37 GQ:39.5 PL:[39.5, 0.0, 49.4] SR:0 DR:15 LR:-39.49 LO:39.56);ALT=A[chr17:65241262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	65346452	+	chr17	65353418	+	.	0	7	6474125_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6474125_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_65341501_65366501_324C;SPAN=6966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:7 DR:0 LR:0.4634 LO:12.88);ALT=C[chr17:65353418[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	65562065	+	chr17	65561042	+	.	13	0	6474833_1	29.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=6474833_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:65561042(-)-17:65562065(+)__17_65562001_65587001D;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:52 GQ:29 PL:[29.0, 0.0, 95.0] SR:0 DR:13 LR:-28.83 LO:30.91);ALT=]chr17:65562065]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	66031956	+	chr17	66033224	+	.	17	5	6476553_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6476553_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_66027501_66052501_359C;SPAN=1268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:98 GQ:32.9 PL:[32.9, 0.0, 204.5] SR:5 DR:17 LR:-32.87 LO:40.05);ALT=G[chr17:66033224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66088392	-	chr17	66089409	+	.	10	0	6476700_1	8.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=6476700_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:66088392(-)-17:66089409(-)__17_66076501_66101501D;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:90 GQ:8.6 PL:[8.6, 0.0, 209.9] SR:0 DR:10 LR:-8.627 LO:19.88);ALT=[chr17:66089409[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	66244317	+	chr17	66246326	+	.	9	0	6477276_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6477276_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:66244317(+)-17:66246326(-)__17_66223501_66248501D;SPAN=2009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:103 GQ:2 PL:[2.0, 0.0, 246.2] SR:0 DR:9 LR:-1.804 LO:16.9);ALT=A[chr17:66246326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66508689	+	chr17	66511532	+	.	56	12	6478114_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6478114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_66493001_66518001_366C;SPAN=2843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:106 GQ:86.9 PL:[169.4, 0.0, 86.9] SR:12 DR:56 LR:-170.7 LO:170.7);ALT=G[chr17:66511532[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66511718	+	chr17	66518895	+	.	3	7	6478248_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6478248_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_66517501_66542501_243C;SPAN=7177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:7 DR:3 LR:-14.27 LO:19.37);ALT=G[chr17:66518895[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	66519098	+	chr17	66520153	+	.	8	0	6478258_1	6.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6478258_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:66519098(+)-17:66520153(-)__17_66517501_66542501D;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=G[chr17:66520153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72462909	+	chr17	72469670	+	.	35	0	6494684_1	92.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6494684_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:72462909(+)-17:72469670(-)__17_72446501_72471501D;SPAN=6761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:87 GQ:92 PL:[92.0, 0.0, 118.4] SR:0 DR:35 LR:-91.97 LO:92.16);ALT=C[chr17:72469670[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72470825	+	chr17	72473575	+	.	0	7	6494775_1	8.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6494775_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_72471001_72496001_71C;SPAN=2750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:56 GQ:8 PL:[8.0, 0.0, 126.8] SR:7 DR:0 LR:-7.935 LO:14.3);ALT=G[chr17:72473575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72733490	+	chr17	72739264	+	.	15	0	6495585_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6495585_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:72733490(+)-17:72739264(-)__17_72716001_72741001D;SPAN=5774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:78 GQ:28.4 PL:[28.4, 0.0, 160.4] SR:0 DR:15 LR:-28.38 LO:33.71);ALT=G[chr17:72739264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72733507	+	chr17	72736905	+	.	25	16	6495587_1	87.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=6495587_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_72716001_72741001_257C;SPAN=3398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:79 GQ:87.5 PL:[87.5, 0.0, 104.0] SR:16 DR:25 LR:-87.53 LO:87.61);ALT=G[chr17:72736905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	72769864	+	chr17	72772404	+	.	9	0	6495633_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6495633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:72769864(+)-17:72772404(-)__17_72765001_72790001D;SPAN=2540;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:89 GQ:5.6 PL:[5.6, 0.0, 210.2] SR:0 DR:9 LR:-5.597 LO:17.5);ALT=A[chr17:72772404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73008967	+	chr17	73015793	+	AATGGTGCAAAGCAAGCCGACAGTGACATCCCTCT	0	18	6496626_1	48.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AATGGTGCAAAGCAAGCCGACAGTGACATCCCTCT;MAPQ=60;MATEID=6496626_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_72985501_73010501_180C;SPAN=6826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:41 GQ:48.5 PL:[48.5, 0.0, 48.5] SR:18 DR:0 LR:-48.31 LO:48.32);ALT=G[chr17:73015793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73038393	+	chr17	73043018	+	.	43	0	6496664_1	99.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6496664_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73038393(+)-17:73043018(-)__17_73034501_73059501D;SPAN=4625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:105 GQ:99 PL:[113.6, 0.0, 140.0] SR:0 DR:43 LR:-113.5 LO:113.7);ALT=A[chr17:73043018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73144767	+	chr17	73150437	+	.	0	58	6496871_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6496871_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73132501_73157501_144C;SPAN=5670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:110 GQ:99 PL:[161.6, 0.0, 105.5] SR:58 DR:0 LR:-162.3 LO:162.3);ALT=C[chr17:73150437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73177284	+	chr17	73178476	+	.	0	9	6497029_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=59;MATEID=6497029_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73157001_73182001_102C;SPAN=1192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:78 GQ:8.6 PL:[8.6, 0.0, 180.2] SR:9 DR:0 LR:-8.577 LO:18.05);ALT=C[chr17:73178476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	114953559	+	chr17	73178992	+	.	40	0	7503369_1	99.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=7503369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73178992(-)-23:114953559(+)__23_114929501_114954501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:0 DR:40 LR:-125.4 LO:125.4);ALT=]chrX:114953559]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	73204715	+	chr17	73205916	+	.	0	5	6497820_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6497820_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73181501_73206501_487C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:66 GQ:1.2 PL:[0.0, 1.2, 161.7] SR:5 DR:0 LR:1.376 LO:9.064);ALT=G[chr17:73205916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73264275	+	chr17	73267222	+	TTGAGTGCTGTCTTCAGCAGCTGCTGGGTCTCTGCATCAAAGGACTGGATTTTATACTCCTCTCTACTGGGCTCCCCCATGACTAGCCAGCCCCGGTAGCTCTTGACTGGGCTGGGAATAAGGACAG	16	22	6497215_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CACCTG;INSERTION=TTGAGTGCTGTCTTCAGCAGCTGCTGGGTCTCTGCATCAAAGGACTGGATTTTATACTCCTCTCTACTGGGCTCCCCCATGACTAGCCAGCCCCGGTAGCTCTTGACTGGGCTGGGAATAAGGACAG;MAPQ=60;MATEID=6497215_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_73255001_73280001_154C;SPAN=2947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:60 GQ:56.3 PL:[89.3, 0.0, 56.3] SR:22 DR:16 LR:-89.78 LO:89.78);ALT=T[chr17:73267222[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73264323	+	chr17	73266288	+	.	17	0	6497216_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6497216_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73264323(+)-17:73266288(-)__17_73255001_73280001D;SPAN=1965;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:70 GQ:37.1 PL:[37.1, 0.0, 132.8] SR:0 DR:17 LR:-37.15 LO:40.17);ALT=T[chr17:73266288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73282922	+	chr17	73285434	+	.	8	0	6497403_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6497403_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73282922(+)-17:73285434(-)__17_73279501_73304501D;SPAN=2512;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:80 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:0 DR:8 LR:-4.734 LO:15.51);ALT=T[chr17:73285434[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73316637	+	chr17	73317740	+	.	3	3	6497676_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6497676_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73304001_73329001_178C;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:72 GQ:0.5 PL:[0.5, 0.0, 172.1] SR:3 DR:3 LR:-0.2994 LO:11.14);ALT=G[chr17:73317740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73328880	+	chr17	73389630	+	.	2	7	6497944_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6497944_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73377501_73402501_11C;SPAN=60750;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:7 DR:2 LR:-16.16 LO:19.94);ALT=T[chr17:73389630[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73389847	+	chr17	73401569	+	.	74	43	6497987_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6497987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73377501_73402501_60C;SPAN=11722;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:138 GQ:74.9 PL:[259.7, 0.0, 74.9] SR:43 DR:74 LR:-265.3 LO:265.3);ALT=C[chr17:73401569[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73663558	+	chr17	73664595	+	.	10	5	6498847_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6498847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73647001_73672001_294C;SPAN=1037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:94 GQ:11 PL:[11.0, 0.0, 215.6] SR:5 DR:10 LR:-10.84 LO:22.13);ALT=G[chr17:73664595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73663589	+	chr17	73667891	+	.	8	0	6498848_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6498848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73663589(+)-17:73667891(-)__17_73647001_73672001D;SPAN=4302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-2.025 LO:15.08);ALT=A[chr17:73667891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73845821	+	chr17	73847647	+	.	0	23	6499581_1	54.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=6499581_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73843001_73868001_274C;SPAN=1826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:81 GQ:54.2 PL:[54.2, 0.0, 140.0] SR:23 DR:0 LR:-53.98 LO:56.19);ALT=C[chr17:73847647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73845874	+	chr17	73851320	+	.	17	0	6499582_1	37.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6499582_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73845874(+)-17:73851320(-)__17_73843001_73868001D;SPAN=5446;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:69 GQ:37.4 PL:[37.4, 0.0, 129.8] SR:0 DR:17 LR:-37.42 LO:40.29);ALT=A[chr17:73851320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73847759	+	chr17	73851320	+	.	19	8	6499590_1	47.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6499590_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73843001_73868001_131C;SPAN=3561;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:83 GQ:47 PL:[47.0, 0.0, 152.6] SR:8 DR:19 LR:-46.83 LO:50.06);ALT=T[chr17:73851320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73898238	+	chr17	73900621	+	.	0	16	6499677_1	29.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6499677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73892001_73917001_304C;SPAN=2383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:85 GQ:29.9 PL:[29.9, 0.0, 175.1] SR:16 DR:0 LR:-29.79 LO:35.79);ALT=G[chr17:73900621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73898283	+	chr17	73900903	+	.	11	0	6499678_1	13.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6499678_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:73898283(+)-17:73900903(-)__17_73892001_73917001D;SPAN=2620;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:0 DR:11 LR:-13.55 LO:22.7);ALT=G[chr17:73900903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	73975593	+	chr17	73982264	+	.	0	15	6500164_1	27.0	.	EVDNC=ASSMB;HOMSEQ=ACAGG;MAPQ=60;MATEID=6500164_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_73965501_73990501_141C;SPAN=6671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:82 GQ:27.5 PL:[27.5, 0.0, 169.4] SR:15 DR:0 LR:-27.3 LO:33.34);ALT=G[chr17:73982264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	74063457	+	chr17	74068388	+	.	9	0	6500642_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6500642_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:74063457(+)-17:74068388(-)__17_74063501_74088501D;SPAN=4931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:0 DR:9 LR:-14.27 LO:19.37);ALT=T[chr17:74068388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	74097945	+	chr17	74099439	+	.	0	7	6500439_1	0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=6500439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_74088001_74113001_366C;SPAN=1494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:7 DR:0 LR:2.902 LO:12.57);ALT=C[chr17:74099439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	74097993	+	chr17	74099742	+	.	10	0	6500440_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6500440_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:74097993(+)-17:74099742(-)__17_74088001_74113001D;SPAN=1749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:0 DR:10 LR:-9.169 LO:19.98);ALT=C[chr17:74099742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	74723004	+	chr17	74729057	+	.	15	0	6502742_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6502742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:74723004(+)-17:74729057(-)__17_74725001_74750001D;SPAN=6053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:38 GQ:39.2 PL:[39.2, 0.0, 52.4] SR:0 DR:15 LR:-39.22 LO:39.33);ALT=C[chr17:74729057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	74725876	+	chr17	74729058	+	.	2	9	6502745_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6502745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_74725001_74750001_297C;SPAN=3182;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:75 GQ:16.1 PL:[16.1, 0.0, 164.6] SR:9 DR:2 LR:-15.99 LO:23.29);ALT=G[chr17:74729058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	75137188	+	chr17	75139645	+	.	8	0	6504094_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6504094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:75137188(+)-17:75139645(-)__17_75117001_75142001D;SPAN=2457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=A[chr17:75139645[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	75137189	+	chr17	75138726	+	.	19	7	6504095_1	41.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6504095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_75117001_75142001_177C;SPAN=1537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:77 GQ:41.9 PL:[41.9, 0.0, 144.2] SR:7 DR:19 LR:-41.86 LO:45.05);ALT=G[chr17:75138726[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	75447658	+	chr17	75478224	+	.	10	0	6505308_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6505308_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:75447658(+)-17:75478224(-)__17_75460001_75485001D;SPAN=30566;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=G[chr17:75478224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	75447661	+	chr17	75483504	+	.	11	0	6505309_1	25.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6505309_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:75447661(+)-17:75483504(-)__17_75460001_75485001D;SPAN=35843;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:0 DR:11 LR:-25.75 LO:26.84);ALT=C[chr17:75483504[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	75478418	+	chr17	75483505	+	.	13	25	6505354_1	85.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6505354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_75460001_75485001_411C;SPAN=5087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:88 GQ:85.1 PL:[85.1, 0.0, 128.0] SR:25 DR:13 LR:-85.09 LO:85.58);ALT=G[chr17:75483505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76122990	+	chr17	76124693	+	.	10	2	6507112_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6507112_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76121501_76146501_58C;SPAN=1703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:58 GQ:20.6 PL:[20.6, 0.0, 119.6] SR:2 DR:10 LR:-20.6 LO:24.64);ALT=G[chr17:76124693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76164798	+	chr17	76166897	+	.	87	22	6507342_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6507342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76146001_76171001_95C;SPAN=2099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:81 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:22 DR:87 LR:-277.3 LO:277.3);ALT=T[chr17:76166897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76181284	+	chr17	76183068	+	.	19	0	6507381_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6507381_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76181284(+)-17:76183068(-)__17_76170501_76195501D;SPAN=1784;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:74 GQ:42.8 PL:[42.8, 0.0, 135.2] SR:0 DR:19 LR:-42.67 LO:45.43);ALT=G[chr17:76183068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76183544	+	chr17	76198576	+	.	13	0	6507650_1	34.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6507650_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76183544(+)-17:76198576(-)__17_76195001_76220001D;SPAN=15032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:32 GQ:34.4 PL:[34.4, 0.0, 41.0] SR:0 DR:13 LR:-34.24 LO:34.3);ALT=G[chr17:76198576[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76187141	+	chr17	76198588	+	CCACCACG	0	7	6507403_1	12.0	.	EVDNC=ASSMB;INSERTION=CCACCACG;MAPQ=60;MATEID=6507403_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76170501_76195501_361C;SPAN=11447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:7 DR:0 LR:-12.54 LO:15.5);ALT=G[chr17:76198588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76374891	+	chr17	76388555	+	.	0	7	6508303_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=6508303_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76366501_76391501_114C;SPAN=13664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:66 GQ:5.3 PL:[5.3, 0.0, 153.8] SR:7 DR:0 LR:-5.226 LO:13.76);ALT=T[chr17:76388555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76704345	+	chr17	76705732	+	.	0	11	6509277_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6509277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_76685001_76710001_289C;SPAN=1387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:79 GQ:14.9 PL:[14.9, 0.0, 176.6] SR:11 DR:0 LR:-14.91 LO:23.02);ALT=T[chr17:76705732[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76704389	+	chr17	76778289	+	.	12	0	6509619_1	34.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6509619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76704389(+)-17:76778289(-)__17_76758501_76783501D;SPAN=73900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:20 GQ:14.3 PL:[34.1, 0.0, 14.3] SR:0 DR:12 LR:-34.64 LO:34.64);ALT=T[chr17:76778289[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76970903	+	chr17	76975905	+	TGCCCGAAGGCAGCTCTGCCCAGAGCCTGGGTGGCGTTCTCGAAGCCCAGGGCCCGGCAGACGACGCTGGCATCAGTCAGGTCCCACAGGTTGTCACACACAGTGCCCCACTGGCCTCTGTAGAAGATCTCCACGCGGCCCTGGTTGGTGGCGCCCCCATCGGCCAGCCGCATGTCACCATCGTTCACGCCTTGGGTTCCTGCAACCAGCAGCCACACCCAGAAGAGCCTCGGAGGGGTCATGGCCGTGCCTGGATGCCCAGAT	2	25	6510169_1	51.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTG;INSERTION=TGCCCGAAGGCAGCTCTGCCCAGAGCCTGGGTGGCGTTCTCGAAGCCCAGGGCCCGGCAGACGACGCTGGCATCAGTCAGGTCCCACAGGTTGTCACACACAGTGCCCCACTGGCCTCTGTAGAAGATCTCCACGCGGCCCTGGTTGGTGGCGCCCCCATCGGCCAGCCGCATGTCACCATCGTTCACGCCTTGGGTTCCTGCAACCAGCAGCCACACCCAGAAGAGCCTCGGAGGGGTCATGGCCGTGCCTGGATGCCCAGAT;MAPQ=60;MATEID=6510169_2;MATENM=0;NM=1;NUMPARTS=4;SCTG=c_17_76954501_76979501_140C;SPAN=5002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:115 GQ:51.5 PL:[51.5, 0.0, 226.4] SR:25 DR:2 LR:-51.37 LO:57.69);ALT=T[chr17:76975905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76972290	+	chr17	76975909	+	.	48	0	6510173_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6510173_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76972290(+)-17:76975909(-)__17_76954501_76979501D;SPAN=3619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:89 GQ:81.5 PL:[134.3, 0.0, 81.5] SR:0 DR:48 LR:-135.0 LO:135.0);ALT=C[chr17:76975909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76973299	+	chr17	76975905	+	.	29	17	6510177_1	87.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=6510177_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_17_76954501_76979501_140C;SPAN=2606;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:92 GQ:87.5 PL:[87.5, 0.0, 133.7] SR:17 DR:29 LR:-87.31 LO:87.89);ALT=G[chr17:76975905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	76994019	+	chr17	77005768	+	.	8	0	6510308_1	18.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6510308_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:76994019(+)-17:77005768(-)__17_76979001_77004001D;SPAN=11749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:31 GQ:18.2 PL:[18.2, 0.0, 54.5] SR:0 DR:8 LR:-18.01 LO:19.15);ALT=C[chr17:77005768[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	77393690	+	chr17	77365465	+	.	49	28	6511543_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6511543_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_17_77371001_77396001_104C;SPAN=28225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:51 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:28 DR:49 LR:-181.5 LO:181.5);ALT=]chr17:77393690]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr17	78237577	+	chr17	78247037	+	.	6	14	6514132_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6514132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_78228501_78253501_354C;SPAN=9460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:77 GQ:38.6 PL:[38.6, 0.0, 147.5] SR:14 DR:6 LR:-38.56 LO:42.19);ALT=G[chr17:78247037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	78965787	+	chr17	78968379	+	.	12	0	6516224_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6516224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:78965787(+)-17:78968379(-)__17_78963501_78988501D;SPAN=2592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:47 GQ:26.9 PL:[26.9, 0.0, 86.3] SR:0 DR:12 LR:-26.88 LO:28.66);ALT=G[chr17:78968379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	78965796	+	chr17	78968818	+	.	12	0	6516225_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6516225_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:78965796(+)-17:78968818(-)__17_78963501_78988501D;SPAN=3022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:0 DR:12 LR:-21.19 LO:26.47);ALT=C[chr17:78968818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79213492	+	chr17	79214785	+	.	39	0	6516554_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6516554_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79213492(+)-17:79214785(-)__17_79208501_79233501D;SPAN=1293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:85 GQ:99 PL:[105.8, 0.0, 99.2] SR:0 DR:39 LR:-105.7 LO:105.7);ALT=G[chr17:79214785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79478667	+	chr17	79479765	+	.	17	0	6517690_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6517690_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79478667(+)-17:79479765(-)__17_79478001_79503001D;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:17 DP:838 GQ:99 PL:[0.0, 170.6, 2376.0] SR:0 DR:17 LR:170.9 LO:20.97);ALT=G[chr17:79479765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79618184	+	chr17	79620188	+	TCCCAGGCCTTCCATTCCAGGGATGTCGTCCCCAA	0	17	6517988_1	33.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TCCCAGGCCTTCCATTCCAGGGATGTCGTCCCCAA;MAPQ=60;MATEID=6517988_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_79600501_79625501_333C;SPAN=2004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:84 GQ:33.5 PL:[33.5, 0.0, 168.8] SR:17 DR:0 LR:-33.36 LO:38.63);ALT=T[chr17:79620188[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79649226	+	chr17	79650577	+	.	14	0	6518261_1	35.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=6518261_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79649226(+)-17:79650577(-)__17_79625001_79650001D;SPAN=1351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:38 GQ:35.9 PL:[35.9, 0.0, 55.7] SR:0 DR:14 LR:-35.92 LO:36.17);ALT=C[chr17:79650577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79781235	+	chr17	79791113	+	.	8	0	6518479_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6518479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79781235(+)-17:79791113(-)__17_79772001_79797001D;SPAN=9878;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=C[chr17:79791113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79782317	+	chr17	79791113	+	.	23	0	6518487_1	59.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6518487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79782317(+)-17:79791113(-)__17_79772001_79797001D;SPAN=8796;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:59 GQ:59.9 PL:[59.9, 0.0, 83.0] SR:0 DR:23 LR:-59.94 LO:60.15);ALT=C[chr17:79791113[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79801968	+	chr17	79803019	+	.	2	9	6518614_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6518614_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCATCA;SCTG=c_17_79796501_79821501_216C;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:2 PL:[2.0, 0.0, 158.0] SR:9 DR:2 LR:-1.908 LO:12.99);ALT=C[chr17:79803019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79801968	+	chr17	79803435	+	GTCATCATCCCCTGCCCCATCCTGGCCACCGCTCTCCAGGAATTTCTTAAAACCATCCAGCGTGCGTTCCCCGTTGTAATCAATG	5	15	6518615_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=GTCATCATCCCCTGCCCCATCCTGGCCACCGCTCTCCAGGAATTTCTTAAAACCATCCAGCGTGCGTTCCCCGTTGTAATCAATG;MAPQ=60;MATEID=6518615_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_79796501_79821501_216C;SPAN=1467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:85 GQ:36.5 PL:[36.5, 0.0, 168.5] SR:15 DR:5 LR:-36.39 LO:41.3);ALT=C[chr17:79803435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79813464	+	chr17	79817057	+	.	0	7	6518645_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6518645_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79796501_79821501_284C;SPAN=3593;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:74 GQ:3.2 PL:[3.2, 0.0, 174.8] SR:7 DR:0 LR:-3.059 LO:13.4);ALT=T[chr17:79817057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79827834	+	chr17	79829171	+	.	112	58	6518996_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=6518996_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79821001_79846001_191C;SPAN=1337;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:94 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:58 DR:112 LR:-373.0 LO:373.0);ALT=C[chr17:79829171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79849982	+	chr17	79851427	+	.	129	6	6518761_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6518761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79845501_79870501_198C;SPAN=1445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:81 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:6 DR:129 LR:-399.4 LO:399.4);ALT=G[chr17:79851427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79849998	+	chr17	79857795	+	.	63	0	6518763_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6518763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79849998(+)-17:79857795(-)__17_79845501_79870501D;SPAN=7797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:124 GQ:99 PL:[174.5, 0.0, 125.0] SR:0 DR:63 LR:-174.8 LO:174.8);ALT=T[chr17:79857795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79852463	+	chr17	79857796	+	.	3	83	6518772_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6518772_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_79845501_79870501_146C;SPAN=5333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:161 GQ:99 PL:[237.2, 0.0, 151.4] SR:83 DR:3 LR:-237.9 LO:237.9);ALT=G[chr17:79857796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79935595	+	chr17	79941429	+	.	9	0	6518953_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6518953_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79935595(+)-17:79941429(-)__17_79919001_79944001D;SPAN=5834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:0 DR:9 LR:-7.222 LO:17.79);ALT=A[chr17:79941429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79977306	+	chr17	79980693	+	.	66	0	6519076_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6519076_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79977306(+)-17:79980693(-)__17_79968001_79993001D;SPAN=3387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:83 GQ:4.1 PL:[195.5, 0.0, 4.1] SR:0 DR:66 LR:-206.2 LO:206.2);ALT=C[chr17:79980693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	79977833	+	chr17	79980599	+	.	15	0	6519080_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6519080_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:79977833(+)-17:79980599(-)__17_79968001_79993001D;SPAN=2766;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:51 GQ:35.9 PL:[35.9, 0.0, 85.4] SR:0 DR:15 LR:-35.7 LO:36.92);ALT=A[chr17:79980599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80009877	+	chr17	80011143	+	.	13	0	6519313_1	31.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6519313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80009877(+)-17:80011143(-)__17_79992501_80017501D;SPAN=1266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:44 GQ:31.1 PL:[31.1, 0.0, 74.0] SR:0 DR:13 LR:-30.99 LO:32.03);ALT=C[chr17:80011143[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80009882	+	chr17	80011740	+	.	36	0	6519314_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6519314_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80009882(+)-17:80011740(-)__17_79992501_80017501D;SPAN=1858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:45 GQ:1.1 PL:[106.7, 0.0, 1.1] SR:0 DR:36 LR:-112.7 LO:112.7);ALT=C[chr17:80011740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80059743	+	chr17	80064146	+	.	48	6	6519145_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6519145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80041501_80066501_279C;SPAN=4403;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:78 GQ:41.6 PL:[147.2, 0.0, 41.6] SR:6 DR:48 LR:-150.5 LO:150.5);ALT=C[chr17:80064146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80186459	+	chr17	80193858	+	.	9	0	6519800_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6519800_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80186459(+)-17:80193858(-)__17_80188501_80213501D;SPAN=7399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:22 GQ:23.9 PL:[23.9, 0.0, 27.2] SR:0 DR:9 LR:-23.75 LO:23.78);ALT=G[chr17:80193858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39044999	+	chr17	80313286	+	GAGAATCATTTGAACCTGGGAGGTAGAGGTTGCA	23	60	6811733_1	99.0	.	DISC_MAPQ=0;EVDNC=TSI_G;HOMSEQ=GTGAGCTGAGATCGCGCCATTGCACTCCA;INSERTION=GAGAATCATTTGAACCTGGGAGGTAGAGGTTGCA;MAPQ=34;MATEID=6811733_2;MATENM=2;NM=2;NUMPARTS=3;SCTG=c_19_39028501_39053501_492C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:32 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:60 DR:23 LR:-211.3 LO:211.3);ALT=]chr19:39044999]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr17	80373506	+	chr17	80376288	+	.	0	16	6520241_1	34.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6520241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80360001_80385001_77C;SPAN=2782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:67 GQ:34.7 PL:[34.7, 0.0, 127.1] SR:16 DR:0 LR:-34.66 LO:37.67);ALT=G[chr17:80376288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80402468	+	chr17	80404498	+	CTGGTCGTGGCCAGCTCTGAAAAGAGTCAGCAGCTTCTTGTAGAGGCTGAACGTCTTCAAAACAACCTTCCCTGTGCTCTTGTCGAAGATGGCTT	0	16	6520343_1	29.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=CTGGTCGTGGCCAGCTCTGAAAAGAGTCAGCAGCTTCTTGTAGAGGCTGAACGTCTTCAAAACAACCTTCCCTGTGCTCTTGTCGAAGATGGCTT;MAPQ=60;MATEID=6520343_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_80384501_80409501_145C;SPAN=2030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:86 GQ:29.6 PL:[29.6, 0.0, 178.1] SR:16 DR:0 LR:-29.52 LO:35.7);ALT=C[chr17:80404498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80402736	+	chr17	80408574	+	.	11	0	6520345_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6520345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80402736(+)-17:80408574(-)__17_80384501_80409501D;SPAN=5838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:83 GQ:14 PL:[14.0, 0.0, 185.6] SR:0 DR:11 LR:-13.82 LO:22.76);ALT=G[chr17:80408574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80403884	+	chr17	80408574	+	.	9	0	6520350_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6520350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80403884(+)-17:80408574(-)__17_80384501_80409501D;SPAN=4690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:81 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-7.764 LO:17.89);ALT=C[chr17:80408574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80404574	+	chr17	80407045	+	CCGCTGTAGTAGGCAGCAGCCAGGCCAATCGACAAGATT	0	12	6520353_1	13.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CCGCTGTAGTAGGCAGCAGCCAGGCCAATCGACAAGATT;MAPQ=60;MATEID=6520353_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_17_80384501_80409501_234C;SPAN=2471;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:96 GQ:13.7 PL:[13.7, 0.0, 218.3] SR:12 DR:0 LR:-13.6 LO:24.51);ALT=T[chr17:80407045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80404629	+	chr17	80408574	+	.	8	0	6520354_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6520354_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80404629(+)-17:80408574(-)__17_80384501_80409501D;SPAN=3945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:0 DR:8 LR:-3.379 LO:15.29);ALT=C[chr17:80408574[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80416702	+	chr17	80422160	+	.	11	0	6520584_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6520584_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80416702(+)-17:80422160(-)__17_80409001_80434001D;SPAN=5458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:81 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:0 DR:11 LR:-14.37 LO:22.89);ALT=G[chr17:80422160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80416707	+	chr17	80417865	+	.	6	5	6520585_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=6520585_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80409001_80434001_218C;SPAN=1158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:5 DR:6 LR:-5.818 LO:15.7);ALT=G[chr17:80417865[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80466975	-	chr17	80468705	+	.	9	0	6520868_1	11.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6520868_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80466975(-)-17:80468705(-)__17_80458001_80483001D;SPAN=1730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:68 GQ:11.3 PL:[11.3, 0.0, 153.2] SR:0 DR:9 LR:-11.29 LO:18.62);ALT=[chr17:80468705[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr17	80601900	+	chr17	80606149	+	.	0	9	6521104_1	24.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6521104_2;MATENM=8;NM=2;NUMPARTS=2;SCTG=c_17_80605001_80630001_366C;SPAN=4249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:20 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:9 DR:0 LR:-24.29 LO:24.29);ALT=C[chr17:80606149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80674706	+	chr17	80676778	+	.	8	0	6521445_1	3.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6521445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80674706(+)-17:80676778(-)__17_80654001_80679001D;SPAN=2072;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:0 DR:8 LR:-3.379 LO:15.29);ALT=C[chr17:80676778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80901928	+	chr17	80904755	+	.	0	11	6522166_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6522166_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80899001_80924001_301C;SPAN=2827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:100 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:11 DR:0 LR:-9.219 LO:21.81);ALT=G[chr17:80904755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80963086	+	chr17	80972330	+	.	0	16	6522285_1	34.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6522285_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_17_80948001_80973001_68C;SPAN=9244;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:68 GQ:34.4 PL:[34.4, 0.0, 130.1] SR:16 DR:0 LR:-34.39 LO:37.55);ALT=T[chr17:80972330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80963133	+	chr17	81006368	+	.	9	0	6522286_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6522286_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80963133(+)-17:81006368(-)__17_80948001_80973001D;SPAN=43235;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:31 GQ:21.5 PL:[21.5, 0.0, 51.2] SR:0 DR:9 LR:-21.31 LO:22.09);ALT=C[chr17:81006368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80972443	+	chr17	81006371	+	.	11	0	6522480_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6522480_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80972443(+)-17:81006371(-)__17_80997001_81022001D;SPAN=33928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:40 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:0 DR:11 LR:-25.47 LO:26.69);ALT=G[chr17:81006371[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr17	80993016	+	chr17	81006399	+	.	11	0	6522482_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6522482_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=17:80993016(+)-17:81006399(-)__17_80997001_81022001D;SPAN=13383;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:45 GQ:24.2 PL:[24.2, 0.0, 83.6] SR:0 DR:11 LR:-24.12 LO:26.03);ALT=T[chr17:81006399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	4535387	+	chr18	4536735	+	AAGGT	0	44	6530649_1	99.0	.	EVDNC=ASSMB;INSERTION=AAGGT;MAPQ=60;MATEID=6530649_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_4532501_4557501_200C;SPAN=1348;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:44 DP:21 GQ:11.7 PL:[128.7, 11.7, 0.0] SR:44 DR:0 LR:-128.7 LO:128.7);ALT=G[chr18:4536735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9102815	+	chr19	53727935	-	.	59	0	6862571_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6862571_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:9102815(+)-19:53727935(+)__19_53704001_53729001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:56 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:0 DR:59 LR:-174.9 LO:174.9);ALT=G]chr19:53727935];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr18	9136963	+	chr18	9182379	+	.	10	5	6537355_1	32.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6537355_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_18_9163001_9188001_100C;SPAN=45416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:27 GQ:32.3 PL:[32.3, 0.0, 32.3] SR:5 DR:10 LR:-32.3 LO:32.3);ALT=G[chr18:9182379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9334918	+	chr18	9337190	+	.	9	4	6537520_1	25.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6537520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_9310001_9335001_158C;SPAN=2272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:28 GQ:25.4 PL:[25.4, 0.0, 41.9] SR:4 DR:9 LR:-25.42 LO:25.66);ALT=G[chr18:9337190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9475691	+	chr18	9512986	+	.	41	30	6537869_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=6537869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_9506001_9531001_226C;SPAN=37295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:56 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:30 DR:41 LR:-171.6 LO:171.6);ALT=T[chr18:9512986[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9513287	+	chr18	9516843	+	.	0	20	6537886_1	52.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6537886_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_9506001_9531001_287C;SPAN=3556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:49 GQ:52.7 PL:[52.7, 0.0, 65.9] SR:20 DR:0 LR:-52.75 LO:52.83);ALT=A[chr18:9516843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9914330	+	chr18	9931807	+	.	33	0	6538777_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6538777_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:9914330(+)-18:9931807(-)__18_9922501_9947501D;SPAN=17477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:39 GQ:3.9 PL:[102.3, 3.9, 0.0] SR:0 DR:33 LR:-105.5 LO:105.5);ALT=A[chr18:9931807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	9950591	+	chr18	9954049	+	.	18	0	6538736_1	37.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6538736_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:9950591(+)-18:9954049(-)__18_9947001_9972001D;SPAN=3458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:82 GQ:37.4 PL:[37.4, 0.0, 159.5] SR:0 DR:18 LR:-37.2 LO:41.62);ALT=T[chr18:9954049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	10222280	+	chr18	10223605	+	.	59	46	6539080_1	99.0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=AA;MAPQ=60;MATEID=6539080_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_10216501_10241501_211C;SPAN=1325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:42 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:46 DR:59 LR:-267.4 LO:267.4);ALT=A[chr18:10223605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	20241677	+	chr18	20245966	+	TAG	12	17	6557975_1	82.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=TAG;MAPQ=40;MATEID=6557975_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_20237001_20262001_90C;SPAN=4289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:27 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:17 DR:12 LR:-82.52 LO:82.52);ALT=A[chr18:20245966[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	20970919	-	chr18	20972171	+	.	5	2	6560009_1	9.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GTGGCTCATGCCTGTAATCC;MAPQ=60;MATEID=6560009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_20972001_20997001_26C;SPAN=1252;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:39 GQ:9.2 PL:[9.2, 0.0, 85.1] SR:2 DR:5 LR:-9.24 LO:12.84);ALT=[chr18:20972171[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	21033466	+	chr18	21042926	+	.	0	31	6560196_1	74.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6560196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21021001_21046001_133C;SPAN=9460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:105 GQ:74 PL:[74.0, 0.0, 179.6] SR:31 DR:0 LR:-73.88 LO:76.37);ALT=G[chr18:21042926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21044592	+	chr18	21046097	+	.	3	5	6560234_1	3.0	.	DISC_MAPQ=50;EVDNC=ASDIS;MAPQ=60;MATEID=6560234_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21045501_21070501_252C;SPAN=1505;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:5 DR:3 LR:-3.23 LO:9.742);ALT=T[chr18:21046097[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21059388	+	chr18	21061134	+	.	2	3	6560283_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6560283_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21045501_21070501_69C;SPAN=1746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:70 GQ:5.7 PL:[0.0, 5.7, 181.5] SR:3 DR:2 LR:5.761 LO:6.746);ALT=G[chr18:21061134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21110577	+	chr18	21111587	+	.	0	4	6560483_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6560483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21094501_21119501_119C;SPAN=1010;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:60 GQ:3 PL:[0.0, 3.0, 151.8] SR:4 DR:0 LR:3.051 LO:7.022);ALT=G[chr18:21111587[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21595002	+	chr18	21599819	+	.	0	10	6561751_1	13.0	.	EVDNC=ASSMB;HOMSEQ=TACAG;MAPQ=60;MATEID=6561751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_21584501_21609501_60C;SPAN=4817;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:74 GQ:13.1 PL:[13.1, 0.0, 164.9] SR:10 DR:0 LR:-12.96 LO:20.79);ALT=G[chr18:21599819[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21903397	+	chr18	21904597	+	.	75	0	6562722_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6562722_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:21903397(+)-18:21904597(-)__18_21903001_21928001D;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:182 GQ:99 PL:[198.5, 0.0, 241.4] SR:0 DR:75 LR:-198.3 LO:198.5);ALT=C[chr18:21904597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	21990742	+	chr18	21992048	+	.	68	50	6562677_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=6562677_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_18_21976501_22001501_37C;SPAN=1306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:44 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:50 DR:68 LR:-267.4 LO:267.4);ALT=C[chr18:21992048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	22445942	-	chr18	22922618	+	.	8	0	6564823_1	15.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=6564823_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:22445942(-)-18:22922618(-)__18_22907501_22932501D;SPAN=476676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.57 LO:18.13);ALT=[chr18:22922618[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr18	22446108	+	chr18	22922452	-	.	11	19	6564825_1	78.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=CCACTGCACTCC;MAPQ=60;MATEID=6564825_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_18_22907501_22932501_58C;SPAN=476344;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:41 GQ:18.8 PL:[78.2, 0.0, 18.8] SR:19 DR:11 LR:-79.8 LO:79.8);ALT=C]chr18:22922452];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr18	23827750	+	chr18	23828894	+	.	4	4	6566881_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTGGGAGGCTGAGG;MAPQ=60;MATEID=6566881_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_23814001_23839001_4C;SPAN=1144;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:76 GQ:3.9 PL:[0.0, 3.9, 191.4] SR:4 DR:4 LR:4.085 LO:8.747);ALT=G[chr18:23828894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43591253	+	chr18	43604575	+	GCTGCTTGAAGACTTCAAGGGCCCGCTTCAGGGTG	0	14	6609027_1	26.0	.	DISC_MAPQ=255;EVDNC=TSI_G;INSERTION=GCTGCTTGAAGACTTCAAGGGCCCGCTTCAGGGTG;MAPQ=60;MATEID=6609027_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_43585501_43610501_183C;SPAN=13322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:75 GQ:26 PL:[26.0, 0.0, 154.7] SR:14 DR:0 LR:-25.89 LO:31.26);ALT=T[chr18:43604575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43604698	+	chr18	43652136	+	.	15	0	6609090_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6609090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:43604698(+)-18:43652136(-)__18_43634501_43659501D;SPAN=47438;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:41 GQ:38.6 PL:[38.6, 0.0, 58.4] SR:0 DR:15 LR:-38.41 LO:38.69);ALT=T[chr18:43652136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43620014	+	chr18	43652122	+	.	23	8	6609091_1	71.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6609091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_43634501_43659501_208C;SPAN=32108;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:39 GQ:22.4 PL:[71.9, 0.0, 22.4] SR:8 DR:23 LR:-73.37 LO:73.37);ALT=C[chr18:43652122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43668224	+	chr18	43669531	+	.	0	13	6609456_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=58;MATEID=6609456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_43659001_43684001_137C;SPAN=1307;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:85 GQ:20 PL:[20.0, 0.0, 185.0] SR:13 DR:0 LR:-19.88 LO:27.78);ALT=C[chr18:43669531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43669964	+	chr18	43671647	+	.	17	30	6609462_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6609462_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_43659001_43684001_274C;SPAN=1683;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:73 GQ:53 PL:[122.3, 0.0, 53.0] SR:30 DR:17 LR:-123.5 LO:123.5);ALT=T[chr18:43671647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43671855	+	chr18	43678166	+	.	100	0	6609467_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6609467_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:43671855(+)-18:43678166(-)__18_43659001_43684001D;SPAN=6311;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:100 DP:91 GQ:27 PL:[297.0, 27.0, 0.0] SR:0 DR:100 LR:-297.1 LO:297.1);ALT=T[chr18:43678166[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43675098	+	chr18	43678136	+	.	13	57	6609477_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=36;MATEID=6609477_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_43659001_43684001_105C;SPAN=3038;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:82 GQ:14.3 PL:[182.6, 0.0, 14.3] SR:57 DR:13 LR:-190.6 LO:190.6);ALT=C[chr18:43678136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	43685334	+	chr18	43698145	+	.	0	20	6609262_1	46.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6609262_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_43683501_43708501_36C;SPAN=12811;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:73 GQ:46.4 PL:[46.4, 0.0, 128.9] SR:20 DR:0 LR:-46.24 LO:48.49);ALT=G[chr18:43698145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	44661077	+	chr18	44676748	+	TTTAAGAGCTTCCTGTGCGCCTGGCACAGCTGCATCTTCAATGTGAAGTGTGCCACTGAGATCTACCAAAACAGCTTTTAATGCACGGCATGCTGCCATCCTTCATTC	13	16	6611754_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TTTAAGAGCTTCCTGTGCGCCTGGCACAGCTGCATCTTCAATGTGAAGTGTGCCACTGAGATCTACCAAAACAGCTTTTAATGCACGGCATGCTGCCATCCTTCATTC;MAPQ=60;MATEID=6611754_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_44663501_44688501_282C;SPAN=15671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:46 GQ:50.3 PL:[60.2, 0.0, 50.3] SR:16 DR:13 LR:-60.19 LO:60.19);ALT=T[chr18:44676748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	44662821	+	chr18	44676748	+	.	11	6	6611755_1	37.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=6611755_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=ACAC;SCTG=c_18_44663501_44688501_282C;SPAN=13927;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:46 GQ:37.1 PL:[37.1, 0.0, 73.4] SR:6 DR:11 LR:-37.05 LO:37.75);ALT=C[chr18:44676748[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	44682605	+	chr18	44683807	+	.	0	29	6611896_1	67.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6611896_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TCATCA;SCTG=c_18_44688001_44713001_116C;SPAN=1202;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:29 DP:0 GQ:7.7 PL:[67.6, 7.7, 0.0] SR:29 DR:0 LR:-67.63 LO:67.63);ALT=T[chr18:44683807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	44682629	+	chr18	44702595	+	.	13	0	6611802_1	35.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6611802_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:44682629(+)-18:44702595(-)__18_44663501_44688501D;SPAN=19966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:28 GQ:32 PL:[35.3, 0.0, 32.0] SR:0 DR:13 LR:-35.33 LO:35.33);ALT=T[chr18:44702595[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	44683908	+	chr18	44702558	+	.	0	43	6611807_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6611807_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_44663501_44688501_121C;SPAN=18650;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:43 DP:51 GQ:6.9 PL:[135.3, 6.9, 0.0] SR:43 DR:0 LR:-137.2 LO:137.2);ALT=A[chr18:44702558[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	45423182	+	chr18	45456730	+	.	3	4	6614076_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6614076_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_45447501_45472501_235C;SPAN=33548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:36 GQ:6.8 PL:[6.8, 0.0, 79.4] SR:4 DR:3 LR:-6.752 LO:10.46);ALT=T[chr18:45456730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	46956819	+	chr18	46986766	+	.	0	9	6617845_1	18.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6617845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_46942001_46967001_331C;SPAN=29947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:9 DR:0 LR:-18.33 LO:20.7);ALT=T[chr18:46986766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47008782	+	chr18	47009953	+	.	11	27	6617933_1	90.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6617933_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_46991001_47016001_126C;SPAN=1171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:80 GQ:90.5 PL:[90.5, 0.0, 103.7] SR:27 DR:11 LR:-90.56 LO:90.61);ALT=T[chr18:47009953[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47008832	+	chr18	47013510	+	.	9	0	6617934_1	1.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6617934_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:47008832(+)-18:47013510(-)__18_46991001_47016001D;SPAN=4678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:104 GQ:1.7 PL:[1.7, 0.0, 249.2] SR:0 DR:9 LR:-1.533 LO:16.86);ALT=C[chr18:47013510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47010142	+	chr18	47013413	+	.	0	18	6617940_1	33.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6617940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_46991001_47016001_315C;SPAN=3271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:96 GQ:33.5 PL:[33.5, 0.0, 198.5] SR:18 DR:0 LR:-33.41 LO:40.23);ALT=C[chr18:47013413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47323966	+	chr18	47329057	+	.	0	16	6618683_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=57;MATEID=6618683_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_47309501_47334501_48C;SPAN=5091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:84 GQ:30.2 PL:[30.2, 0.0, 172.1] SR:16 DR:0 LR:-30.06 LO:35.88);ALT=T[chr18:47329057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47323999	+	chr18	47339833	+	.	9	0	6619094_1	19.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=6619094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:47323999(+)-18:47339833(-)__18_47334001_47359001D;SPAN=15834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:38 GQ:19.4 PL:[19.4, 0.0, 72.2] SR:0 DR:9 LR:-19.41 LO:21.15);ALT=C[chr18:47339833[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47329225	+	chr18	47339836	+	.	32	8	6619096_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=6619096_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_47334001_47359001_192C;SPAN=10611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:8 DR:32 LR:-115.5 LO:115.5);ALT=T[chr18:47339836[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	47694973	+	chr18	47698387	+	CTGG	0	39	6619787_1	99.0	.	EVDNC=ASSMB;INSERTION=CTGG;MAPQ=60;MATEID=6619787_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_47677001_47702001_219C;SPAN=3414;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:48 GQ:0.2 PL:[115.7, 0.0, 0.2] SR:39 DR:0 LR:-122.7 LO:122.7);ALT=C[chr18:47698387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	48405680	+	chr18	48422178	+	.	19	17	6621626_1	82.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6621626_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_48387501_48412501_187C;SPAN=16498;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:26 GQ:7.5 PL:[82.5, 7.5, 0.0] SR:17 DR:19 LR:-82.52 LO:82.52);ALT=T[chr18:48422178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	51681684	+	chr18	51686131	+	.	17	5	6628692_1	40.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTACCTG;MAPQ=60;MATEID=6628692_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_51670501_51695501_46C;SPAN=4447;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:72 GQ:40.1 PL:[40.1, 0.0, 132.5] SR:5 DR:17 LR:-39.91 LO:42.8);ALT=G[chr18:51686131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	51952968	+	chr18	51956960	+	.	0	41	6629716_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGCCA;MAPQ=60;MATEID=6629716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_51940001_51965001_206C;SPAN=3992;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:29 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:41 DR:0 LR:-118.8 LO:118.8);ALT=A[chr18:51956960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	52942985	+	chr18	52988899	+	TGCATGAAGAAGGAGCTAGGGAAAGTGCTGGTTGCTGGTTTGGAGGAAGGATAGCCTGGCGAGTCCCTATTGTAGTCGGCAGTGCTTGCTGATGGAGCATAG	0	11	6631369_1	26.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=TGCATGAAGAAGGAGCTAGGGAAAGTGCTGGTTGCTGGTTTGGAGGAAGGATAGCCTGGCGAGTCCCTATTGTAGTCGGCAGTGCTTGCTGATGGAGCATAG;MAPQ=60;MATEID=6631369_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_52969001_52994001_78C;SPAN=45914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:37 GQ:26.3 PL:[26.3, 0.0, 62.6] SR:11 DR:0 LR:-26.29 LO:27.14);ALT=T[chr18:52988899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	54291694	+	chr18	54293591	+	.	0	7	6634355_1	13.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6634355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_54292001_54317001_151C;SPAN=1897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:35 GQ:13.7 PL:[13.7, 0.0, 69.8] SR:7 DR:0 LR:-13.62 LO:15.86);ALT=T[chr18:54293591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	54293689	+	chr18	54305571	+	.	0	26	6634358_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CACC;MAPQ=60;MATEID=6634358_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_54292001_54317001_247C;SPAN=11882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:96 GQ:59.9 PL:[59.9, 0.0, 172.1] SR:26 DR:0 LR:-59.82 LO:62.88);ALT=C[chr18:54305571[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	54946737	+	chr18	54948718	+	.	53	46	6635909_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=6635909_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_18_54929001_54954001_164C;SPAN=1981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:40 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:46 DR:53 LR:-244.3 LO:244.3);ALT=A[chr18:54948718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	55283210	+	chr18	55287800	+	.	0	13	6636607_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CCTT;MAPQ=60;MATEID=6636607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_55272001_55297001_56C;SPAN=4590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:79 GQ:21.5 PL:[21.5, 0.0, 170.0] SR:13 DR:0 LR:-21.51 LO:28.24);ALT=T[chr18:55287800[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	55287885	+	chr18	55288940	+	.	2	3	6636628_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6636628_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_55272001_55297001_364C;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:74 GQ:3.3 PL:[0.0, 3.3, 184.8] SR:3 DR:2 LR:3.543 LO:8.807);ALT=T[chr18:55288940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	56807210	+	chr18	56819765	+	.	8	0	6640951_1	15.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6640951_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:56807210(+)-18:56819765(-)__18_56815501_56840501D;SPAN=12555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:39 GQ:15.8 PL:[15.8, 0.0, 78.5] SR:0 DR:8 LR:-15.84 LO:18.23);ALT=T[chr18:56819765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	56807267	+	chr18	56816741	+	.	20	8	6640952_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAG;MAPQ=60;MATEID=6640952_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_56815501_56840501_166C;SPAN=9474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:43 GQ:41.3 PL:[61.1, 0.0, 41.3] SR:8 DR:20 LR:-61.13 LO:61.13);ALT=G[chr18:56816741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	56816854	+	chr18	56819766	+	.	0	17	6640960_1	35.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6640960_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_56815501_56840501_167C;SPAN=2912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:77 GQ:35.3 PL:[35.3, 0.0, 150.8] SR:17 DR:0 LR:-35.26 LO:39.36);ALT=G[chr18:56819766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	56819917	+	chr18	56825862	+	AGATAATGGAGACATCAAATTTCTGACTAAAGGAGATAATAATGAAGTTGATGATAGAGGCTTGTACAAAGAAGGCCAGAACTGGCTGGAAAAGAAGGACGTGGTGGGAAGAGCAAGAGGGTTTTTACCATATGTTGGTATGGTCACCATAATAATGAATGACTATCCAAAATTCA	0	15	6640973_1	32.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGATAATGGAGACATCAAATTTCTGACTAAAGGAGATAATAATGAAGTTGATGATAGAGGCTTGTACAAAGAAGGCCAGAACTGGCTGGAAAAGAAGGACGTGGTGGGAAGAGCAAGAGGGTTTTTACCATATGTTGGTATGGTCACCATAATAATGAATGACTATCCAAAATTCA;MAPQ=60;MATEID=6640973_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_18_56815501_56840501_103C;SPAN=5945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:15 DR:0 LR:-31.91 LO:35.06);ALT=A[chr18:56825862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	57013284	+	chr18	57016345	+	GGCTCTTTTCCAGGTTCAGTCAACTGGAAAGTCAGAAAAGAAAGGACATCATGGTCAT	3	11	6641420_1	20.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GGCTCTTTTCCAGGTTCAGTCAACTGGAAAGTCAGAAAAGAAAGGACATCATGGTCAT;MAPQ=60;MATEID=6641420_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_57011501_57036501_104C;SPAN=3061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:73 GQ:20 PL:[20.0, 0.0, 155.3] SR:11 DR:3 LR:-19.83 LO:26.06);ALT=C[chr18:57016345[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	57016468	+	chr18	57020430	+	.	0	7	6641429_1	0	.	EVDNC=ASSMB;HOMSEQ=TTAC;MAPQ=60;MATEID=6641429_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_57011501_57036501_181C;SPAN=3962;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:89 GQ:0.9 PL:[0.0, 0.9, 217.8] SR:7 DR:0 LR:1.005 LO:12.81);ALT=C[chr18:57020430[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	57022890	+	chr18	57026263	+	.	0	21	6641445_1	48.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6641445_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_57011501_57036501_221C;SPAN=3373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:77 GQ:48.5 PL:[48.5, 0.0, 137.6] SR:21 DR:0 LR:-48.46 LO:50.87);ALT=T[chr18:57026263[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	57567467	+	chr18	57569876	+	.	34	43	6642667_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6642667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_57550501_57575501_291C;SPAN=2409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:83 GQ:20.6 PL:[179.0, 0.0, 20.6] SR:43 DR:34 LR:-185.9 LO:185.9);ALT=G[chr18:57569876[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	17863746	+	chr18	57777462	+	.	7	55	7209434_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;HOMSEQ=TCAGCCTCCCGAGTAGCTGGGAT;MAPQ=60;MATEID=7209434_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_17860501_17885501_271C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:58 DP:31 GQ:15.6 PL:[171.6, 15.6, 0.0] SR:55 DR:7 LR:-171.6 LO:171.6);ALT=]chr22:17863746]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr18	74092261	+	chr18	74153200	+	.	4	2	6678931_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6678931_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_74137001_74162001_228C;SPAN=60939;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:36 GQ:3.5 PL:[3.5, 0.0, 82.7] SR:2 DR:4 LR:-3.451 LO:7.95);ALT=T[chr18:74153200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	74104825	+	chr18	74106794	+	.	24	0	6678857_1	64.0	.	DISC_MAPQ=34;EVDNC=DSCRD;IMPRECISE;MAPQ=34;MATEID=6678857_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:74104825(+)-18:74106794(-)__18_74088001_74113001D;SPAN=1969;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:56 GQ:64.1 PL:[64.1, 0.0, 70.7] SR:0 DR:24 LR:-64.05 LO:64.08);ALT=G[chr18:74106794[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	74778399	+	chr18	74844663	+	.	8	0	6680916_1	19.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6680916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:74778399(+)-18:74844663(-)__18_74823001_74848001D;SPAN=66264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:25 GQ:19.7 PL:[19.7, 0.0, 39.5] SR:0 DR:8 LR:-19.64 LO:20.05);ALT=A[chr18:74844663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	74817292	+	chr18	74844656	+	.	17	0	6680918_1	49.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6680918_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:74817292(+)-18:74844656(-)__18_74823001_74848001D;SPAN=27364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:24 GQ:6.8 PL:[49.7, 0.0, 6.8] SR:0 DR:17 LR:-51.26 LO:51.26);ALT=T[chr18:74844656[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	75266998	+	chr18	75268160	+	.	59	41	6681908_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6681908_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_75264001_75289001_115C;SPAN=1162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:42 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:41 DR:59 LR:-250.9 LO:250.9);ALT=T[chr18:75268160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76197188	+	chr18	76198342	+	.	13	0	6683961_1	31.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6683961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:76197188(+)-18:76198342(-)__18_76195001_76220001D;SPAN=1154;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:43 GQ:31.4 PL:[31.4, 0.0, 71.0] SR:0 DR:13 LR:-31.26 LO:32.19);ALT=G[chr18:76198342[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76202137	+	chr18	76203341	+	.	45	34	6683978_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAAAGATTGATCAAGG;MAPQ=60;MATEID=6683978_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_18_76195001_76220001_177C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:69 DP:39 GQ:18.6 PL:[204.6, 18.6, 0.0] SR:34 DR:45 LR:-204.7 LO:204.7);ALT=G[chr18:76203341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76290700	+	chr18	76294730	+	.	0	25	6684276_1	72.0	.	EVDNC=ASSMB;HOMSEQ=CTC;MAPQ=60;MATEID=6684276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_76293001_76318001_217C;SPAN=4030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:25 DP:16 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:25 DR:0 LR:-72.62 LO:72.62);ALT=C[chr18:76294730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76295468	+	chr18	76296725	+	.	61	38	6684283_1	99.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=6684283_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_18_76293001_76318001_81C;SPAN=1257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:39 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:38 DR:61 LR:-241.0 LO:241.0);ALT=C[chr18:76296725[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	76728685	+	chr22	50933882	+	.	10	0	7344245_1	24.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7344245_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:76728685(+)-22:50933882(-)__22_50911001_50936001D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:33 GQ:24.2 PL:[24.2, 0.0, 53.9] SR:0 DR:10 LR:-24.07 LO:24.77);ALT=G[chr22:50933882[;VARTYPE=BND:TRX-ht;JOINTYPE=ht
chr18	77309950	+	chr18	77312062	+	.	76	18	6686927_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GACAAAGCCTCACAGACCCCCAGACAGGG;MAPQ=60;MATEID=6686927_2;MATENM=4;NM=0;NUMPARTS=2;SCTG=c_18_77297501_77322501_163C;SPAN=2112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:35 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:18 DR:76 LR:-260.8 LO:260.8);ALT=G[chr18:77312062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	77733858	+	chr18	77748239	+	.	3	4	6687938_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6687938_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_77738501_77763501_232C;SPAN=14381;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:40 GQ:12.2 PL:[12.2, 0.0, 84.8] SR:4 DR:3 LR:-12.27 LO:15.41);ALT=T[chr18:77748239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	77737703	+	chr18	77748238	+	.	0	7	6687940_1	12.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6687940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_18_77738501_77763501_181C;SPAN=10535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:7 DR:0 LR:-12.54 LO:15.5);ALT=T[chr18:77748238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr18	77794653	+	chr18	77797329	+	AAAAAAGGTTTGGTATGAAAGTCCTTCCTTGGGTTCTCACTC	11	15	6687890_1	41.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AAAAAAGGTTTGGTATGAAAGTCCTTCCTTGGGTTCTCACTC;MAPQ=60;MATEID=6687890_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_18_77787501_77812501_275C;SPAN=2676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:80 GQ:41 PL:[41.0, 0.0, 153.2] SR:15 DR:11 LR:-41.05 LO:44.68);ALT=A[chr18:77797329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	481584	+	chr19	480453	+	.	25	0	6690454_1	58.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6690454_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:480453(-)-19:481584(+)__19_465501_490501D;SPAN=1131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:91 GQ:58.1 PL:[58.1, 0.0, 160.4] SR:0 DR:25 LR:-57.87 LO:60.65);ALT=]chr19:481584]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	572701	+	chr19	579502	+	CT	101	22	6690845_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CT;MAPQ=60;MATEID=6690845_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_563501_588501_54C;SPAN=6801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:109 DP:75 GQ:29.4 PL:[323.4, 29.4, 0.0] SR:22 DR:101 LR:-323.5 LO:323.5);ALT=G[chr19:579502[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	572750	+	chr19	580378	+	.	20	0	6690846_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6690846_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:572750(+)-19:580378(-)__19_563501_588501D;SPAN=7628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:71 GQ:47 PL:[47.0, 0.0, 122.9] SR:0 DR:20 LR:-46.78 LO:48.78);ALT=T[chr19:580378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	605301	+	chr19	608432	+	.	18	14	6690637_1	71.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GCTT;MAPQ=60;MATEID=6690637_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_588001_613001_169C;SPAN=3131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:66 GQ:71.3 PL:[71.3, 0.0, 87.8] SR:14 DR:18 LR:-71.25 LO:71.35);ALT=T[chr19:608432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	608623	+	chr19	605529	+	.	18	26	6690639_1	99.0	.	DISC_MAPQ=33;EVDNC=ASDIS;MAPQ=17;MATEID=6690639_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_588001_613001_329C;SPAN=3094;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:67 GQ:47.9 PL:[113.9, 0.0, 47.9] SR:26 DR:18 LR:-115.3 LO:115.3);ALT=]chr19:608623]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	652346	+	chr19	663107	+	.	9	0	6690908_1	24.0	.	DISC_MAPQ=39;EVDNC=DSCRD;IMPRECISE;MAPQ=39;MATEID=6690908_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:652346(+)-19:663107(-)__19_661501_686501D;SPAN=10761;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:21 GQ:24.2 PL:[24.2, 0.0, 24.2] SR:0 DR:9 LR:-24.02 LO:24.03);ALT=C[chr19:663107[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	652885	+	chr19	663046	+	.	13	12	6690909_1	46.0	.	DISC_MAPQ=44;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=6690909_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_19_661501_686501_26C;SPAN=10161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:14 DP:16 GQ:4.2 PL:[46.2, 4.2, 0.0] SR:12 DR:13 LR:-45.42 LO:45.42);ALT=C[chr19:663046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	685923	+	chr19	686924	+	.	17	28	6690973_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6690973_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_661501_686501_249C;SPAN=1001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:62 GQ:39.5 PL:[108.8, 0.0, 39.5] SR:28 DR:17 LR:-110.3 LO:110.3);ALT=C[chr19:686924[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	687189	+	chr19	694814	+	CGCAGCAGGCAGATGTCGTTGGCGTGGGTCATGGGGTGGTAGTCGGGGTGCGTGGTGAGAGCATCGATGCCAAACACCTGCTGGGTGGGCTCCGCAGTACTCAGGACGTGGGCGCCCAGCACCACCAGGCCAGTGCGGAGGTCT	0	176	6691076_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CGCAGCAGGCAGATGTCGTTGGCGTGGGTCATGGGGTGGTAGTCGGGGTGCGTGGTGAGAGCATCGATGCCAAACACCTGCTGGGTGGGCTCCGCAGTACTCAGGACGTGGGCGCCCAGCACCACCAGGCCAGTGCGGAGGTCT;MAPQ=60;MATEID=6691076_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_19_686001_711001_342C;SPAN=7625;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:176 DP:195 GQ:52.6 PL:[577.6, 52.6, 0.0] SR:176 DR:0 LR:-577.6 LO:577.6);ALT=C[chr19:694814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	687189	+	chr19	691858	+	.	27	16	6691075_1	81.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6691075_2;MATENM=1;NM=1;NUMPARTS=3;REPSEQ=GCAGCA;SCTG=c_19_686001_711001_342C;SPAN=4669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:113 GQ:81.5 PL:[81.5, 0.0, 120.5] SR:16 DR:27 LR:-81.27 LO:81.82);ALT=C[chr19:691858[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	687236	+	chr19	695386	+	.	9	0	6691077_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691077_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:687236(+)-19:695386(-)__19_686001_711001D;SPAN=8150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:253 GQ:38.5 PL:[0.0, 38.5, 689.8] SR:0 DR:9 LR:38.84 LO:13.3);ALT=C[chr19:695386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	692005	+	chr19	694814	+	.	8	148	6691098_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6691098_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_686001_711001_342C;SPAN=2809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:153 DP:252 GQ:99 PL:[437.0, 0.0, 172.9] SR:148 DR:8 LR:-442.9 LO:442.9);ALT=G[chr19:694814[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	692052	+	chr19	695350	+	.	110	0	6691099_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691099_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:692052(+)-19:695350(-)__19_686001_711001D;SPAN=3298;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:110 DP:122 GQ:32.7 PL:[359.7, 32.7, 0.0] SR:0 DR:110 LR:-359.8 LO:359.8);ALT=G[chr19:695350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	797540	+	chr19	804030	+	.	19	0	6691587_1	41.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6691587_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:797540(+)-19:804030(-)__19_784001_809001D;SPAN=6490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:78 GQ:41.6 PL:[41.6, 0.0, 147.2] SR:0 DR:19 LR:-41.59 LO:44.92);ALT=C[chr19:804030[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	808763	+	chr19	810543	+	.	2	2	6691364_1	0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6691364_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_808501_833501_26C;SPAN=1780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:68 GQ:5.1 PL:[0.0, 5.1, 174.9] SR:2 DR:2 LR:5.219 LO:6.798);ALT=G[chr19:810543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	828387	+	chr19	829562	+	.	0	162	6691417_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6691417_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_808501_833501_76C;SPAN=1175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:162 DP:201 GQ:5.2 PL:[480.5, 0.0, 5.2] SR:162 DR:0 LR:-508.4 LO:508.4);ALT=G[chr19:829562[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	828432	+	chr19	830704	+	.	12	0	6691418_1	16.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6691418_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:828432(+)-19:830704(-)__19_808501_833501D;SPAN=2272;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:0 DR:12 LR:-16.31 LO:25.12);ALT=G[chr19:830704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	841082	+	chr19	843467	+	.	12	0	6691656_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691656_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:841082(+)-19:843467(-)__19_833001_858001D;SPAN=2385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:0 DR:12 LR:-16.31 LO:25.12);ALT=C[chr19:843467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	861957	+	chr19	863090	+	.	0	94	6691756_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6691756_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_857501_882501_38C;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:94 DP:201 GQ:99 PL:[256.1, 0.0, 229.7] SR:94 DR:0 LR:-255.9 LO:255.9);ALT=G[chr19:863090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	891186	+	chr19	893114	+	.	17	0	6691473_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:891186(+)-19:893114(-)__19_882001_907001D;SPAN=1928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:65 GQ:38.6 PL:[38.6, 0.0, 117.8] SR:0 DR:17 LR:-38.51 LO:40.81);ALT=C[chr19:893114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	902130	+	chr19	913086	+	.	0	14	6691500_1	31.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6691500_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_882001_907001_68C;SPAN=10956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:54 GQ:31.7 PL:[31.7, 0.0, 97.7] SR:14 DR:0 LR:-31.58 LO:33.55);ALT=C[chr19:913086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	902618	+	chr19	913104	+	.	65	0	6691503_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6691503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:902618(+)-19:913104(-)__19_882001_907001D;SPAN=10486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:33 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=C[chr19:913104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	984564	+	chr19	985863	+	.	19	17	6691983_1	76.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6691983_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_19_980001_1005001_42C;SPAN=1299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:85 GQ:76.1 PL:[76.1, 0.0, 128.9] SR:17 DR:19 LR:-76.0 LO:76.78);ALT=G[chr19:985863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	992122	+	chr19	994016	+	.	2	4	6692008_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=6692008_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_980001_1005001_224C;SPAN=1894;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:79 GQ:8.1 PL:[0.0, 8.1, 207.9] SR:4 DR:2 LR:8.199 LO:6.531);ALT=G[chr19:994016[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1026723	+	chr19	1031069	+	.	78	21	6692493_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6692493_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1029001_1054001_204C;SPAN=4346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:40 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:21 DR:78 LR:-250.9 LO:250.9);ALT=G[chr19:1031069[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1026733	+	chr19	1032390	+	.	26	0	6692495_1	75.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6692495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1026733(+)-19:1032390(-)__19_1029001_1054001D;SPAN=5657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:38 GQ:16.1 PL:[75.5, 0.0, 16.1] SR:0 DR:26 LR:-77.64 LO:77.64);ALT=G[chr19:1032390[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1031191	+	chr19	1032391	+	.	0	57	6692496_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6692496_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1029001_1054001_31C;SPAN=1200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:90 GQ:54.8 PL:[163.7, 0.0, 54.8] SR:57 DR:0 LR:-166.8 LO:166.8);ALT=C[chr19:1032391[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1084345	+	chr19	1085657	+	.	2	2	6692319_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6692319_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1078001_1103001_286C;SPAN=1312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:84 GQ:9.3 PL:[0.0, 9.3, 221.1] SR:2 DR:2 LR:9.554 LO:6.423);ALT=G[chr19:1085657[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1091909	+	chr19	1093903	+	.	2	35	6692347_1	93.0	.	DISC_MAPQ=33;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6692347_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1078001_1103001_113C;SPAN=1994;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:107 GQ:93.2 PL:[93.2, 0.0, 165.8] SR:35 DR:2 LR:-93.15 LO:94.29);ALT=G[chr19:1093903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1091930	+	chr19	1095276	+	.	18	0	6692348_1	35.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6692348_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1091930(+)-19:1095276(-)__19_1078001_1103001D;SPAN=3346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:0 DR:18 LR:-35.58 LO:40.99);ALT=C[chr19:1095276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1094082	+	chr19	1095258	+	.	0	14	6692357_1	20.0	.	EVDNC=ASSMB;HOMSEQ=CTGCA;MAPQ=60;MATEID=6692357_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_1078001_1103001_261C;SPAN=1176;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:94 GQ:20.9 PL:[20.9, 0.0, 205.7] SR:14 DR:0 LR:-20.75 LO:29.74);ALT=A[chr19:1095258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1104126	+	chr19	1105184	+	.	173	16	6692418_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6692418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1102501_1127501_158C;SPAN=1058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:184 DP:119 GQ:49.6 PL:[544.6, 49.6, 0.0] SR:16 DR:173 LR:-544.6 LO:544.6);ALT=G[chr19:1105184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1104161	+	chr19	1105653	+	.	13	0	6692419_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6692419_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1104161(+)-19:1105653(-)__19_1102501_1127501D;SPAN=1492;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:75 GQ:22.7 PL:[22.7, 0.0, 158.0] SR:0 DR:13 LR:-22.59 LO:28.56);ALT=A[chr19:1105653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1242608	+	chr19	1244095	+	.	3	102	6693260_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6693260_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_1225001_1250001_147C;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:115 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:102 DR:3 LR:-338.6 LO:338.6);ALT=G[chr19:1244095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1255694	+	chr19	1256999	+	GGAT	4	2	6692800_1	0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=GGAT;MAPQ=60;MATEID=6692800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1249501_1274501_319C;SPAN=1305;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:72 GQ:2.7 PL:[0.0, 2.7, 178.2] SR:2 DR:4 LR:3.002 LO:8.869);ALT=G[chr19:1256999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1269410	+	chr19	1270926	+	.	55	12	6692834_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6692834_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1249501_1274501_58C;SPAN=1516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:94 GQ:53.9 PL:[172.7, 0.0, 53.9] SR:12 DR:55 LR:-175.9 LO:175.9);ALT=G[chr19:1270926[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1269417	+	chr19	1271135	+	.	116	0	6692835_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6692835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1269417(+)-19:1271135(-)__19_1249501_1274501D;SPAN=1718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:127 GQ:34.2 PL:[376.2, 34.2, 0.0] SR:0 DR:116 LR:-376.3 LO:376.3);ALT=C[chr19:1271135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1272052	+	chr19	1274305	+	.	2	16	6692883_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GGT;MAPQ=60;MATEID=6692883_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_19_1274001_1299001_83C;SPAN=2253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:41 GQ:45.2 PL:[45.2, 0.0, 51.8] SR:16 DR:2 LR:-45.01 LO:45.06);ALT=T[chr19:1274305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1275831	+	chr19	1277180	+	.	0	24	6692890_1	54.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=6692890_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1274001_1299001_157C;SPAN=1349;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:90 GQ:54.8 PL:[54.8, 0.0, 163.7] SR:24 DR:0 LR:-54.84 LO:57.85);ALT=T[chr19:1277180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1276104	+	chr19	1277178	+	.	0	7	6692892_1	0	.	EVDNC=ASSMB;HOMSEQ=CCAGGT;MAPQ=60;MATEID=6692892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1274001_1299001_296C;SPAN=1074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:7 DR:0 LR:0.1925 LO:12.92);ALT=T[chr19:1277178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1276121	+	chr19	1278774	+	.	9	0	6692893_1	6.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6692893_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1276121(+)-19:1278774(-)__19_1274001_1299001D;SPAN=2653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:86 GQ:6.5 PL:[6.5, 0.0, 201.2] SR:0 DR:9 LR:-6.41 LO:17.64);ALT=G[chr19:1278774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1277298	+	chr19	1278775	+	.	7	14	6692896_1	46.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6692896_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_1274001_1299001_107C;SPAN=1477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:84 GQ:46.7 PL:[46.7, 0.0, 155.6] SR:14 DR:7 LR:-46.56 LO:49.93);ALT=G[chr19:1278775[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1379243	-	chr19	1380319	+	.	8	0	6693382_1	1.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6693382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1379243(-)-19:1380319(-)__19_1372001_1397001D;SPAN=1076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:0 DR:8 LR:-1.483 LO:15.0);ALT=[chr19:1380319[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	1383993	+	chr19	1388541	+	.	85	0	6693399_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6693399_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1383993(+)-19:1388541(-)__19_1372001_1397001D;SPAN=4548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:120 GQ:43.4 PL:[248.0, 0.0, 43.4] SR:0 DR:85 LR:-256.3 LO:256.3);ALT=G[chr19:1388541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1383995	+	chr19	1390866	+	.	37	0	6693400_1	94.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6693400_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1383995(+)-19:1390866(-)__19_1372001_1397001D;SPAN=6871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:103 GQ:94.4 PL:[94.4, 0.0, 153.8] SR:0 DR:37 LR:-94.23 LO:95.06);ALT=A[chr19:1390866[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1388592	+	chr19	1390869	+	CACCCAGCCTGCCCTGCCAAAGGCCAGAGCCGTGGCTCCCAAACCCAGCAGCCGGGGCGAGTATGTGGTGGCCAAGCTGGATGACCTCGTCAACTGGGCCCGCCG	24	155	6693413_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CACCCAGCCTGCCCTGCCAAAGGCCAGAGCCGTGGCTCCCAAACCCAGCAGCCGGGGCGAGTATGTGGTGGCCAAGCTGGATGACCTCGTCAACTGGGCCCGCCG;MAPQ=60;MATEID=6693413_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_1372001_1397001_146C;SPAN=2277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:166 DP:138 GQ:44.8 PL:[491.8, 44.8, 0.0] SR:155 DR:24 LR:-491.8 LO:491.8);ALT=G[chr19:1390869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1391051	+	chr19	1393239	+	CTACGACCAGATGCCGGAGCCGCGCTACGTGGTCTCCATGGGG	0	48	6693422_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTACGACCAGATGCCGGAGCCGCGCTACGTGGTCTCCATGGGG;MAPQ=60;MATEID=6693422_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_1372001_1397001_17C;SPAN=2188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:115 GQ:99 PL:[127.4, 0.0, 150.5] SR:48 DR:0 LR:-127.3 LO:127.4);ALT=T[chr19:1393239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1391164	+	chr19	1393239	+	.	7	42	6693423_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6693423_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_1372001_1397001_17C;SPAN=2075;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:112 GQ:99 PL:[128.3, 0.0, 141.5] SR:42 DR:7 LR:-128.1 LO:128.2);ALT=G[chr19:1393239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1393330	+	chr19	1395387	+	.	0	91	6693432_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6693432_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1372001_1397001_201C;SPAN=2057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:105 GQ:18.3 PL:[290.4, 18.3, 0.0] SR:91 DR:0 LR:-293.9 LO:293.9);ALT=G[chr19:1395387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1399939	+	chr19	1401294	+	.	0	23	6693293_1	58.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6693293_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1396501_1421501_284C;SPAN=1355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:64 GQ:58.7 PL:[58.7, 0.0, 95.0] SR:23 DR:0 LR:-58.58 LO:59.1);ALT=T[chr19:1401294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1407802	+	chr19	1418201	+	AAGCTCTTCGTGGGCGGTCTTGACTGGAGCACGACCCA	17	29	6693318_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAGCTCTTCGTGGGCGGTCTTGACTGGAGCACGACCCA;MAPQ=60;MATEID=6693318_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_1396501_1421501_23C;SPAN=10399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:79 GQ:90.8 PL:[100.7, 0.0, 90.8] SR:29 DR:17 LR:-100.8 LO:100.8);ALT=G[chr19:1418201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1407802	+	chr19	1417498	+	.	6	19	6693317_1	50.0	.	DISC_MAPQ=50;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6693317_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_19_1396501_1421501_23C;SPAN=9696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:56 GQ:50.9 PL:[50.9, 0.0, 83.9] SR:19 DR:6 LR:-50.85 LO:51.32);ALT=G[chr19:1417498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1432689	+	chr19	1434735	+	.	6	8	6693556_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6693556_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1421001_1446001_39C;SPAN=2046;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:8 DR:6 LR:-16.26 LO:23.36);ALT=G[chr19:1434735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1475259	+	chr19	1478773	+	.	8	10	6693701_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6693701_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1470001_1495001_295C;SPAN=3514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:84 GQ:33.5 PL:[33.5, 0.0, 168.8] SR:10 DR:8 LR:-33.36 LO:38.63);ALT=T[chr19:1478773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1475308	+	chr19	1479117	+	.	15	0	6693702_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6693702_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1475308(+)-19:1479117(-)__19_1470001_1495001D;SPAN=3809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:74 GQ:29.6 PL:[29.6, 0.0, 148.4] SR:0 DR:15 LR:-29.47 LO:34.09);ALT=G[chr19:1479117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1598215	+	chr19	1599409	+	.	0	145	6694009_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=6694009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1592501_1617501_49C;SPAN=1194;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:145 DP:303 GQ:99 PL:[396.7, 0.0, 337.3] SR:145 DR:0 LR:-396.8 LO:396.8);ALT=C[chr19:1599409[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1598263	+	chr19	1605361	+	.	61	0	6694010_1	99.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6694010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:1598263(+)-19:1605361(-)__19_1592501_1617501D;SPAN=7098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:91 GQ:41.6 PL:[176.9, 0.0, 41.6] SR:0 DR:61 LR:-181.2 LO:181.2);ALT=G[chr19:1605361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	1599560	+	chr19	1605358	+	.	75	24	6694017_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6694017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_1592501_1617501_289C;SPAN=5798;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:114 GQ:25.4 PL:[249.8, 0.0, 25.4] SR:24 DR:75 LR:-260.2 LO:260.2);ALT=C[chr19:1605358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2078679	+	chr19	2085172	+	.	2	7	6695954_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6695954_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2082501_2107501_182C;SPAN=6493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:34 GQ:17.3 PL:[17.3, 0.0, 63.5] SR:7 DR:2 LR:-17.2 LO:18.78);ALT=C[chr19:2085172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2234301	+	chr19	2236190	+	.	10	0	6696048_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6696048_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2234301(+)-19:2236190(-)__19_2229501_2254501D;SPAN=1889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:73 GQ:13.4 PL:[13.4, 0.0, 161.9] SR:0 DR:10 LR:-13.23 LO:20.85);ALT=T[chr19:2236190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2236932	+	chr19	2243377	+	.	46	0	6696056_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6696056_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2236932(+)-19:2243377(-)__19_2229501_2254501D;SPAN=6445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:75 GQ:49.1 PL:[131.6, 0.0, 49.1] SR:0 DR:46 LR:-133.5 LO:133.5);ALT=C[chr19:2243377[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2236946	+	chr19	2244540	+	.	11	0	6696057_1	15.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6696057_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2236946(+)-19:2244540(-)__19_2229501_2254501D;SPAN=7594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:76 GQ:15.8 PL:[15.8, 0.0, 167.6] SR:0 DR:11 LR:-15.72 LO:23.22);ALT=G[chr19:2244540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2269743	+	chr19	2271382	+	.	0	202	6696468_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6696468_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2254001_2279001_304C;SPAN=1639;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:202 DP:335 GQ:99 PL:[576.2, 0.0, 236.2] SR:202 DR:0 LR:-583.7 LO:583.7);ALT=G[chr19:2271382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2269744	+	chr19	2271779	+	.	34	4	6696469_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6696469_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2254001_2279001_360C;SPAN=2035;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:216 GQ:99 PL:[109.9, 0.0, 413.6] SR:4 DR:34 LR:-109.8 LO:119.8);ALT=G[chr19:2271779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2270247	+	chr19	2271381	+	.	111	0	6696475_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6696475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2270247(+)-19:2271381(-)__19_2254001_2279001D;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:195 GQ:99 PL:[313.7, 0.0, 158.6] SR:0 DR:111 LR:-316.3 LO:316.3);ALT=G[chr19:2271381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2321823	+	chr19	2324124	+	.	0	71	6696368_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6696368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2303001_2328001_60C;SPAN=2301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:175 GQ:99 PL:[187.1, 0.0, 236.6] SR:71 DR:0 LR:-187.0 LO:187.3);ALT=T[chr19:2324124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2324198	+	chr19	2328386	+	.	0	73	6696586_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTT;MAPQ=60;MATEID=6696586_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2327501_2352501_344C;SPAN=4188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:73 DP:45 GQ:19.5 PL:[214.5, 19.5, 0.0] SR:73 DR:0 LR:-214.6 LO:214.6);ALT=T[chr19:2328386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2328778	+	chr19	2334597	+	.	8	0	6696591_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6696591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2328778(+)-19:2334597(-)__19_2327501_2352501D;SPAN=5819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=A[chr19:2334597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2334720	+	chr19	2337442	+	.	0	10	6696608_1	11.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6696608_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_2327501_2352501_333C;SPAN=2722;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:82 GQ:11 PL:[11.0, 0.0, 185.9] SR:10 DR:0 LR:-10.79 LO:20.31);ALT=A[chr19:2337442[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2349583	+	chr19	2348175	+	.	44	0	6696649_1	99.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6696649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2348175(-)-19:2349583(+)__19_2327501_2352501D;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:73 GQ:49.7 PL:[125.6, 0.0, 49.7] SR:0 DR:44 LR:-127.1 LO:127.1);ALT=]chr19:2349583]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	2737680	+	chr19	2739942	+	.	58	0	6697898_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6697898_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2737680(+)-19:2739942(-)__19_2719501_2744501D;SPAN=2262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:81 GQ:24.5 PL:[169.7, 0.0, 24.5] SR:0 DR:58 LR:-175.4 LO:175.4);ALT=T[chr19:2739942[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2767686	+	chr19	2768967	+	.	0	16	6698087_1	34.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6698087_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_19_2744001_2769001_227C;SPAN=1281;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:68 GQ:34.4 PL:[34.4, 0.0, 130.1] SR:16 DR:0 LR:-34.39 LO:37.55);ALT=T[chr19:2768967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2767735	+	chr19	2783228	+	.	12	0	6698088_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6698088_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2767735(+)-19:2783228(-)__19_2744001_2769001D;SPAN=15493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:16 GQ:2.3 PL:[35.3, 0.0, 2.3] SR:0 DR:12 LR:-36.79 LO:36.79);ALT=A[chr19:2783228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2769087	+	chr19	2783228	+	.	11	0	6698092_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6698092_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2769087(+)-19:2783228(-)__19_2744001_2769001D;SPAN=14141;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:3 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:11 LR:-29.71 LO:29.71);ALT=T[chr19:2783228[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	2785625	+	chr19	2790416	+	.	13	0	6697997_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6697997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:2785625(+)-19:2790416(-)__19_2768501_2793501D;SPAN=4791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:81 GQ:21.2 PL:[21.2, 0.0, 173.0] SR:0 DR:13 LR:-20.97 LO:28.08);ALT=A[chr19:2790416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3054194	+	chr19	3055662	+	.	3	10	6699051_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6699051_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=TT;SCTG=c_19_3038001_3063001_339C;SPAN=1468;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:85 GQ:16.7 PL:[16.7, 0.0, 188.3] SR:10 DR:3 LR:-16.58 LO:25.19);ALT=T[chr19:3055662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3054194	+	chr19	3061158	+	CTTGGGAGAGGTAGGGCAGGACCTGGGCACAAATCCCGTTCAGCCTTTTGACGATCTCAGCCTGTTTGTGCATCTCGATGTTCAAGCCGTAGGACATCTCGTAGTACATCACATAGTGACGCTGCATCTCTGACTTCTCACTGGCCAACTTGTCACATTCGAGCTTGAGG	4	39	6699052_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTTGGGAGAGGTAGGGCAGGACCTGGGCACAAATCCCGTTCAGCCTTTTGACGATCTCAGCCTGTTTGTGCATCTCGATGTTCAAGCCGTAGGACATCTCGTAGTACATCACATAGTGACGCTGCATCTCTGACTTCTCACTGGCCAACTTGTCACATTCGAGCTTGAGG;MAPQ=60;MATEID=6699052_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_19_3038001_3063001_339C;SPAN=6964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:77 GQ:74.9 PL:[111.2, 0.0, 74.9] SR:39 DR:4 LR:-111.5 LO:111.5);ALT=T[chr19:3061158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3057743	+	chr19	3061158	+	.	5	26	6699068_1	79.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6699068_2;MATENM=0;NM=0;NUMPARTS=5;REPSEQ=GG;SCTG=c_19_3038001_3063001_339C;SPAN=3415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:74 GQ:79.1 PL:[79.1, 0.0, 98.9] SR:26 DR:5 LR:-78.98 LO:79.13);ALT=G[chr19:3061158[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3057790	+	chr19	3062195	+	.	9	0	6699070_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6699070_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3057790(+)-19:3062195(-)__19_3038001_3063001D;SPAN=4405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:60 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:0 DR:9 LR:-13.45 LO:19.15);ALT=A[chr19:3062195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3061256	+	chr19	3062697	+	.	7	8	6699654_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6699654_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_3062501_3087501_19C;SPAN=1441;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:10 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:8 DR:7 LR:-29.71 LO:29.71);ALT=C[chr19:3062697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3136594	+	chr19	3148588	+	.	6	5	6699888_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6699888_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3136001_3161001_375C;SPAN=11994;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:5 DR:6 LR:3.123 LO:14.39);ALT=G[chr19:3148588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3148773	+	chr19	3150127	+	.	3	3	6699930_1	0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6699930_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_3136001_3161001_65C;SPAN=1354;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:127 GQ:21 PL:[0.0, 21.0, 349.8] SR:3 DR:3 LR:21.2 LO:5.697);ALT=G[chr19:3150127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3150283	+	chr19	3151705	+	.	3	2	6699939_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6699939_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_3136001_3161001_450C;SPAN=1422;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:2 DR:3 LR:6.844 LO:6.647);ALT=A[chr19:3151705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3151834	+	chr19	3155820	+	.	5	4	6699942_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6699942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3136001_3161001_195C;SPAN=3986;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:78 GQ:5.3 PL:[5.3, 0.0, 183.5] SR:4 DR:5 LR:-5.276 LO:15.61);ALT=G[chr19:3155820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3155950	+	chr19	3157724	+	.	2	7	6699954_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6699954_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3136001_3161001_357C;SPAN=1774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:7 DR:2 LR:-5.326 LO:17.45);ALT=G[chr19:3157724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3157880	+	chr19	3162790	+	.	2	2	6699961_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6699961_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3136001_3161001_416C;SPAN=4910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:46 GQ:0.8 PL:[0.8, 0.0, 109.7] SR:2 DR:2 LR:-0.7415 LO:7.501);ALT=G[chr19:3162790[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3173297	+	chr19	3175785	+	TGCCTGTGCCCCTCATGGGACGCCTGCGTTCTCGTGGGATGCCTGTACCC	9	21	6699496_1	99.0	.	DISC_MAPQ=31;EVDNC=TSI_G;HOMSEQ=GCCTGTGCCCTCATGGGACACCTGTGTTCTCATGGGATGCCTGTGCCCCTCATGGGACGCCTG;INSERTION=TGCCTGTGCCCCTCATGGGACGCCTGCGTTCTCGTGGGATGCCTGTACCC;MAPQ=8;MATEID=6699496_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_19_3160501_3185501_58C;SECONDARY;SPAN=2488;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:34 GQ:9 PL:[99.0, 9.0, 0.0] SR:21 DR:9 LR:-97.74 LO:97.74);ALT=A[chr19:3175785[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3173297	+	chr19	3175777	+	.	9	6	6699495_1	41.0	.	DISC_MAPQ=31;EVDNC=TSI_L;HOMSEQ=CCTGTGTTCTCATGGGA;MAPQ=8;MATEID=6699495_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_3160501_3185501_58C;SPAN=2480;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:30 GQ:31.4 PL:[41.3, 0.0, 31.4] SR:6 DR:9 LR:-41.46 LO:41.46);ALT=A[chr19:3175777[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3186213	+	chr19	3192467	+	.	0	7	6699292_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6699292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3185001_3210001_136C;SPAN=6254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:7 DR:0 LR:-2.246 LO:13.27);ALT=G[chr19:3192467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3359728	+	chr19	3381710	+	.	13	0	6700474_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6700474_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3359728(+)-19:3381710(-)__19_3381001_3406001D;SPAN=21982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:41 GQ:32 PL:[32.0, 0.0, 65.0] SR:0 DR:13 LR:-31.81 LO:32.52);ALT=G[chr19:3381710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3366695	+	chr19	3381724	+	.	16	0	6700475_1	41.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6700475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3366695(+)-19:3381724(-)__19_3381001_3406001D;SPAN=15029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:43 GQ:41.3 PL:[41.3, 0.0, 61.1] SR:0 DR:16 LR:-41.17 LO:41.42);ALT=C[chr19:3381724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3435206	+	chr19	3449010	+	.	3	3	6700555_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6700555_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGAGGA;SCTG=c_19_3430001_3455001_37C;SPAN=13804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:75 GQ:7 PL:[0.0, 7.0, 148.2] SR:3 DR:3 LR:7.309 LO:5.331);ALT=G[chr19:3449010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3456633	+	chr19	3462747	+	.	0	8	6700769_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6700769_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3454501_3479501_319C;SPAN=6114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:63 GQ:9.5 PL:[9.5, 0.0, 141.5] SR:8 DR:0 LR:-9.34 LO:16.4);ALT=G[chr19:3462747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3474996	+	chr19	3478417	+	.	51	6	6700826_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6700826_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_3454501_3479501_216C;SPAN=3421;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:81 GQ:27.8 PL:[166.4, 0.0, 27.8] SR:6 DR:51 LR:-171.5 LO:171.5);ALT=T[chr19:3478417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3475042	+	chr19	3478813	+	.	23	0	6700827_1	54.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6700827_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3475042(+)-19:3478813(-)__19_3454501_3479501D;SPAN=3771;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:80 GQ:54.2 PL:[54.2, 0.0, 140.0] SR:0 DR:23 LR:-54.25 LO:56.34);ALT=C[chr19:3478813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3496916	+	chr19	3500561	+	.	14	0	6700660_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6700660_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3496916(+)-19:3500561(-)__19_3479001_3504001D;SPAN=3645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:0 DR:14 LR:-23.73 LO:30.57);ALT=A[chr19:3500561[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3573045	+	chr19	3574278	+	.	14	0	6701131_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6701131_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3573045(+)-19:3574278(-)__19_3552501_3577501D;SPAN=1233;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:68 GQ:27.8 PL:[27.8, 0.0, 136.7] SR:0 DR:14 LR:-27.79 LO:31.93);ALT=T[chr19:3574278[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3762772	+	chr19	3767257	+	.	8	0	6701649_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6701649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3762772(+)-19:3767257(-)__19_3748501_3773501D;SPAN=4485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=C[chr19:3767257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3762816	+	chr19	3765160	+	.	83	45	6701650_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCAG;MAPQ=60;MATEID=6701650_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_3748501_3773501_150C;SPAN=2344;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:100 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:45 DR:83 LR:-303.7 LO:303.7);ALT=G[chr19:3765160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3765330	+	chr19	3767266	+	CTGTTT	4	36	6701658_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGTTT;MAPQ=60;MATEID=6701658_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3748501_3773501_74C;SPAN=1936;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:99 GQ:98.6 PL:[98.6, 0.0, 141.5] SR:36 DR:4 LR:-98.62 LO:99.04);ALT=G[chr19:3767266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3978172	+	chr19	3979327	+	.	26	30	6702652_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6702652_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_19_3969001_3994001_188C;SPAN=1155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:123 GQ:99 PL:[138.5, 0.0, 158.3] SR:30 DR:26 LR:-138.3 LO:138.4);ALT=T[chr19:3979327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3978172	+	chr19	3979806	+	TGATGGGGATGCAGGCGTGGTCCTCCTCCAGGTCCTTCAGGCAGATCTCCAGGTGCAGCTCGCCGGCGCCCGCGATGATGTGCTCTCCCGACTCCTCGATGATGCA	13	50	6702653_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TGATGGGGATGCAGGCGTGGTCCTCCTCCAGGTCCTTCAGGCAGATCTCCAGGTGCAGCTCGCCGGCGCCCGCGATGATGTGCTCTCCCGACTCCTCGATGATGCA;MAPQ=60;MATEID=6702653_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_3969001_3994001_188C;SPAN=1634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:102 GQ:84.8 PL:[160.7, 0.0, 84.8] SR:50 DR:13 LR:-161.7 LO:161.7);ALT=T[chr19:3979806[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3983336	+	chr19	3985399	+	.	75	0	6702679_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6702679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:3983336(+)-19:3985399(-)__19_3969001_3994001D;SPAN=2063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:245 GQ:99 PL:[181.3, 0.0, 412.4] SR:0 DR:75 LR:-181.2 LO:186.2);ALT=G[chr19:3985399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	3984349	+	chr19	3985372	+	.	161	23	6702686_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TCACC;MAPQ=60;MATEID=6702686_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_3969001_3994001_329C;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:168 DP:110 GQ:45.4 PL:[498.4, 45.4, 0.0] SR:23 DR:161 LR:-498.4 LO:498.4);ALT=C[chr19:3985372[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4179289	+	chr19	4180778	+	.	0	8	6703168_1	0	.	EVDNC=ASSMB;HOMSEQ=CCTGAAG;MAPQ=60;MATEID=6703168_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_4165001_4190001_131C;SPAN=1489;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:116 GQ:4.8 PL:[0.0, 4.8, 290.4] SR:8 DR:0 LR:5.019 LO:14.16);ALT=G[chr19:4180778[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4179330	+	chr19	4182470	+	.	8	0	6703169_1	2.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6703169_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4179330(+)-19:4182470(-)__19_4165001_4190001D;SPAN=3140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:87 GQ:2.9 PL:[2.9, 0.0, 207.5] SR:0 DR:8 LR:-2.838 LO:15.21);ALT=A[chr19:4182470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4180908	+	chr19	4182471	+	.	16	2	6703174_1	29.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6703174_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_4165001_4190001_11C;SPAN=1563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:101 GQ:29 PL:[29.0, 0.0, 213.8] SR:2 DR:16 LR:-28.75 LO:37.11);ALT=T[chr19:4182471[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4448413	+	chr19	4452361	+	.	3	2	6704228_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6704228_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_4434501_4459501_187C;SPAN=3948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:92 GQ:8.1 PL:[0.0, 8.1, 237.6] SR:2 DR:3 LR:8.42 LO:8.321);ALT=C[chr19:4452361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4660015	+	chr19	4670172	+	GTAGGCCATGGCGTACTCAATCTCAGCGCCCCGCACCTCTGCCTTGAACTGTGTGAAGTACAGATAGGACTTCCCCTGGGGCCTCCAGATGGTGCAGGTGAAGTGCTGGTGGTCTTCGCTGGTCCCCAGACTCATCTGCCATTGCTCATTGGTCCCTCCTTGAGAGGCGTAAGTGAACATACACGTATATTTGT	0	94	6704942_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=GTAGGCCATGGCGTACTCAATCTCAGCGCCCCGCACCTCTGCCTTGAACTGTGTGAAGTACAGATAGGACTTCCCCTGGGGCCTCCAGATGGTGCAGGTGAAGTGCTGGTGGTCTTCGCTGGTCCCCAGACTCATCTGCCATTGCTCATTGGTCCCTCCTTGAGAGGCGTAAGTGAACATACACGTATATTTGT;MAPQ=60;MATEID=6704942_2;MATENM=0;NM=0;NUMPARTS=5;SCTG=c_19_4655001_4680001_79C;SPAN=10157;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:81 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:94 DR:0 LR:-277.3 LO:277.3);ALT=A[chr19:4670172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4660812	+	chr19	4670178	+	.	11	0	6704946_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6704946_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4660812(+)-19:4670178(-)__19_4655001_4680001D;SPAN=9366;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:97 GQ:10.1 PL:[10.1, 0.0, 224.6] SR:0 DR:11 LR:-10.03 LO:21.97);ALT=G[chr19:4670178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4665004	+	chr19	4670171	+	.	37	0	6704965_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6704965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4665004(+)-19:4670171(-)__19_4655001_4680001D;SPAN=5167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:80 GQ:93.8 PL:[100.4, 0.0, 93.8] SR:0 DR:37 LR:-100.5 LO:100.5);ALT=C[chr19:4670171[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4666183	-	chr19	4667686	+	.	8	0	6704969_1	8.0	.	DISC_MAPQ=49;EVDNC=DSCRD;IMPRECISE;MAPQ=49;MATEID=6704969_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4666183(-)-19:4667686(-)__19_4655001_4680001D;SPAN=1503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:66 GQ:8.6 PL:[8.6, 0.0, 150.5] SR:0 DR:8 LR:-8.527 LO:16.22);ALT=[chr19:4667686[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	4668715	+	chr19	4670269	+	.	57	0	6704978_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6704978_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4668715(+)-19:4670269(-)__19_4655001_4680001D;SPAN=1554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:75 GQ:12.8 PL:[167.9, 0.0, 12.8] SR:0 DR:57 LR:-175.5 LO:175.5);ALT=A[chr19:4670269[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4818541	+	chr19	4831625	+	.	11	0	6705509_1	26.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6705509_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4818541(+)-19:4831625(-)__19_4826501_4851501D;SPAN=13084;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:0 DR:11 LR:-26.02 LO:26.98);ALT=G[chr19:4831625[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4847903	+	chr19	4852028	+	.	3	2	6705619_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6705619_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_4851001_4876001_246C;SPAN=4125;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:59 GQ:0.5 PL:[0.5, 0.0, 142.4] SR:2 DR:3 LR:-0.5205 LO:9.318);ALT=C[chr19:4852028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4860038	+	chr19	4861341	+	.	7	18	6705651_1	62.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6705651_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_4851001_4876001_265C;SPAN=1303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:76 GQ:62 PL:[62.0, 0.0, 121.4] SR:18 DR:7 LR:-61.94 LO:63.03);ALT=T[chr19:4861341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4860074	+	chr19	4867619	+	.	62	0	6705652_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6705652_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4860074(+)-19:4867619(-)__19_4851001_4876001D;SPAN=7545;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:101 GQ:65.3 PL:[177.5, 0.0, 65.3] SR:0 DR:62 LR:-180.0 LO:180.0);ALT=G[chr19:4867619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	4909596	+	chr19	4910885	+	.	11	0	6705854_1	17.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6705854_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:4909596(+)-19:4910885(-)__19_4900001_4925001D;SPAN=1289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:72 GQ:17 PL:[17.0, 0.0, 155.6] SR:0 DR:11 LR:-16.8 LO:23.5);ALT=C[chr19:4910885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5488255	+	chr19	5487054	+	.	16	5	6707906_1	53.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=GCCCAGGCTGGAGTGCAGTGGCGC;MAPQ=59;MATEID=6707906_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5488001_5513001_76C;SPAN=1201;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:45 GQ:53.9 PL:[53.9, 0.0, 53.9] SR:5 DR:16 LR:-53.83 LO:53.83);ALT=]chr19:5488255]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	5598897	+	chr19	5600140	+	.	3	4	6708235_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6708235_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5586001_5611001_174C;SPAN=1243;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:92 GQ:8.1 PL:[0.0, 8.1, 237.6] SR:4 DR:3 LR:8.42 LO:8.321);ALT=T[chr19:5600140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5600271	+	chr19	5604594	+	.	3	5	6708241_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6708241_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5586001_5611001_45C;SPAN=4323;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:74 GQ:0 PL:[0.0, 0.0, 178.2] SR:5 DR:3 LR:0.2424 LO:11.06);ALT=T[chr19:5604594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5604951	+	chr19	5610004	+	.	0	7	6708254_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCTTC;MAPQ=60;MATEID=6708254_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_5586001_5611001_362C;SPAN=5053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:85 GQ:0.2 PL:[0.2, 0.0, 204.8] SR:7 DR:0 LR:-0.07842 LO:12.95);ALT=C[chr19:5610004[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5621409	+	chr19	5622540	+	.	0	4	6708310_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6708310_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5610501_5635501_355C;SPAN=1131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:88 GQ:10.5 PL:[0.0, 10.5, 234.3] SR:4 DR:0 LR:10.64 LO:6.34);ALT=T[chr19:5622540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5623406	+	chr19	5626414	+	.	5	7	6708315_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6708315_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_5610501_5635501_261C;SPAN=3008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:7 DR:5 LR:-14.86 LO:21.25);ALT=G[chr19:5626414[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5661820	+	chr19	5664032	+	.	2	2	6708511_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6708511_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5659501_5684501_307C;SPAN=2212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:106 GQ:15.3 PL:[0.0, 15.3, 287.1] SR:2 DR:2 LR:15.51 LO:6.013);ALT=G[chr19:5664032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5678709	+	chr19	5680466	+	.	20	0	6708569_1	41.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6708569_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:5678709(+)-19:5680466(-)__19_5659501_5684501D;SPAN=1757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:90 GQ:41.6 PL:[41.6, 0.0, 176.9] SR:0 DR:20 LR:-41.64 LO:46.37);ALT=A[chr19:5680466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5894865	+	chr19	5896464	+	.	9	100	6709400_1	99.0	.	DISC_MAPQ=39;EVDNC=ASDIS;MAPQ=60;MATEID=6709400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5880001_5905001_275C;SPAN=1599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:107 DP:177 GQ:99 PL:[305.3, 0.0, 123.8] SR:100 DR:9 LR:-309.4 LO:309.4);ALT=G[chr19:5896464[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5894913	+	chr19	5903707	+	.	8	0	6709402_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6709402_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:5894913(+)-19:5903707(-)__19_5880001_5905001D;SPAN=8794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:146 GQ:12.9 PL:[0.0, 12.9, 379.5] SR:0 DR:8 LR:13.15 LO:13.34);ALT=A[chr19:5903707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5896795	+	chr19	5903677	+	.	47	0	6709409_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6709409_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:5896795(+)-19:5903677(-)__19_5880001_5905001D;SPAN=6882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:132 GQ:99 PL:[119.6, 0.0, 198.8] SR:0 DR:47 LR:-119.4 LO:120.5);ALT=G[chr19:5903677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5897009	+	chr19	5903622	+	.	0	66	6709411_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6709411_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5880001_5905001_28C;SPAN=6613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:172 GQ:99 PL:[171.5, 0.0, 244.1] SR:66 DR:0 LR:-171.3 LO:172.0);ALT=C[chr19:5903622[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	5978525	+	chr19	5980510	+	.	11	13	6709625_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6709625_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_5978001_6003001_254C;SPAN=1985;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:68 GQ:44.3 PL:[44.3, 0.0, 120.2] SR:13 DR:11 LR:-44.3 LO:46.26);ALT=G[chr19:5980510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6078400	+	chr19	6110432	+	.	13	0	6710036_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6710036_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:6078400(+)-19:6110432(-)__19_6100501_6125501D;SPAN=32032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:0 DR:13 LR:-33.7 LO:33.85);ALT=G[chr19:6110432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6362556	+	chr19	6364462	+	.	0	11	6711074_1	14.0	.	EVDNC=ASSMB;HOMSEQ=GGTG;MAPQ=60;MATEID=6711074_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_6345501_6370501_102C;SPAN=1906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:81 GQ:14.6 PL:[14.6, 0.0, 179.6] SR:11 DR:0 LR:-14.37 LO:22.89);ALT=G[chr19:6364462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6366374	+	chr19	6368548	+	.	2	7	6711098_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6711098_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_6345501_6370501_171C;SPAN=2174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:71 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:7 DR:2 LR:-7.172 LO:15.95);ALT=G[chr19:6368548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6373036	+	chr19	6374213	+	.	67	89	6711229_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6711229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_6370001_6395001_254C;SPAN=1177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:124 DP:137 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:89 DR:67 LR:-406.0 LO:406.0);ALT=G[chr19:6374213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	6381862	+	chr19	6383321	+	.	2	5	6711260_1	0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6711260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_6370001_6395001_21C;SPAN=1459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:77 GQ:0.9 PL:[0.0, 0.9, 188.1] SR:5 DR:2 LR:1.055 LO:10.95);ALT=C[chr19:6383321[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7414403	+	chr19	7427665	+	.	11	0	6714733_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6714733_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7414403(+)-19:7427665(-)__19_7423501_7448501D;SPAN=13262;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:46 GQ:23.9 PL:[23.9, 0.0, 86.6] SR:0 DR:11 LR:-23.85 LO:25.91);ALT=C[chr19:7427665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7429286	+	chr19	7427996	+	.	27	0	6714751_1	64.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6714751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7427996(-)-19:7429286(+)__19_7423501_7448501D;SPAN=1290;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:90 GQ:64.7 PL:[64.7, 0.0, 153.8] SR:0 DR:27 LR:-64.74 LO:66.74);ALT=]chr19:7429286]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	7587667	+	chr19	7589844	+	.	13	6	6715179_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6715179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_7570501_7595501_145C;SPAN=2177;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:107 GQ:20.6 PL:[20.6, 0.0, 238.4] SR:6 DR:13 LR:-20.53 LO:31.44);ALT=G[chr19:7589844[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7694784	+	chr19	7696355	+	.	18	0	6715766_1	39.0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=6715766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7694784(+)-19:7696355(-)__19_7693001_7718001D;SPAN=1571;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:75 GQ:39.2 PL:[39.2, 0.0, 141.5] SR:0 DR:18 LR:-39.1 LO:42.43);ALT=G[chr19:7696355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7702099	+	chr19	7705613	+	.	15	0	6715785_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6715785_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7702099(+)-19:7705613(-)__19_7693001_7718001D;SPAN=3514;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:106 GQ:20.9 PL:[20.9, 0.0, 235.4] SR:0 DR:15 LR:-20.8 LO:31.5);ALT=T[chr19:7705613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7702112	+	chr19	7703898	+	.	28	0	6715786_1	66.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6715786_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7702112(+)-19:7703898(-)__19_7693001_7718001D;SPAN=1786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:95 GQ:66.8 PL:[66.8, 0.0, 162.5] SR:0 DR:28 LR:-66.69 LO:68.95);ALT=G[chr19:7703898[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7702112	+	chr19	7704615	+	.	35	0	6715787_1	91.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6715787_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:7702112(+)-19:7704615(-)__19_7693001_7718001D;SPAN=2503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:90 GQ:91.1 PL:[91.1, 0.0, 127.4] SR:0 DR:35 LR:-91.15 LO:91.48);ALT=G[chr19:7704615[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	7745936	+	chr19	7747126	+	.	115	7	6715859_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6715859_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_7742001_7767001_141C;SPAN=1190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:118 DP:120 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:7 DR:115 LR:-356.5 LO:356.5);ALT=G[chr19:7747126[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8046073	+	chr19	8070379	+	CTACTTTATCCCGAATAAGTTTTGCAGATTCAACTTCACCAATGCTGCTGAACAGGCTTCGTAACTCATCCTGGGTCATGTTCTGAGGGAGGTAGTTGACGATCAAATTCGTTCTCCCGATGTCACCCCTGCAGTCTTCGGCCATGTGGTCTTCATAACCATTAGACATTGTATTTTTCAAAAAT	0	33	6717079_1	95.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=CTACTTTATCCCGAATAAGTTTTGCAGATTCAACTTCACCAATGCTGCTGAACAGGCTTCGTAACTCATCCTGGGTCATGTTCTGAGGGAGGTAGTTGACGATCAAATTCGTTCTCCCGATGTCACCCCTGCAGTCTTCGGCCATGTGGTCTTCATAACCATTAGACATTGTATTTTTCAAAAAT;MAPQ=60;MATEID=6717079_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8060501_8085501_245C;SPAN=24306;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:6 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:33 DR:0 LR:-95.72 LO:95.72);ALT=G[chr19:8070379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8056718	+	chr19	8070379	+	.	52	20	6717081_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6717081_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8060501_8085501_245C;SPAN=13661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:61 DP:6 GQ:16.2 PL:[178.2, 16.2, 0.0] SR:20 DR:52 LR:-178.2 LO:178.2);ALT=G[chr19:8070379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8376481	+	chr19	8381380	+	.	2	73	6718251_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6718251_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8379001_8404001_307C;SPAN=4899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:74 DP:68 GQ:19.8 PL:[217.8, 19.8, 0.0] SR:73 DR:2 LR:-217.9 LO:217.9);ALT=T[chr19:8381380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8376524	+	chr19	8386191	+	.	18	0	6718252_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6718252_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:8376524(+)-19:8386191(-)__19_8379001_8404001D;SPAN=9667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:44 GQ:47.6 PL:[47.6, 0.0, 57.5] SR:0 DR:18 LR:-47.5 LO:47.57);ALT=T[chr19:8386191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8381530	+	chr19	8386192	+	GCTTGGAGATCTCCTGGTAGCGTAGCTGCAGCTTCCCCTGCAGGTCATG	74	28	6718260_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GCTTGGAGATCTCCTGGTAGCGTAGCTGCAGCTTCCCCTGCAGGTCATG;MAPQ=60;MATEID=6718260_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8379001_8404001_277C;SPAN=4662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:99 GQ:6.9 PL:[254.1, 6.9, 0.0] SR:28 DR:74 LR:-264.3 LO:264.3);ALT=C[chr19:8386192[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8455340	+	chr19	8464745	+	.	85	4	6718532_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6718532_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8452501_8477501_184C;SPAN=9405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:94 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:4 DR:85 LR:-277.3 LO:277.3);ALT=G[chr19:8464745[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8455378	+	chr19	8466969	+	.	15	0	6718533_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6718533_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:8455378(+)-19:8466969(-)__19_8452501_8477501D;SPAN=11591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:89 GQ:25.4 PL:[25.4, 0.0, 190.4] SR:0 DR:15 LR:-25.4 LO:32.75);ALT=G[chr19:8466969[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8464944	+	chr19	8466970	+	.	0	32	6718564_1	76.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6718564_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8452501_8477501_93C;SPAN=2026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:108 GQ:76.4 PL:[76.4, 0.0, 185.3] SR:32 DR:0 LR:-76.37 LO:78.89);ALT=T[chr19:8466970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8509995	+	chr19	8520288	+	.	41	16	6718641_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6718641_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8501501_8526501_363C;SPAN=10293;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:89 GQ:88.1 PL:[127.7, 0.0, 88.1] SR:16 DR:41 LR:-128.1 LO:128.1);ALT=G[chr19:8520288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8520458	+	chr19	8528477	+	TTGGTGAGGTAACATACGTGGAGCTCTTAATGGACGCTGAAGGAAAGTCAAGGGGATGTGC	8	34	6718695_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTGGTGAGGTAACATACGTGGAGCTCTTAATGGACGCTGAAGGAAAGTCAAGGGGATGTGC;MAPQ=60;MATEID=6718695_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8526001_8551001_306C;SPAN=8019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:53 GQ:18.8 PL:[107.9, 0.0, 18.8] SR:34 DR:8 LR:-111.1 LO:111.1);ALT=G[chr19:8528477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8520458	+	chr19	8527411	+	.	6	21	6718694_1	64.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6718694_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8526001_8551001_306C;SPAN=6953;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:42 GQ:35 PL:[64.7, 0.0, 35.0] SR:21 DR:6 LR:-64.93 LO:64.93);ALT=G[chr19:8527411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8528571	+	chr19	8531119	+	ATTTGCTACAAATACTGTGCTTCCAAGTCTTCCAGCCTGTAATGCATGGATAATCTCATTTGGGATGTTGGGATTATTTAGGATACTGGGTGGGATAGTAATCATTCCTGGGCCACCTGGTCCCATACCCATCCCACCAGTCGTAGCCATCACCTTTTGCATTGCTCTCCTGGCATGTTCACCATCAGGAT	5	12	6718703_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=ATTTGCTACAAATACTGTGCTTCCAAGTCTTCCAGCCTGTAATGCATGGATAATCTCATTTGGGATGTTGGGATTATTTAGGATACTGGGTGGGATAGTAATCATTCCTGGGCCACCTGGTCCCATACCCATCCCACCAGTCGTAGCCATCACCTTTTGCATTGCTCTCCTGGCATGTTCACCATCAGGAT;MAPQ=60;MATEID=6718703_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_8526001_8551001_394C;SPAN=2548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:89 GQ:18.8 PL:[18.8, 0.0, 197.0] SR:12 DR:5 LR:-18.8 LO:27.5);ALT=G[chr19:8531119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8531272	+	chr19	8532419	+	.	2	11	6718714_1	15.0	.	DISC_MAPQ=49;EVDNC=TSI_L;MAPQ=60;MATEID=6718714_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TATA;SCTG=c_19_8526001_8551001_187C;SPAN=1147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:11 DR:2 LR:-15.23 LO:24.87);ALT=T[chr19:8532419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8531272	+	chr19	8536210	+	CTATGTTCAATGGCCAGCTGCTATTTGATAGACCAATGCACGTCAAGATGGATGAGAGGGCCTTACCAAAAGGAGATTTCTTCCCTCCTGAGCGTCCACAACAACTTCCCC	5	21	6718715_1	54.0	.	DISC_MAPQ=43;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=CTATGTTCAATGGCCAGCTGCTATTTGATAGACCAATGCACGTCAAGATGGATGAGAGGGCCTTACCAAAAGGAGATTTCTTCCCTCCTGAGCGTCCACAACAACTTCCCC;MAPQ=60;MATEID=6718715_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_8526001_8551001_187C;SPAN=4938;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:78 GQ:54.8 PL:[54.8, 0.0, 134.0] SR:21 DR:5 LR:-54.79 LO:56.65);ALT=T[chr19:8536210[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8539181	+	chr19	8550484	+	.	9	0	6718888_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6718888_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:8539181(+)-19:8550484(-)__19_8550501_8575501D;SPAN=11303;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:36 GQ:20 PL:[20.0, 0.0, 66.2] SR:0 DR:9 LR:-19.96 LO:21.4);ALT=T[chr19:8550484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8564665	+	chr19	8567448	+	.	53	4	6718945_1	99.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6718945_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_8550501_8575501_130C;SPAN=2783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:106 GQ:99 PL:[152.9, 0.0, 103.4] SR:4 DR:53 LR:-153.3 LO:153.3);ALT=C[chr19:8567448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8592369	+	chr19	8595080	+	.	3	6	6718855_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6718855_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8575001_8600001_319C;SPAN=2711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:95 GQ:2.4 PL:[0.0, 2.4, 234.3] SR:6 DR:3 LR:2.631 LO:12.6);ALT=T[chr19:8595080[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8595458	+	chr19	8601136	+	.	2	2	6718860_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6718860_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_8575001_8600001_6C;SPAN=5678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:40 GQ:2.3 PL:[2.3, 0.0, 94.7] SR:2 DR:2 LR:-2.367 LO:7.756);ALT=C[chr19:8601136[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8619675	+	chr19	8642234	+	.	12	0	6719435_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6719435_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:8619675(+)-19:8642234(-)__19_8599501_8624501D;SPAN=22559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:49 GQ:26.3 PL:[26.3, 0.0, 92.3] SR:0 DR:12 LR:-26.34 LO:28.41);ALT=C[chr19:8642234[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	8620712	+	chr19	8642224	+	.	24	0	6719437_1	70.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6719437_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:8620712(+)-19:8642224(-)__19_8599501_8624501D;SPAN=21512;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:32 GQ:4.7 PL:[70.7, 0.0, 4.7] SR:0 DR:24 LR:-73.59 LO:73.59);ALT=C[chr19:8642224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9274508	+	chr19	9042090	+	.	36	0	6721691_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6721691_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:9042090(-)-19:9274508(+)__19_9261001_9286001D;SPAN=232418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:36 DP:16 GQ:9.6 PL:[105.6, 9.6, 0.0] SR:0 DR:36 LR:-105.6 LO:105.6);ALT=]chr19:9274508]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	9042204	+	chr19	9284364	+	.	9	53	6721693_1	99.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6721693_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_19_9261001_9286001_246C;SPAN=242160;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:20 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:53 DR:9 LR:-161.7 LO:161.7);ALT=A[chr19:9284364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9222962	+	chr19	9225122	+	.	22	21	6722817_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CATGCCTGTAATCCCAGC;MAPQ=60;MATEID=6722817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_9212001_9237001_96C;SPAN=2160;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:68 GQ:47.6 PL:[116.9, 0.0, 47.6] SR:21 DR:22 LR:-118.5 LO:118.5);ALT=C[chr19:9225122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9274510	+	chr19	9284364	+	CATCTGCCACCATGCCCGGCTAATTTTTTTGTGTATTTTTAGTA	17	74	6721726_1	99.0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=GAGA;INSERTION=CATCTGCCACCATGCCCGGCTAATTTTTTTGTGTATTTTTAGTA;MAPQ=0;MATEID=6721726_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_19_9261001_9286001_246C;SECONDARY;SPAN=9854;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:36 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:74 DR:17 LR:-244.3 LO:244.3);ALT=G[chr19:9284364[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9925250	-	chr19	9926301	+	.	8	0	6725282_1	7.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=6725282_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:9925250(-)-19:9926301(-)__19_9922501_9947501D;SPAN=1051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.443 LO:16.0);ALT=[chr19:9926301[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	9938694	+	chr19	9940639	+	.	21	0	6725322_1	43.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6725322_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:9938694(+)-19:9940639(-)__19_9922501_9947501D;SPAN=1945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:97 GQ:43.1 PL:[43.1, 0.0, 191.6] SR:0 DR:21 LR:-43.04 LO:48.41);ALT=A[chr19:9940639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9946079	+	chr19	9949109	+	.	97	4	6725345_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6725345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_9922501_9947501_61C;SPAN=3030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:54 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:4 DR:97 LR:-290.5 LO:290.5);ALT=G[chr19:9949109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9946094	+	chr19	9958704	+	.	8	0	6725346_1	11.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6725346_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:9946094(+)-19:9958704(-)__19_9922501_9947501D;SPAN=12610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:0 DR:8 LR:-11.51 LO:16.91);ALT=G[chr19:9958704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	9949325	+	chr19	9958705	+	.	2	34	6725192_1	86.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6725192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_9947001_9972001_121C;SPAN=9380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:107 GQ:86.6 PL:[86.6, 0.0, 172.4] SR:34 DR:2 LR:-86.55 LO:88.13);ALT=G[chr19:9958705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10227866	+	chr19	10229344	+	.	5	25	6726420_1	39.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6726420_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCTCCT;SCTG=c_19_10216501_10241501_325C;SPAN=1478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:113 GQ:39.9 PL:[39.9, 0.0, 162.1] SR:25 DR:5 LR:-39.64 LO:44.75);ALT=T[chr19:10229344[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10227866	+	chr19	10229544	+	TCCTCCTTGCGACAGCCTTTGAAGCCTTCCGGGTCTCAATCCTGAAGGTGCGGACAAT	9	104	6726421_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TCCTCCTTGCGACAGCCTTTGAAGCCTTCCGGGTCTCAATCCTGAAGGTGCGGACAAT;MAPQ=60;MATEID=6726421_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_10216501_10241501_325C;SPAN=1678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:112 DP:115 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:104 DR:9 LR:-340.0 LO:340.0);ALT=T[chr19:10229544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10227917	+	chr19	10230515	+	.	15	0	6726422_1	8.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6726422_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10227917(+)-19:10230515(-)__19_10216501_10241501D;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:150 GQ:8.9 PL:[8.9, 0.0, 355.4] SR:0 DR:15 LR:-8.876 LO:29.09);ALT=C[chr19:10230515[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10229453	+	chr19	10230513	+	.	35	0	6726433_1	80.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6726433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10229453(+)-19:10230513(-)__19_10216501_10241501D;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:132 GQ:80 PL:[80.0, 0.0, 238.4] SR:0 DR:35 LR:-79.77 LO:84.27);ALT=C[chr19:10230513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10277361	+	chr19	10283765	+	GGTTCTTTGGTTTGACTTCGGAGTCTCTTTTCTT	0	16	6726520_1	32.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGTTCTTTGGTTTGACTTCGGAGTCTCTTTTCTT;MAPQ=60;MATEID=6726520_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_10265501_10290501_70C;SPAN=6404;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:77 GQ:32 PL:[32.0, 0.0, 154.1] SR:16 DR:0 LR:-31.96 LO:36.56);ALT=T[chr19:10283765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10283851	+	chr19	10287968	+	GTTCTCTGGATGTAACTCTACGTCTCTTCTCATCCTGGTCTTTGTCTTCTTCCTTGATGGACTCATCCGATTTGGCTCTTTCAGACTCTTCCTGAGGTTTCCGTTTGGCAGGG	0	63	6726545_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GTTCTCTGGATGTAACTCTACGTCTCTTCTCATCCTGGTCTTTGTCTTCTTCCTTGATGGACTCATCCGATTTGGCTCTTTCAGACTCTTCCTGAGGTTTCCGTTTGGCAGGG;MAPQ=60;MATEID=6726545_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_10265501_10290501_109C;SPAN=4117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:97 GQ:53 PL:[181.7, 0.0, 53.0] SR:63 DR:0 LR:-185.5 LO:185.5);ALT=C[chr19:10287968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10288043	+	chr19	10291026	+	.	0	25	6726557_1	68.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6726557_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10265501_10290501_348C;SPAN=2983;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:53 GQ:58.4 PL:[68.3, 0.0, 58.4] SR:25 DR:0 LR:-68.19 LO:68.19);ALT=G[chr19:10291026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10291618	+	chr19	10305517	+	.	70	0	6726615_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6726615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10291618(+)-19:10305517(-)__19_10290001_10315001D;SPAN=13899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:89 GQ:8.9 PL:[206.9, 0.0, 8.9] SR:0 DR:70 LR:-217.9 LO:217.9);ALT=A[chr19:10305517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10381896	+	chr19	10385438	+	.	9	0	6727189_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6727189_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10381896(+)-19:10385438(-)__19_10363501_10388501D;SPAN=3542;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:74 GQ:9.8 PL:[9.8, 0.0, 168.2] SR:0 DR:9 LR:-9.661 LO:18.26);ALT=T[chr19:10385438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10446652	+	chr19	10449357	+	.	0	9	6727343_1	11.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6727343_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_10437001_10462001_86C;SPAN=2705;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:9 DR:0 LR:-11.02 LO:18.56);ALT=C[chr19:10449357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10446700	+	chr19	10450235	+	.	8	0	6727344_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6727344_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10446700(+)-19:10450235(-)__19_10437001_10462001D;SPAN=3535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:111 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.665 LO:14.32);ALT=C[chr19:10450235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10461839	+	chr19	10463110	+	.	3	2	6727414_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6727414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10437001_10462001_232C;SPAN=1271;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:38 GQ:6.2 PL:[6.2, 0.0, 85.4] SR:2 DR:3 LR:-6.21 LO:10.33);ALT=C[chr19:10463110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10504147	+	chr19	10505707	+	.	13	0	6727683_1	19.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6727683_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10504147(+)-19:10505707(-)__19_10486001_10511001D;SPAN=1560;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:0 DR:13 LR:-19.34 LO:27.64);ALT=C[chr19:10505707[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10506882	+	chr19	10514053	+	.	144	67	6727689_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6727689_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10486001_10511001_172C;SPAN=7171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:178 DP:60 GQ:48.1 PL:[528.1, 48.1, 0.0] SR:67 DR:144 LR:-528.1 LO:528.1);ALT=G[chr19:10514053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10610789	+	chr19	10613947	+	.	8	0	6727726_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6727726_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10610789(+)-19:10613947(-)__19_10608501_10633501D;SPAN=3158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:74 GQ:6.5 PL:[6.5, 0.0, 171.5] SR:0 DR:8 LR:-6.36 LO:15.8);ALT=G[chr19:10613947[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10678096	+	chr19	10679187	+	.	7	8	6728186_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=6728186_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10657501_10682501_353C;SPAN=1091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:95 GQ:7.4 PL:[7.4, 0.0, 221.9] SR:8 DR:7 LR:-7.272 LO:19.63);ALT=G[chr19:10679187[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10765135	+	chr19	10781233	+	.	21	0	6728496_1	52.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6728496_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:10765135(+)-19:10781233(-)__19_10780001_10805001D;SPAN=16098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:62 GQ:52.7 PL:[52.7, 0.0, 95.6] SR:0 DR:21 LR:-52.52 LO:53.28);ALT=C[chr19:10781233[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10765163	+	chr19	10781649	+	AGTTGAAGTATTGATAACACCAAGGAACTCTATCACAATTTGAAAAGATAAGCAAAAGTTTGATTTCCAGACACTACAGAAGAAGTAAAAAT	0	57	6728597_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AGTTGAAGTATTGATAACACCAAGGAACTCTATCACAATTTGAAAAGATAAGCAAAAGTTTGATTTCCAGACACTACAGAAGAAGTAAAAAT;MAPQ=60;MATEID=6728597_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_10755501_10780501_233C;SPAN=16486;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:57 DP:26 GQ:15.3 PL:[168.3, 15.3, 0.0] SR:57 DR:0 LR:-168.3 LO:168.3);ALT=G[chr19:10781649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	10959216	+	chr19	10960934	+	.	6	6	6729202_1	7.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6729202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_10951501_10976501_233C;SPAN=1718;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:6 DR:6 LR:-6.951 LO:17.74);ALT=G[chr19:10960934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11071851	+	chr19	11094799	+	.	19	8	6729967_1	63.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6729967_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11049501_11074501_25C;SPAN=22948;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:34 GQ:17.3 PL:[63.5, 0.0, 17.3] SR:8 DR:19 LR:-64.73 LO:64.73);ALT=G[chr19:11094799[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11100119	+	chr19	11101823	+	.	2	4	6729671_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6729671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11098501_11123501_292C;SPAN=1704;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:87 GQ:3.6 PL:[0.0, 3.6, 217.8] SR:4 DR:2 LR:3.764 LO:10.62);ALT=G[chr19:11101823[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11102000	+	chr19	11105501	+	.	3	5	6729679_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6729679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11098501_11123501_120C;SPAN=3501;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:5 DR:3 LR:0.4634 LO:12.88);ALT=G[chr19:11105501[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11105678	+	chr19	11106888	+	.	4	16	6729692_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6729692_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11098501_11123501_180C;SPAN=1210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:100 GQ:38.9 PL:[38.9, 0.0, 203.9] SR:16 DR:4 LR:-38.93 LO:45.33);ALT=G[chr19:11106888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11170864	+	chr19	11172458	+	.	4	8	6729989_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6729989_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11172001_11197001_318C;SPAN=1594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:59 GQ:17 PL:[17.0, 0.0, 125.9] SR:8 DR:4 LR:-17.03 LO:21.86);ALT=G[chr19:11172458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11448186	+	chr19	11450195	+	.	10	0	6730841_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6730841_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:11448186(+)-19:11450195(-)__19_11441501_11466501D;SPAN=2009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.75 LO:21.78);ALT=T[chr19:11450195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11453801	+	chr19	11455928	+	.	7	17	6730860_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGGC;MAPQ=60;MATEID=6730860_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11441501_11466501_87C;SPAN=2127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:115 GQ:48.2 PL:[48.2, 0.0, 229.7] SR:17 DR:7 LR:-48.07 LO:54.89);ALT=C[chr19:11455928[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11457331	+	chr19	11460611	+	.	28	0	6730873_1	69.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6730873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:11457331(+)-19:11460611(-)__19_11441501_11466501D;SPAN=3280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:85 GQ:69.5 PL:[69.5, 0.0, 135.5] SR:0 DR:28 LR:-69.4 LO:70.61);ALT=T[chr19:11460611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11547327	+	chr19	11548694	+	.	0	6	6731342_1	0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6731342_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11539501_11564501_197C;SPAN=1367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:93 GQ:5.1 PL:[0.0, 5.1, 234.3] SR:6 DR:0 LR:5.39 LO:10.44);ALT=G[chr19:11548694[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11560243	+	chr19	11561459	+	.	8	16	6731379_1	45.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6731379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11539501_11564501_60C;SPAN=1216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:77 GQ:45.2 PL:[45.2, 0.0, 140.9] SR:16 DR:8 LR:-45.16 LO:47.94);ALT=G[chr19:11561459[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11625039	+	chr19	11629888	+	.	0	14	6731810_1	18.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=6731810_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_11613001_11638001_259C;SPAN=4849;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:104 GQ:18.2 PL:[18.2, 0.0, 232.7] SR:14 DR:0 LR:-18.04 LO:29.08);ALT=G[chr19:11629888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11625085	+	chr19	11639874	+	.	18	0	6731811_1	46.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6731811_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:11625085(+)-19:11639874(-)__19_11613001_11638001D;SPAN=14789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:47 GQ:46.7 PL:[46.7, 0.0, 66.5] SR:0 DR:18 LR:-46.68 LO:46.89);ALT=G[chr19:11639874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11630040	+	chr19	11639881	+	.	11	0	6731829_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6731829_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:11630040(+)-19:11639881(-)__19_11613001_11638001D;SPAN=9841;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:0 DR:11 LR:-20.87 LO:24.74);ALT=G[chr19:11639881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	11664943	+	chr19	11670004	+	.	9	0	6731965_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6731965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:11664943(+)-19:11670004(-)__19_11662001_11687001D;SPAN=5061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=C[chr19:11670004[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12098639	+	chr19	12112588	+	.	10	10	6733244_1	43.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6733244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12078501_12103501_6C;SPAN=13949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:47 GQ:43.4 PL:[43.4, 0.0, 69.8] SR:10 DR:10 LR:-43.38 LO:43.74);ALT=G[chr19:12112588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12098639	+	chr19	12114205	+	AAATAAATGGAAAGACCAGAATATTGAAGATCACTACAGAAATCTA	14	22	6733569_1	85.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGGGTCAGGCATGGTGGCTCACACCTGTAATCCCAGCACTTTGGGA;INSERTION=AAATAAATGGAAAGACCAGAATATTGAAGATCACTACAGAAATCTA;MAPQ=60;MATEID=6733569_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_12103001_12128001_254C;SECONDARY;SPAN=15566;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:37 GQ:3.2 PL:[85.7, 0.0, 3.2] SR:22 DR:14 LR:-90.16 LO:90.16);ALT=G[chr19:12114205[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77359862	+	chr19	12670380	+	.	134	0	7455522_1	99.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=7455522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12670380(-)-23:77359862(+)__23_77346501_77371501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:134 DP:50 GQ:36 PL:[396.0, 36.0, 0.0] SR:0 DR:134 LR:-396.1 LO:396.1);ALT=]chrX:77359862]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	12694884	+	chr19	12698931	+	.	89	76	6735358_1	99.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=GCCTCCCA;MAPQ=0;MATEID=6735358_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12691001_12716001_27C;SPAN=4047;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:32 GQ:37.9 PL:[415.9, 37.9, 0.0] SR:76 DR:89 LR:-415.9 LO:415.9);ALT=A[chr19:12698931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12761038	+	chr19	12762967	+	.	11	10	6735746_1	43.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6735746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12740001_12765001_202C;SPAN=1929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:83 GQ:43.7 PL:[43.7, 0.0, 155.9] SR:10 DR:11 LR:-43.53 LO:47.18);ALT=T[chr19:12762967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12763276	+	chr19	12766508	+	.	8	4	6735753_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6735753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12740001_12765001_82C;SPAN=3232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:4 DR:8 LR:-20.82 LO:23.18);ALT=T[chr19:12766508[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12788212	+	chr19	12790271	+	.	2	5	6735495_1	4.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6735495_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_12789001_12814001_10C;SPAN=2059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:44 GQ:4.7 PL:[4.7, 0.0, 100.4] SR:5 DR:2 LR:-4.584 LO:9.99);ALT=T[chr19:12790271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12791186	+	chr19	12792585	+	.	8	0	6735503_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6735503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12791186(+)-19:12792585(-)__19_12789001_12814001D;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:91 GQ:2 PL:[2.0, 0.0, 216.5] SR:0 DR:8 LR:-1.754 LO:15.04);ALT=G[chr19:12792585[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12841884	+	chr19	12845125	+	CATCCTCCGTCTTCTGCTTCTTGGCTACTATTCCCGTCTTGAGGGCTAGTTTGTTCCCGCCTCTGCGTTTGCCC	8	23	6735862_1	73.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=CATCCTCCGTCTTCTGCTTCTTGGCTACTATTCCCGTCTTGAGGGCTAGTTTGTTCCCGCCTCTGCGTTTGCCC;MAPQ=60;MATEID=6735862_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_12838001_12863001_109C;SPAN=3241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:84 GQ:73.1 PL:[73.1, 0.0, 129.2] SR:23 DR:8 LR:-72.97 LO:73.87);ALT=T[chr19:12845125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12842412	+	chr19	12845134	+	.	10	0	6735865_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6735865_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12842412(+)-19:12845134(-)__19_12838001_12863001D;SPAN=2722;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:101 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.647 LO:19.35);ALT=T[chr19:12845134[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12849473	+	chr19	12856190	+	.	0	8	6735889_1	5.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6735889_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_12838001_12863001_125C;SPAN=6717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:76 GQ:5.9 PL:[5.9, 0.0, 177.5] SR:8 DR:0 LR:-5.818 LO:15.7);ALT=G[chr19:12856190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	12885761	+	chr19	12889159	+	.	13	0	6736093_1	33.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6736093_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:12885761(+)-19:12889159(-)__19_12887001_12912001D;SPAN=3398;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:34 GQ:33.8 PL:[33.8, 0.0, 47.0] SR:0 DR:13 LR:-33.7 LO:33.85);ALT=G[chr19:12889159[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13041565	+	chr19	13044362	+	.	41	19	6736517_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=6736517_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_13034001_13059001_196C;SPAN=2797;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:95 GQ:99 PL:[129.5, 0.0, 99.8] SR:19 DR:41 LR:-129.6 LO:129.6);ALT=T[chr19:13044362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13051703	+	chr19	13054348	+	.	0	25	6736548_1	56.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=6736548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_13034001_13059001_78C;SPAN=2645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:97 GQ:56.3 PL:[56.3, 0.0, 178.4] SR:25 DR:0 LR:-56.25 LO:59.83);ALT=T[chr19:13054348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13056774	+	chr19	13058660	+	.	82	0	6736751_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6736751_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:13056774(+)-19:13058660(-)__19_13058501_13083501D;SPAN=1886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:38 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:0 DR:82 LR:-241.0 LO:241.0);ALT=C[chr19:13058660[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13056837	+	chr19	13058989	+	AAGGTGCTAAAGGAGAAGATAGAAGCTGAGAAGGGTCGTGATGCCTTCCCCGTGGCTGGACAGAAACTCATCTATGCCGGCAAGATCTTGAGTGACGATGTCCCTATCAGGGACTATCGCATCGATGAGAAGAACTTTGTGGTCGTCATGGTGACCA	0	72	6736753_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAGGTGCTAAAGGAGAAGATAGAAGCTGAGAAGGGTCGTGATGCCTTCCCCGTGGCTGGACAGAAACTCATCTATGCCGGCAAGATCTTGAGTGACGATGTCCCTATCAGGGACTATCGCATCGATGAGAAGAACTTTGTGGTCGTCATGGTGACCA;MAPQ=60;MATEID=6736753_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_13058501_13083501_171C;SPAN=2152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:72 DP:60 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:72 DR:0 LR:-211.3 LO:211.3);ALT=G[chr19:13058989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13065342	+	chr19	13067676	+	.	0	20	6736777_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6736777_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_13058501_13083501_9C;SPAN=2334;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:109 GQ:36.5 PL:[36.5, 0.0, 227.9] SR:20 DR:0 LR:-36.49 LO:44.49);ALT=T[chr19:13067676[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13212010	+	chr19	13213343	+	.	13	17	6737196_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6737196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_13205501_13230501_131C;SPAN=1333;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:89 GQ:55.1 PL:[55.1, 0.0, 160.7] SR:17 DR:13 LR:-55.11 LO:57.99);ALT=C[chr19:13213343[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13256211	+	chr19	13260312	+	CTCTGTTATTCCTCTCCAAAAATGCTACGGCTGTTGGGCTGACCATATGGTCCTTCATTT	4	12	6737348_1	21.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCTGGA;INSERTION=CTCTGTTATTCCTCTCCAAAAATGCTACGGCTGTTGGGCTGACCATATGGTCCTTCATTT;MAPQ=60;MATEID=6737348_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_13254501_13279501_282C;SPAN=4101;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:90 GQ:21.8 PL:[21.8, 0.0, 196.7] SR:12 DR:4 LR:-21.83 LO:30.03);ALT=T[chr19:13260312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13775699	+	chr19	13776846	+	.	14	0	6738953_1	29.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6738953_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:13775699(+)-19:13776846(-)__19_13769001_13794001D;SPAN=1147;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:62 GQ:29.6 PL:[29.6, 0.0, 118.7] SR:0 DR:14 LR:-29.42 LO:32.57);ALT=A[chr19:13776846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13858810	+	chr19	13862463	+	.	8	0	6739650_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6739650_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:13858810(+)-19:13862463(-)__19_13842501_13867501D;SPAN=3653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=C[chr19:13862463[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13885390	+	chr19	13888864	+	CGTGTTATCGCTCCCAGGAAGGCGCGCGTCGTGCAGCAGCAAAAGCTCAAGA	0	76	6739545_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CGTGTTATCGCTCCCAGGAAGGCGCGCGTCGTGCAGCAGCAAAAGCTCAAGA;MAPQ=60;MATEID=6739545_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_13867001_13892001_36C;SPAN=3474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:76 DP:109 GQ:43.1 PL:[221.3, 0.0, 43.1] SR:76 DR:0 LR:-228.1 LO:228.1);ALT=T[chr19:13888864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	13885521	+	chr19	13888864	+	.	105	63	6739548_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6739548_2;MATENM=0;NM=1;NUMPARTS=3;REPSEQ=GAAGAA;SCTG=c_19_13867001_13892001_36C;SPAN=3343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:140 DP:121 GQ:37.7 PL:[327.7, 37.7, 0.0] SR:63 DR:105 LR:-327.7 LO:327.7);ALT=G[chr19:13888864[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14063404	+	chr19	14065149	+	.	8	0	6740421_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6740421_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14063404(+)-19:14065149(-)__19_14038501_14063501D;SPAN=1745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=G[chr19:14065149[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14248069	+	chr19	14265964	+	.	15	0	6741052_1	39.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6741052_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14248069(+)-19:14265964(-)__19_14234501_14259501D;SPAN=17895;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:38 GQ:39.2 PL:[39.2, 0.0, 52.4] SR:0 DR:15 LR:-39.22 LO:39.33);ALT=C[chr19:14265964[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14266291	+	chr19	14281934	+	.	0	8	6740927_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=6740927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14259001_14284001_221C;SPAN=15643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:8 DR:0 LR:-3.109 LO:15.25);ALT=G[chr19:14281934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14492357	+	chr19	14499261	+	.	65	33	6742295_1	99.0	.	DISC_MAPQ=41;EVDNC=ASDIS;HOMSEQ=G;MAPQ=58;MATEID=6742295_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_19_14479501_14504501_10C;SPAN=6904;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:106 GQ:21.9 PL:[300.3, 21.9, 0.0] SR:33 DR:65 LR:-302.1 LO:302.1);ALT=G[chr19:14499261[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14499260	-	chr19	14887590	+	.	47	0	6742323_1	99.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6742323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14499260(-)-19:14887590(-)__19_14479501_14504501D;SPAN=388330;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:55 GQ:8.1 PL:[148.5, 8.1, 0.0] SR:0 DR:47 LR:-150.8 LO:150.8);ALT=[chr19:14887590[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	14499630	+	chr19	14501735	+	.	0	31	6742330_1	72.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=45;MATEID=6742330_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14479501_14504501_32C;SPAN=2105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:110 GQ:72.5 PL:[72.5, 0.0, 194.6] SR:31 DR:0 LR:-72.53 LO:75.61);ALT=G[chr19:14501735[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14501734	-	chr19	14887593	+	.	11	0	6742345_1	21.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6742345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14501734(-)-19:14887593(-)__19_14479501_14504501D;SPAN=385859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=[chr19:14887593[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	14523525	+	chr19	14530081	+	.	10	0	6742375_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6742375_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14523525(+)-19:14530081(-)__19_14528501_14553501D;SPAN=6556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:64 GQ:15.8 PL:[15.8, 0.0, 137.9] SR:0 DR:10 LR:-15.67 LO:21.47);ALT=T[chr19:14530081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14524083	+	chr19	14530081	+	.	37	0	6742376_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6742376_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14524083(+)-19:14530081(-)__19_14528501_14553501D;SPAN=5998;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:64 GQ:48.8 PL:[104.9, 0.0, 48.8] SR:0 DR:37 LR:-105.8 LO:105.8);ALT=G[chr19:14530081[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14627860	+	chr19	14628950	+	.	0	174	6742657_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6742657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14626501_14651501_12C;SPAN=1090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:174 DP:156 GQ:46.9 PL:[514.9, 46.9, 0.0] SR:174 DR:0 LR:-514.9 LO:514.9);ALT=T[chr19:14628950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14640506	+	chr19	14674611	+	.	10	0	6742700_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6742700_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14640506(+)-19:14674611(-)__19_14626501_14651501D;SPAN=34105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:50 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.46 LO:22.66);ALT=G[chr19:14674611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14640525	+	chr19	14673984	+	GGAGATTCTGGACGCAAAGACAAGGGAGAAGCTGTGTTTCTTGGACA	6	10	6742582_1	35.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=GGAGATTCTGGACGCAAAGACAAGGGAGAAGCTGTGTTTCTTGGACA;MAPQ=60;MATEID=6742582_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_14651001_14676001_334C;SPAN=33459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:42 GQ:35 PL:[35.0, 0.0, 64.7] SR:10 DR:6 LR:-34.84 LO:35.4);ALT=T[chr19:14673984[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14640525	+	chr19	14673333	+	.	5	10	6742701_1	34.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=ACCTCG;MAPQ=60;MATEID=6742701_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_19_14626501_14651501_27C;SPAN=32808;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:43 GQ:34.7 PL:[34.7, 0.0, 67.7] SR:10 DR:5 LR:-34.56 LO:35.22);ALT=T[chr19:14673333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14677746	+	chr19	14682701	+	.	0	80	6742782_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6742782_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_14675501_14700501_96C;SPAN=4955;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:80 DP:129 GQ:83.9 PL:[229.1, 0.0, 83.9] SR:80 DR:0 LR:-232.8 LO:232.8);ALT=C[chr19:14682701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14732345	+	chr19	14734127	+	.	63	36	6743190_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=TAAAACTCCTGGACTT;MAPQ=60;MATEID=6743190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_14724501_14749501_298C;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:87 DP:127 GQ:54.8 PL:[252.8, 0.0, 54.8] SR:36 DR:63 LR:-259.9 LO:259.9);ALT=T[chr19:14734127[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	14884916	+	chr19	14887592	+	.	13	0	6743487_1	17.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6743487_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:14884916(+)-19:14887592(-)__19_14871501_14896501D;SPAN=2676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:93 GQ:17.9 PL:[17.9, 0.0, 206.0] SR:0 DR:13 LR:-17.72 LO:27.23);ALT=A[chr19:14887592[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15046392	+	chr19	15049478	+	.	15	14	6744070_1	70.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=T;MAPQ=60;MATEID=6744070_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_15043001_15068001_117C;SPAN=3086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:46 GQ:40.4 PL:[70.1, 0.0, 40.4] SR:14 DR:15 LR:-70.45 LO:70.45);ALT=T[chr19:15049478[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15330770	-	chr19	15332033	+	.	10	0	6745218_1	7.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6745218_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:15330770(-)-19:15332033(-)__19_15312501_15337501D;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:94 GQ:7.7 PL:[7.7, 0.0, 218.9] SR:0 DR:10 LR:-7.543 LO:19.68);ALT=[chr19:15332033[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	15367988	+	chr19	15374230	+	.	4	14	6744762_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTGG;MAPQ=60;MATEID=6744762_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_15361501_15386501_155C;SPAN=6242;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:76 GQ:38.9 PL:[38.9, 0.0, 144.5] SR:14 DR:4 LR:-38.83 LO:42.31);ALT=G[chr19:15374230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15367988	+	chr19	15375215	+	AGCTTGCGGGCCATGGCCACCACCTCATGGTCAGGAGGGTTGTACTTATAGCAGTTGGAGAACATCAATCGGACGTCAGCACCAAACTCCTGAGCATCACGGTACTCACGGGCCTCCAGTTTAGA	5	19	6744763_1	49.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=AGCTTGCGGGCCATGGCCACCACCTCATGGTCAGGAGGGTTGTACTTATAGCAGTTGGAGAACATCAATCGGACGTCAGCACCAAACTCCTGAGCATCACGGTACTCACGGGCCTCCAGTTTAGA;MAPQ=60;MATEID=6744763_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_15361501_15386501_155C;SPAN=7227;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:73 GQ:49.7 PL:[49.7, 0.0, 125.6] SR:19 DR:5 LR:-49.54 LO:51.45);ALT=G[chr19:15375215[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15376456	+	chr19	15378226	+	.	16	5	6744793_1	33.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6744793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_15361501_15386501_9C;SPAN=1770;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:83 GQ:33.8 PL:[33.8, 0.0, 165.8] SR:5 DR:16 LR:-33.63 LO:38.73);ALT=T[chr19:15378226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15484869	+	chr19	15490522	+	.	8	0	6745714_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6745714_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:15484869(+)-19:15490522(-)__19_15484001_15509001D;SPAN=5653;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:80 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:0 DR:8 LR:-4.734 LO:15.51);ALT=T[chr19:15490522[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15514528	+	chr19	15521330	+	CTATTTGTCCCAGAGTTCCAAGTTCCATAT	0	9	6745431_1	3.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CTATTTGTCCCAGAGTTCCAAGTTCCATAT;MAPQ=60;MATEID=6745431_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_15508501_15533501_158C;SPAN=6802;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:98 GQ:3.2 PL:[3.2, 0.0, 234.2] SR:9 DR:0 LR:-3.158 LO:17.1);ALT=T[chr19:15521330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	15514587	+	chr19	15529720	+	.	10	0	6745432_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6745432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:15514587(+)-19:15529720(-)__19_15508501_15533501D;SPAN=15133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:0 DR:10 LR:-8.898 LO:19.93);ALT=A[chr19:15529720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16187508	+	chr19	16192723	+	.	0	67	6747796_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6747796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16170001_16195001_100C;SPAN=5215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:72 GQ:19.2 PL:[211.2, 19.2, 0.0] SR:67 DR:0 LR:-211.3 LO:211.3);ALT=G[chr19:16192723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16222810	+	chr19	16232557	+	.	28	0	6747566_1	70.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6747566_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16222810(+)-19:16232557(-)__19_16219001_16244001D;SPAN=9747;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:81 GQ:70.7 PL:[70.7, 0.0, 123.5] SR:0 DR:28 LR:-70.48 LO:71.35);ALT=C[chr19:16232557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16222836	+	chr19	16229034	+	.	24	23	6747567_1	74.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6747567_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=GG;SCTG=c_19_16219001_16244001_376C;SPAN=6198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:81 GQ:74 PL:[74.0, 0.0, 120.2] SR:23 DR:24 LR:-73.78 LO:74.45);ALT=G[chr19:16229034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16222836	+	chr19	16236279	+	AATTGACTTTAAAATTAGGACCATAGAGCTCGATGGCAAGAGAATTAAACTGCAGATATGGGACACAGCCGGTCAGGAACGGTTTCGGACGATCACAACGGCCTACTACAGGGGTGCAAT	11	55	6747568_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=GG;INSERTION=AATTGACTTTAAAATTAGGACCATAGAGCTCGATGGCAAGAGAATTAAACTGCAGATATGGGACACAGCCGGTCAGGAACGGTTTCGGACGATCACAACGGCCTACTACAGGGGTGCAAT;MAPQ=60;MATEID=6747568_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_16219001_16244001_376C;SPAN=13443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:94 GQ:57.2 PL:[169.4, 0.0, 57.2] SR:55 DR:11 LR:-172.2 LO:172.2);ALT=G[chr19:16236279[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16254586	+	chr19	16259529	+	.	66	14	6747887_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCCAGGT;MAPQ=60;MATEID=6747887_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16243501_16268501_339C;SPAN=4943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:136 GQ:99 PL:[200.9, 0.0, 128.3] SR:14 DR:66 LR:-201.7 LO:201.7);ALT=T[chr19:16259529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16254627	+	chr19	16263361	+	.	67	0	6747889_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6747889_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16254627(+)-19:16263361(-)__19_16243501_16268501D;SPAN=8734;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:118 GQ:96.8 PL:[189.2, 0.0, 96.8] SR:0 DR:67 LR:-190.8 LO:190.8);ALT=G[chr19:16263361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16259686	+	chr19	16263362	+	.	7	86	6747914_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6747914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16243501_16268501_358C;SPAN=3676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:92 DP:152 GQ:99 PL:[262.7, 0.0, 104.3] SR:86 DR:7 LR:-266.1 LO:266.1);ALT=G[chr19:16263362[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16264018	+	chr19	16265257	+	.	0	16	6747940_1	15.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=6747940_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16243501_16268501_346C;SPAN=1239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:139 GQ:15.2 PL:[15.2, 0.0, 322.1] SR:16 DR:0 LR:-15.16 LO:32.06);ALT=G[chr19:16265257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16265302	+	chr19	16268018	+	.	4	5	6748091_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6748091_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16268001_16293001_370C;SPAN=2716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:42 GQ:15.2 PL:[15.2, 0.0, 84.5] SR:5 DR:4 LR:-15.03 LO:17.94);ALT=G[chr19:16268018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16308881	+	chr19	16314268	+	.	37	20	6748229_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6748229_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16292501_16317501_235C;SPAN=5387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:84 GQ:69.8 PL:[132.5, 0.0, 69.8] SR:20 DR:37 LR:-133.4 LO:133.4);ALT=T[chr19:16314268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16435814	+	chr19	16437665	+	.	31	19	6748677_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGGTGAG;MAPQ=60;MATEID=6748677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16415001_16440001_342C;SPAN=1851;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:108 GQ:99 PL:[129.2, 0.0, 132.5] SR:19 DR:31 LR:-129.2 LO:129.2);ALT=G[chr19:16437665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16758122	+	chr19	16770894	+	.	22	0	6749765_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6749765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16758122(+)-19:16770894(-)__19_16758001_16783001D;SPAN=12772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:99 GQ:45.8 PL:[45.8, 0.0, 194.3] SR:0 DR:22 LR:-45.8 LO:51.0);ALT=T[chr19:16770894[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16764981	+	chr19	16770893	+	.	20	0	6749783_1	41.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6749783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16764981(+)-19:16770893(-)__19_16758001_16783001D;SPAN=5912;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:93 GQ:41 PL:[41.0, 0.0, 182.9] SR:0 DR:20 LR:-40.82 LO:46.04);ALT=T[chr19:16770893[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	16865939	+	chr19	16864680	+	.	25	0	6749868_1	61.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6749868_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:16864680(-)-19:16865939(+)__19_16856001_16881001D;SPAN=1259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:77 GQ:61.7 PL:[61.7, 0.0, 124.4] SR:0 DR:25 LR:-61.66 LO:62.85);ALT=]chr19:16865939]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	16940708	+	chr19	16942303	+	.	0	7	6750491_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6750491_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_16929501_16954501_273C;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:66 GQ:5.3 PL:[5.3, 0.0, 153.8] SR:7 DR:0 LR:-5.226 LO:13.76);ALT=G[chr19:16942303[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17186684	+	chr19	17212468	+	.	12	2	6751301_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6751301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_17199001_17224001_259C;SPAN=25784;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:2 DR:12 LR:-27.96 LO:29.21);ALT=G[chr19:17212468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17378336	+	chr19	17379601	+	.	84	3	6752067_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6752067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_17370501_17395501_112C;SPAN=1265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:84 DP:81 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:3 DR:84 LR:-247.6 LO:247.6);ALT=G[chr19:17379601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17387719	+	chr19	17389652	+	.	7	9	6752103_1	30.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6752103_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_17370501_17395501_241C;SPAN=1933;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:69 GQ:30.8 PL:[30.8, 0.0, 136.4] SR:9 DR:7 LR:-30.82 LO:34.61);ALT=G[chr19:17389652[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17403663	+	chr19	17407523	+	.	0	7	6752192_1	2.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6752192_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_17395001_17420001_239C;SPAN=3860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:7 DR:0 LR:-2.246 LO:13.27);ALT=G[chr19:17407523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18800243	+	chr19	17424254	+	.	8	0	6757385_1	20.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=6757385_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:17424254(-)-19:18800243(+)__19_18791501_18816501D;SPAN=1375989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:22 GQ:20.6 PL:[20.6, 0.0, 30.5] SR:0 DR:8 LR:-20.45 LO:20.61);ALT=]chr19:18800243]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	17514635	+	chr19	17516100	+	CAGTCGCTCCACCTCTGCAGACGCGTCCTGAAGCTTATGGTTTAATGTAGTGATCTCTCCCTCAAGCTCCTCCACTTTCTTTTGTCCTTGGGCCTTCTCTGCATCCAGGGAAGCCATTAGGGCCAT	0	32	6752608_1	80.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CAGTCGCTCCACCTCTGCAGACGCGTCCTGAAGCTTATGGTTTAATGTAGTGATCTCTCCCTCAAGCTCCTCCACTTTCTTTTGTCCTTGGGCCTTCTCTGCATCCAGGGAAGCCATTAGGGCCAT;MAPQ=60;MATEID=6752608_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_17493001_17518001_54C;SPAN=1465;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:93 GQ:80.6 PL:[80.6, 0.0, 143.3] SR:32 DR:0 LR:-80.44 LO:81.46);ALT=T[chr19:17516100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17622769	+	chr19	17628094	+	ACGCATCTTCTCTCCAGACTGCCGATCCCAGAAAGCCAGGTGATCACCATTAACCCCGAGCTGCCTGTGGAGGAGGCGGCTGAGGACTACGCCAAGAAGCTGAGA	2	83	6752912_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=ACGCATCTTCTCTCCAGACTGCCGATCCCAGAAAGCCAGGTGATCACCATTAACCCCGAGCTGCCTGTGGAGGAGGCGGCTGAGGACTACGCCAAGAAGCTGAGA;MAPQ=60;MATEID=6752912_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_17615501_17640501_48C;SPAN=5325;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:84 DP:108 GQ:13.7 PL:[248.0, 0.0, 13.7] SR:83 DR:2 LR:-260.5 LO:260.5);ALT=G[chr19:17628094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17622769	+	chr19	17626981	+	.	17	70	6752911_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6752911_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_17615501_17640501_48C;SPAN=4212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:86 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:70 DR:17 LR:-254.2 LO:254.2);ALT=G[chr19:17626981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17627090	+	chr19	17628094	+	.	3	12	6752923_1	20.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAGG;MAPQ=60;MATEID=6752923_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_17615501_17640501_48C;SPAN=1004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:97 GQ:20 PL:[20.0, 0.0, 214.7] SR:12 DR:3 LR:-19.93 LO:29.53);ALT=G[chr19:17628094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	17628659	+	chr19	17631751	+	.	11	17	6752935_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6752935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_17615501_17640501_271C;SPAN=3092;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:108 GQ:53.3 PL:[53.3, 0.0, 208.4] SR:17 DR:11 LR:-53.27 LO:58.47);ALT=G[chr19:17631751[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18043907	+	chr19	18047229	+	.	8	0	6754373_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6754373_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18043907(+)-19:18047229(-)__19_18032001_18057001D;SPAN=3322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:121 GQ:6 PL:[0.0, 6.0, 303.6] SR:0 DR:8 LR:6.374 LO:14.01);ALT=G[chr19:18047229[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18043908	+	chr19	18053462	+	.	40	0	6754374_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6754374_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18043908(+)-19:18053462(-)__19_18032001_18057001D;SPAN=9554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:82 GQ:86.9 PL:[110.0, 0.0, 86.9] SR:0 DR:40 LR:-109.9 LO:109.9);ALT=C[chr19:18053462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18047389	+	chr19	18053463	+	.	30	56	6754392_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6754392_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_18032001_18057001_180C;SPAN=6074;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:71 DP:112 GQ:65.6 PL:[204.2, 0.0, 65.6] SR:56 DR:30 LR:-207.8 LO:207.8);ALT=G[chr19:18053463[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18284783	+	chr19	18285848	+	.	82	66	6755349_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6755349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18277001_18302001_56C;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:118 DP:152 GQ:18.5 PL:[348.5, 0.0, 18.5] SR:66 DR:82 LR:-365.7 LO:365.7);ALT=G[chr19:18285848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18286507	+	chr19	18287950	+	.	7	7	6755357_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6755357_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18277001_18302001_112C;SPAN=1443;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:7 DR:7 LR:-9.982 LO:20.14);ALT=A[chr19:18287950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18418367	+	chr19	18420485	+	.	10	10	6755746_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=6755746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18399501_18424501_334C;SPAN=2118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:82 GQ:34.1 PL:[34.1, 0.0, 162.8] SR:10 DR:10 LR:-33.9 LO:38.83);ALT=T[chr19:18420485[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18420672	+	chr19	18423413	+	.	4	112	6755753_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6755753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18399501_18424501_50C;SPAN=2741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:140 GQ:1.5 PL:[343.2, 1.5, 0.0] SR:112 DR:4 LR:-363.4 LO:363.4);ALT=C[chr19:18423413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18420721	+	chr19	18433825	+	.	79	0	6755900_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6755900_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18420721(+)-19:18433825(-)__19_18424001_18449001D;SPAN=13104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:49 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:0 DR:79 LR:-234.4 LO:234.4);ALT=C[chr19:18433825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18423513	+	chr19	18426834	+	.	3	39	6755767_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6755767_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_18399501_18424501_202C;SPAN=3321;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:53 GQ:2.3 PL:[124.4, 0.0, 2.3] SR:39 DR:3 LR:-131.1 LO:131.1);ALT=C[chr19:18426834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18423569	+	chr19	18433825	+	.	93	0	6755769_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6755769_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18423569(+)-19:18433825(-)__19_18399501_18424501D;SPAN=10256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:31 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:93 LR:-274.0 LO:274.0);ALT=C[chr19:18433825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18426933	+	chr19	18433827	+	.	10	0	6755914_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6755914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18426933(+)-19:18433827(-)__19_18424001_18449001D;SPAN=6894;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:100 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.918 LO:19.39);ALT=G[chr19:18433827[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18451533	+	chr19	18466701	+	.	9	0	6756124_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6756124_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18451533(+)-19:18466701(-)__19_18448501_18473501D;SPAN=15168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-8.035 LO:17.94);ALT=G[chr19:18466701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18466821	+	chr19	18468190	+	.	0	6	6756193_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6756193_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18448501_18473501_63C;SPAN=1369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:83 GQ:2.4 PL:[0.0, 2.4, 204.6] SR:6 DR:0 LR:2.681 LO:10.75);ALT=G[chr19:18468190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18650531	+	chr19	18652488	+	.	0	11	6756962_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6756962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18644501_18669501_132C;SPAN=1957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:93 GQ:11.3 PL:[11.3, 0.0, 212.6] SR:11 DR:0 LR:-11.12 LO:22.18);ALT=C[chr19:18652488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18652807	+	chr19	18654295	+	.	137	12	6756974_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6756974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18644501_18669501_231C;SPAN=1488;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:143 DP:97 GQ:38.5 PL:[422.5, 38.5, 0.0] SR:12 DR:137 LR:-422.5 LO:422.5);ALT=T[chr19:18654295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18668725	+	chr19	18672843	+	.	20	5	6757073_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6757073_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18669001_18694001_54C;SPAN=4118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:40 GQ:32 PL:[65.0, 0.0, 32.0] SR:5 DR:20 LR:-65.7 LO:65.7);ALT=G[chr19:18672843[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18668772	+	chr19	18675678	+	.	53	0	6757075_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6757075_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18668772(+)-19:18675678(-)__19_18669001_18694001D;SPAN=6906;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:55 GQ:14.7 PL:[161.7, 14.7, 0.0] SR:0 DR:53 LR:-161.7 LO:161.7);ALT=A[chr19:18675678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18672968	+	chr19	18675679	+	.	3	44	6757093_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6757093_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18669001_18694001_223C;SPAN=2711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:102 GQ:99 PL:[124.4, 0.0, 121.1] SR:44 DR:3 LR:-124.2 LO:124.2);ALT=G[chr19:18675679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18675832	+	chr19	18679212	+	ACGCTGAAAGGGAAACTGGCCAGGCAGCACCCAGAGGCCTTCAGCC	2	16	6757101_1	26.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=ACGCTGAAAGGGAAACTGGCCAGGCAGCACCCAGAGGCCTTCAGCC;MAPQ=60;MATEID=6757101_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_18669001_18694001_284C;SPAN=3380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:96 GQ:26.9 PL:[26.9, 0.0, 205.1] SR:16 DR:2 LR:-26.81 LO:34.85);ALT=G[chr19:18679212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18682754	+	chr19	18684094	+	.	26	0	6757133_1	50.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6757133_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18682754(+)-19:18684094(-)__19_18669001_18694001D;SPAN=1340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:133 GQ:50 PL:[50.0, 0.0, 271.1] SR:0 DR:26 LR:-49.79 LO:58.63);ALT=G[chr19:18684094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18682766	+	chr19	18685677	+	.	35	0	6757135_1	55.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6757135_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:18682766(+)-19:18685677(-)__19_18669001_18694001D;SPAN=2911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:220 GQ:55.9 PL:[55.9, 0.0, 478.4] SR:0 DR:35 LR:-55.93 LO:75.45);ALT=G[chr19:18685677[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18684558	+	chr19	18685678	+	.	24	85	6757139_1	99.0	.	DISC_MAPQ=29;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6757139_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18669001_18694001_351C;SPAN=1120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:328 GQ:99 PL:[261.1, 0.0, 535.1] SR:85 DR:24 LR:-261.0 LO:266.2);ALT=G[chr19:18685678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18700496	+	chr19	18701663	+	.	6	24	6757301_1	65.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6757301_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18693501_18718501_98C;SPAN=1167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:89 GQ:65 PL:[65.0, 0.0, 150.8] SR:24 DR:6 LR:-65.02 LO:66.9);ALT=G[chr19:18701663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	18701744	+	chr19	18702918	+	.	4	57	6757305_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6757305_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_18693501_18718501_230C;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:118 GQ:99 PL:[162.8, 0.0, 123.2] SR:57 DR:4 LR:-163.1 LO:163.1);ALT=G[chr19:18702918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19010538	+	chr19	19014076	+	GGCCTGGTACTCCTTGATGAAGGGATGGGACCTGTGGGCATCCTTCAGCTGGGACAGGTATCGGTTTGTCACCTCAGGGGGCTTGCCCAGGTGCTGGGACAGGACGATGAGGTTGACCAGCGTCTCTGGGTAGCCACTAT	0	137	6758066_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=GGCCTGGTACTCCTTGATGAAGGGATGGGACCTGTGGGCATCCTTCAGCTGGGACAGGTATCGGTTTGTCACCTCAGGGGGCTTGCCCAGGTGCTGGGACAGGACGATGAGGTTGACCAGCGTCTCTGGGTAGCCACTAT;MAPQ=60;MATEID=6758066_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_18987501_19012501_151C;SPAN=3538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:137 DP:59 GQ:36.9 PL:[405.9, 36.9, 0.0] SR:137 DR:0 LR:-406.0 LO:406.0);ALT=T[chr19:19014076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19011260	+	chr19	19014076	+	.	3	16	6758069_1	45.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=6758069_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_18987501_19012501_151C;SPAN=2816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:51 GQ:45.8 PL:[45.8, 0.0, 75.5] SR:16 DR:3 LR:-45.6 LO:46.07);ALT=T[chr19:19014076[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19017923	+	chr19	19021779	+	.	5	45	6758101_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6758101_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_19012001_19037001_289C;SPAN=3856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:49 DP:104 GQ:99 PL:[133.7, 0.0, 117.2] SR:45 DR:5 LR:-133.6 LO:133.6);ALT=T[chr19:19021779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19017972	+	chr19	19030105	+	.	28	0	6758103_1	68.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6758103_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19017972(+)-19:19030105(-)__19_19012001_19037001D;SPAN=12133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:89 GQ:68.3 PL:[68.3, 0.0, 147.5] SR:0 DR:28 LR:-68.32 LO:69.92);ALT=C[chr19:19030105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19021941	+	chr19	19030031	+	.	90	0	6758114_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6758114_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19021941(+)-19:19030031(-)__19_19012001_19037001D;SPAN=8090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:90 DP:93 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:0 DR:90 LR:-274.0 LO:274.0);ALT=G[chr19:19030031[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19023906	+	chr19	19030103	+	.	81	0	6758130_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6758130_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19023906(+)-19:19030103(-)__19_19012001_19037001D;SPAN=6197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:85 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:0 DR:81 LR:-250.9 LO:250.9);ALT=C[chr19:19030103[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19040400	+	chr19	19042131	+	.	10	0	6758309_1	5.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6758309_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19040400(+)-19:19042131(-)__19_19036501_19061501D;SPAN=1731;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:104 GQ:5 PL:[5.0, 0.0, 245.9] SR:0 DR:10 LR:-4.834 LO:19.21);ALT=G[chr19:19042131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19049859	+	chr19	19051859	+	.	34	8	6758350_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6758350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_19036501_19061501_239C;SPAN=2000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:61 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:8 DR:34 LR:-107.1 LO:107.1);ALT=C[chr19:19051859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19144806	+	chr19	19153516	+	.	8	0	6758510_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6758510_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19144806(+)-19:19153516(-)__19_19134501_19159501D;SPAN=8710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:81 GQ:4.7 PL:[4.7, 0.0, 189.5] SR:0 DR:8 LR:-4.463 LO:15.47);ALT=G[chr19:19153516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19309041	+	chr19	19312456	+	AATGGAGGGACGCCACTGCTGTACGCTGTGCGCGGGAACCACGTGAAATGCGTTGAGGCCTTGCTGGCCCGAGGCGCTGACCTCACCACCGAAGCCGACTCTGGCTACACCCCGATGGACCTTGCCGTGGCCCTGGGATACCGGAA	0	44	6759521_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AATGGAGGGACGCCACTGCTGTACGCTGTGCGCGGGAACCACGTGAAATGCGTTGAGGCCTTGCTGGCCCGAGGCGCTGACCTCACCACCGAAGCCGACTCTGGCTACACCCCGATGGACCTTGCCGTGGCCCTGGGATACCGGAA;MAPQ=60;MATEID=6759521_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_19306001_19331001_79C;SPAN=3415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:91 GQ:97.7 PL:[120.8, 0.0, 97.7] SR:44 DR:0 LR:-120.7 LO:120.7);ALT=G[chr19:19312456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19627142	+	chr19	19638087	+	CTACAGCATGCTGGCCATAGGGATTGGAACCCTGATCTACGGGCACTGGAGCATAATGAAGTGGAACCGTGAGCG	0	188	6760415_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CTACAGCATGCTGGCCATAGGGATTGGAACCCTGATCTACGGGCACTGGAGCATAATGAAGTGGAACCGTGAGCG;MAPQ=60;MATEID=6760415_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_19624501_19649501_44C;SPAN=10945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:188 DP:182 GQ:50.8 PL:[557.8, 50.8, 0.0] SR:188 DR:0 LR:-557.8 LO:557.8);ALT=G[chr19:19638087[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19627142	+	chr19	19636990	+	.	87	42	6760414_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6760414_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_19_19624501_19649501_44C;SPAN=9848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:173 DP:102 GQ:46.6 PL:[511.6, 46.6, 0.0] SR:42 DR:87 LR:-511.6 LO:511.6);ALT=G[chr19:19636990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	19627192	+	chr19	19638507	+	.	29	0	6760416_1	51.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6760416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:19627192(+)-19:19638507(-)__19_19624501_19649501D;SPAN=11315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:165 GQ:51.2 PL:[51.2, 0.0, 348.2] SR:0 DR:29 LR:-51.03 LO:63.9);ALT=G[chr19:19638507[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	20801300	+	chr19	20883926	-	.	11	0	6763923_1	21.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=6763923_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:20801300(+)-19:20883926(+)__19_20874001_20899001D;SPAN=82626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=A]chr19:20883926];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	21106210	+	chr19	21116829	+	.	10	3	6764531_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=13;MATEID=6764531_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_21094501_21119501_372C;SPAN=10619;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:77 GQ:15.5 PL:[15.5, 0.0, 170.6] SR:3 DR:10 LR:-15.45 LO:23.15);ALT=G[chr19:21116829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21203610	+	chr19	21205594	+	.	0	7	6764817_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6764817_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_21192501_21217501_317C;SPAN=1984;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:7 DR:0 LR:-0.6203 LO:13.03);ALT=G[chr19:21205594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21324990	+	chr19	21326353	+	.	13	6	6765243_1	26.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6765243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_21315001_21340001_219C;SPAN=1363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:85 GQ:26.6 PL:[26.6, 0.0, 178.4] SR:6 DR:13 LR:-26.49 LO:33.08);ALT=G[chr19:21326353[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21492144	+	chr19	21512010	+	.	2	3	6765799_1	7.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6765799_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_21486501_21511501_174C;SPAN=19866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:34 GQ:7.4 PL:[7.4, 0.0, 73.4] SR:3 DR:2 LR:-7.294 LO:10.59);ALT=C[chr19:21512010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21541946	+	chr19	21544567	+	.	8	4	6765705_1	11.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6765705_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_21535501_21560501_221C;SPAN=2621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:81 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:4 DR:8 LR:-11.07 LO:20.36);ALT=G[chr19:21544567[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	21903056	+	chr19	21905568	+	.	22	11	6767557_1	89.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TGTTAT;MAPQ=60;MATEID=6767557_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_21878501_21903501_310C;SPAN=2512;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:31 DP:11 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:11 DR:22 LR:-89.12 LO:89.12);ALT=T[chr19:21905568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	22989471	+	chr19	22444405	+	GGAGGGACAAGCGGGCGGAGAAGGGGCGGCCCT	0	17	6770380_1	46.0	.	EVDNC=ASSMB;INSERTION=GGAGGGACAAGCGGGCGGAGAAGGGGCGGCCCT;MAPQ=60;MATEID=6770380_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_22981001_23006001_290C;SPAN=545066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:35 GQ:36.8 PL:[46.7, 0.0, 36.8] SR:17 DR:0 LR:-46.68 LO:46.68);ALT=]chr19:22989471]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	22444698	+	chr19	22989451	-	.	13	0	6770382_1	32.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6770382_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:22444698(+)-19:22989451(+)__19_22981001_23006001D;SPAN=544753;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:38 GQ:32.6 PL:[32.6, 0.0, 59.0] SR:0 DR:13 LR:-32.62 LO:33.05);ALT=G]chr19:22989451];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	22444851	-	chr19	22989327	+	.	10	0	6770383_1	21.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6770383_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:22444851(-)-19:22989327(-)__19_22981001_23006001D;SPAN=544476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:43 GQ:21.5 PL:[21.5, 0.0, 80.9] SR:0 DR:10 LR:-21.36 LO:23.41);ALT=[chr19:22989327[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	23140838	+	chr19	23142919	+	.	14	0	6770778_1	34.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6770778_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:23140838(+)-19:23142919(-)__19_23128001_23153001D;SPAN=2081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:43 GQ:34.7 PL:[34.7, 0.0, 67.7] SR:0 DR:14 LR:-34.56 LO:35.22);ALT=A[chr19:23142919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	23805793	+	chr19	23808308	+	.	23	28	6772745_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=GGGTTCAAGCAATTCTCCTGCCTCAGCCTCCC;MAPQ=60;MATEID=6772745_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_19_23789501_23814501_162C;SPAN=2515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:48 DP:26 GQ:12.9 PL:[141.9, 12.9, 0.0] SR:28 DR:23 LR:-141.9 LO:141.9);ALT=C[chr19:23808308[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24270079	+	chr19	24289348	+	.	8	0	6774524_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6774524_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:24270079(+)-19:24289348(-)__19_24279501_24304501D;SPAN=19269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:35 GQ:17 PL:[17.0, 0.0, 66.5] SR:0 DR:8 LR:-16.93 LO:18.66);ALT=T[chr19:24289348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24270140	+	chr19	24288741	+	.	8	3	6774525_1	26.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6774525_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_19_24279501_24304501_152C;SECONDARY;SPAN=18601;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:38 GQ:26 PL:[26.0, 0.0, 65.6] SR:3 DR:8 LR:-26.02 LO:26.98);ALT=G[chr19:24288741[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24459052	+	chr19	24464776	+	GA	25	22	6774958_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;INSERTION=GA;MAPQ=60;MATEID=6774958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_24451001_24476001_96C;SPAN=5724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:50 GQ:12.8 PL:[108.5, 0.0, 12.8] SR:22 DR:25 LR:-113.0 LO:113.0);ALT=T[chr19:24464776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	24595035	+	chr19	24596046	+	.	38	23	6775996_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=CTCTTTTTGTAGAATCT;MAPQ=60;MATEID=6775996_2;MATENM=3;NM=1;NUMPARTS=2;SCTG=c_19_24573501_24598501_452C;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:72 GQ:13.7 PL:[158.9, 0.0, 13.7] SR:23 DR:38 LR:-165.6 LO:165.6);ALT=T[chr19:24596046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	29699068	+	chr19	29703968	+	.	17	0	6781391_1	32.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=6781391_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:29699068(+)-19:29703968(-)__19_29694001_29719001D;SPAN=4900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:89 GQ:32 PL:[32.0, 0.0, 183.8] SR:0 DR:17 LR:-32.01 LO:38.15);ALT=G[chr19:29703968[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	29950197	+	chr19	29956168	+	.	0	33	6782174_1	95.0	.	EVDNC=ASSMB;HOMSEQ=AAAAAAGAAATTA;MAPQ=60;MATEID=6782174_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_29939001_29964001_164C;SPAN=5971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:33 DP:29 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:33 DR:0 LR:-95.72 LO:95.72);ALT=A[chr19:29956168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	30099656	+	chr19	30101312	+	.	12	0	6782290_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6782290_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:30099656(+)-19:30101312(-)__19_30086001_30111001D;SPAN=1656;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:87 GQ:16.1 PL:[16.1, 0.0, 194.3] SR:0 DR:12 LR:-16.04 LO:25.06);ALT=T[chr19:30101312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	30388804	+	chr19	30393101	+	.	80	41	6783648_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=TAATTTTTATTTTT;MAPQ=60;MATEID=6783648_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_30380001_30405001_173C;SPAN=4297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:94 DP:78 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:41 DR:80 LR:-277.3 LO:277.3);ALT=T[chr19:30393101[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	31307588	+	chr19	31306230	+	.	8	1	6785730_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CATTCTCAG;MAPQ=0;MATEID=6785730_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=ACAC;SCTG=c_19_31286501_31311501_129C;SECONDARY;SPAN=1358;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:92 GQ:1.7 PL:[1.7, 0.0, 219.5] SR:1 DR:8 LR:-1.483 LO:15.0);ALT=]chr19:31307588]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	31951354	+	chr19	31955460	+	CAGATATTATTGTAACAATAATATAAACAATAGCAAGCTTTGACCCACTATGGTTAACTCAGGAAGATAGAATGGATTCAACATTAGCGAATCTATCTTATAATTAACTAACTTAAAAGATTGAACAGAAAAAAATGTGATAATCACAAAAGATGATAGATTTTAATATCCA	0	56	6787299_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TTCTT;INSERTION=CAGATATTATTGTAACAATAATATAAACAATAGCAAGCTTTGACCCACTATGGTTAACTCAGGAAGATAGAATGGATTCAACATTAGCGAATCTATCTTATAATTAACTAACTTAAAAGATTGAACAGAAAAAAATGTGATAATCACAAAAGATGATAGATTTTAATATCCA;MAPQ=60;MATEID=6787299_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_31948001_31973001_259C;SPAN=4106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:56 DP:36 GQ:15 PL:[165.0, 15.0, 0.0] SR:56 DR:0 LR:-165.0 LO:165.0);ALT=G[chr19:31955460[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	31951388	+	chr19	31955024	+	.	8	0	6787300_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6787300_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:31951388(+)-19:31955024(-)__19_31948001_31973001D;SPAN=3636;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=T[chr19:31955024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	33072234	+	chr19	33076721	+	.	10	0	6790136_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6790136_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:33072234(+)-19:33076721(-)__19_33075001_33100001D;SPAN=4487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:44 GQ:21.2 PL:[21.2, 0.0, 83.9] SR:0 DR:10 LR:-21.09 LO:23.3);ALT=G[chr19:33076721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34002064	+	chr19	34003498	+	.	0	16	6793244_1	29.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=6793244_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_33981501_34006501_351C;SPAN=1434;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:86 GQ:29.6 PL:[29.6, 0.0, 178.1] SR:16 DR:0 LR:-29.52 LO:35.7);ALT=G[chr19:34003498[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34003674	+	chr19	34012649	+	.	13	0	6793249_1	29.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6793249_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:34003674(+)-19:34012649(-)__19_33981501_34006501D;SPAN=8975;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:49 GQ:29.6 PL:[29.6, 0.0, 89.0] SR:0 DR:13 LR:-29.64 LO:31.3);ALT=A[chr19:34012649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34663668	+	chr19	34685381	+	.	10	11	6795239_1	47.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6795239_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_34643001_34668001_359C;SPAN=21713;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:43 GQ:47.9 PL:[47.9, 0.0, 54.5] SR:11 DR:10 LR:-47.77 LO:47.81);ALT=G[chr19:34685381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34710814	+	chr19	34712406	+	.	10	0	6795158_1	10.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=6795158_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:34710814(+)-19:34712406(-)__19_34692001_34717001D;SPAN=1592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:0 DR:10 LR:-9.982 LO:20.14);ALT=G[chr19:34712406[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34856237	+	chr19	34857685	+	.	18	0	6795685_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6795685_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:34856237(+)-19:34857685(-)__19_34839001_34864001D;SPAN=1448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:97 GQ:33.2 PL:[33.2, 0.0, 201.5] SR:0 DR:18 LR:-33.14 LO:40.14);ALT=C[chr19:34857685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34857341	+	chr19	34859486	+	CCAAGTCCAGGGGCGTGGAGGCCGCCCGGGAGCGGATGTTCAATGGTGAGAAGATCAACTACACCG	2	46	6795689_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=CCAAGTCCAGGGGCGTGGAGGCCGCCCGGGAGCGGATGTTCAATGGTGAGAAGATCAACTACACCG;MAPQ=60;MATEID=6795689_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_34839001_34864001_210C;SPAN=2145;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:96 GQ:99 PL:[125.9, 0.0, 106.1] SR:46 DR:2 LR:-125.9 LO:125.9);ALT=G[chr19:34859486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34857757	+	chr19	34859486	+	.	2	14	6795690_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6795690_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_34839001_34864001_210C;SPAN=1729;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:83 GQ:30.5 PL:[30.5, 0.0, 169.1] SR:14 DR:2 LR:-30.33 LO:35.97);ALT=G[chr19:34859486[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34884972	+	chr19	34887203	+	.	2	3	6795991_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6795991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_34863501_34888501_195C;SPAN=2231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:74 GQ:3.3 PL:[0.0, 3.3, 184.8] SR:3 DR:2 LR:3.543 LO:8.807);ALT=G[chr19:34887203[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34887562	+	chr19	34890110	+	.	4	3	6796001_1	12.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6796001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_34863501_34888501_380C;SPAN=2548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:38 GQ:12.8 PL:[12.8, 0.0, 78.8] SR:3 DR:4 LR:-12.81 LO:15.58);ALT=G[chr19:34890110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	34919475	+	chr19	34921480	+	.	14	16	6796291_1	48.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6796291_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_34912501_34937501_343C;SPAN=2005;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:90 GQ:48.2 PL:[48.2, 0.0, 170.3] SR:16 DR:14 LR:-48.24 LO:52.06);ALT=G[chr19:34921480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35491415	+	chr19	35500022	+	.	15	0	6797529_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6797529_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:35491415(+)-19:35500022(-)__19_35476001_35501001D;SPAN=8607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:67 GQ:31.4 PL:[31.4, 0.0, 130.4] SR:0 DR:15 LR:-31.36 LO:34.83);ALT=A[chr19:35500022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35645762	+	chr19	35651609	+	.	28	0	6798450_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6798450_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:35645762(+)-19:35651609(-)__19_35623001_35648001D;SPAN=5847;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:56 GQ:57.5 PL:[77.3, 0.0, 57.5] SR:0 DR:28 LR:-77.39 LO:77.39);ALT=G[chr19:35651609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35645772	+	chr19	35648322	+	ATGTCGCCCTCTGGTCGCCTGTGTCTTCTCACCATCGTTGGCCTGATTCTCCCCACCAG	73	73	6798452_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGTCGCCCTCTGGTCGCCTGTGTCTTCTCACCATCGTTGGCCTGATTCTCCCCACCAG;MAPQ=60;MATEID=6798452_2;MATENM=0;NM=1;NUMPARTS=3;SCTG=c_19_35623001_35648001_50C;SPAN=2550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:146 DP:53 GQ:39.4 PL:[432.4, 39.4, 0.0] SR:73 DR:73 LR:-432.4 LO:432.4);ALT=G[chr19:35648322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35648404	+	chr19	35651611	+	ATGCAGTCTACACAGAACTCCAGCCCACCTCTCCGACCCCAACCTGGCCTGCTGAT	0	191	6798290_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATGCAGTCTACACAGAACTCCAGCCCACCTCTCCGACCCCAACCTGGCCTGCTGAT;MAPQ=60;MATEID=6798290_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_35647501_35672501_155C;SPAN=3207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:191 DP:267 GQ:89.5 PL:[558.2, 0.0, 89.5] SR:191 DR:0 LR:-577.5 LO:577.5);ALT=G[chr19:35651611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35651704	+	chr19	35655056	+	.	2	43	6798297_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6798297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_35647501_35672501_204C;SPAN=3352;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:122 GQ:99 PL:[112.4, 0.0, 181.7] SR:43 DR:2 LR:-112.2 LO:113.1);ALT=G[chr19:35655056[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35655151	+	chr19	35657153	+	TTCATGAGGATGACCCCTTCTTCTAT	5	46	6798310_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;INSERTION=TTCATGAGGATGACCCCTTCTTCTAT;MAPQ=60;MATEID=6798310_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TT;SCTG=c_19_35647501_35672501_257C;SPAN=2002;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:98 GQ:99 PL:[128.6, 0.0, 108.8] SR:46 DR:5 LR:-128.7 LO:128.7);ALT=T[chr19:35657153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35655203	+	chr19	35660468	+	.	13	0	6798312_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6798312_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:35655203(+)-19:35660468(-)__19_35647501_35672501D;SPAN=5265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:102 GQ:15.5 PL:[15.5, 0.0, 230.0] SR:0 DR:13 LR:-15.28 LO:26.67);ALT=T[chr19:35660468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	35657231	+	chr19	35660469	+	TTCATGAGGATGACCCCTTCTTCTAT	14	44	6798320_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=GTG;INSERTION=TTCATGAGGATGACCCCTTCTTCTAT;MAPQ=60;MATEID=6798320_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_19_35647501_35672501_257C;SPAN=3238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:58 DP:120 GQ:99 PL:[158.9, 0.0, 132.5] SR:44 DR:14 LR:-159.1 LO:159.1);ALT=G[chr19:35660469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36139306	+	chr19	36145472	+	ATTCAGCACCATGGCGGAAGACATGGAGACCAAAATCAAGAACTACAAGACCGCCCCTTTTGACAGCCGCTTCCCCAACCAGAACCAGACTAGAAACTGCTGGCAGAACTACCTG	97	188	6800245_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATTCAGCACCATGGCGGAAGACATGGAGACCAAAATCAAGAACTACAAGACCGCCCCTTTTGACAGCCGCTTCCCCAACCAGAACCAGACTAGAAACTGCTGGCAGAACTACCTG;MAPQ=60;MATEID=6800245_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36137501_36162501_282C;SPAN=6166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:266 DP:218 GQ:71.8 PL:[788.8, 71.8, 0.0] SR:188 DR:97 LR:-788.9 LO:788.9);ALT=G[chr19:36145472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36139306	+	chr19	36142133	+	.	56	9	6800244_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6800244_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_36137501_36162501_282C;SPAN=2827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:159 GQ:79.1 PL:[306.8, 0.0, 79.1] SR:9 DR:56 LR:-314.3 LO:314.3);ALT=G[chr19:36142133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36139353	+	chr19	36149493	+	.	17	0	6800246_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6800246_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36139353(+)-19:36149493(-)__19_36137501_36162501D;SPAN=10140;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:172 GQ:9.7 PL:[9.7, 0.0, 405.8] SR:0 DR:17 LR:-9.518 LO:32.87);ALT=A[chr19:36149493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36142251	+	chr19	36145472	+	.	2	172	6800257_1	99.0	.	DISC_MAPQ=54;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6800257_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_19_36137501_36162501_282C;SPAN=3221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:174 DP:229 GQ:43.6 PL:[512.3, 0.0, 43.6] SR:172 DR:2 LR:-535.6 LO:535.6);ALT=G[chr19:36145472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36142253	+	chr19	36149495	+	.	3	2	6800258_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=6800258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_36137501_36162501_113C;SPAN=7242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:230 GQ:45.7 PL:[0.0, 45.7, 650.2] SR:2 DR:3 LR:45.81 LO:6.317);ALT=T[chr19:36149495[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36230671	+	chr19	36231924	+	.	0	5	6799891_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6799891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_36211001_36236001_225C;SPAN=1253;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:82 GQ:5.4 PL:[0.0, 5.4, 207.9] SR:5 DR:0 LR:5.711 LO:8.577);ALT=C[chr19:36231924[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36231023	+	chr19	36233290	+	.	18	0	6799893_1	34.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6799893_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36231023(+)-19:36233290(-)__19_36211001_36236001D;SPAN=2267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:92 GQ:34.7 PL:[34.7, 0.0, 186.5] SR:0 DR:18 LR:-34.49 LO:40.6);ALT=C[chr19:36233290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36232120	+	chr19	36233290	+	.	77	0	6799896_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6799896_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36232120(+)-19:36233290(-)__19_36211001_36236001D;SPAN=1170;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:87 GQ:20.1 PL:[250.8, 20.1, 0.0] SR:0 DR:77 LR:-251.3 LO:251.3);ALT=C[chr19:36233290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36233707	+	chr19	36234708	+	.	0	5	6799902_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=6799902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_36211001_36236001_52C;SPAN=1001;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:75 GQ:3.6 PL:[0.0, 3.6, 188.1] SR:5 DR:0 LR:3.814 LO:8.777);ALT=G[chr19:36234708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36393538	+	chr19	36394671	+	TGGCTGCAGCTCAGACGACTCCAGGAGAGAGATCATCACTCCCTGCCTTTTACCCTGGCACTT	0	164	6801065_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=TGGCTGCAGCTCAGACGACTCCAGGAGAGAGATCATCACTCCCTGCCTTTTACCCTGGCACTT;MAPQ=60;MATEID=6801065_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36382501_36407501_230C;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:164 DP:241 GQ:99 PL:[476.3, 0.0, 106.6] SR:164 DR:0 LR:-489.0 LO:489.0);ALT=G[chr19:36394671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36393600	+	chr19	36395019	+	.	15	0	6801067_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6801067_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36393600(+)-19:36395019(-)__19_36382501_36407501D;SPAN=1419;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:180 GQ:0.7 PL:[0.7, 0.0, 436.4] SR:0 DR:15 LR:-0.7486 LO:27.84);ALT=C[chr19:36395019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36395538	+	chr19	36398348	+	GATAAGGCGACTCGGTCTCAGTGATACGCTGTTTCCGGGTCGCTG	6	110	6801076_1	99.0	.	DISC_MAPQ=40;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GATAAGGCGACTCGGTCTCAGTGATACGCTGTTTCCGGGTCGCTG;MAPQ=60;MATEID=6801076_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36382501_36407501_142C;SPAN=2810;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:116 DP:580 GQ:99 PL:[225.8, 0.0, 1183.0] SR:110 DR:6 LR:-225.8 LO:262.9);ALT=T[chr19:36398348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36395585	+	chr19	36399110	+	.	8	0	6801078_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6801078_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:36395585(+)-19:36399110(-)__19_36382501_36407501D;SPAN=3525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:309 GQ:57.2 PL:[0.0, 57.2, 864.8] SR:0 DR:8 LR:57.31 LO:10.71);ALT=A[chr19:36399110[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36607088	+	chr19	36611612	+	.	0	28	6801864_1	65.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6801864_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_36603001_36628001_370C;SPAN=4524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:101 GQ:65.3 PL:[65.3, 0.0, 177.5] SR:28 DR:0 LR:-65.07 LO:68.06);ALT=T[chr19:36611612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36612622	+	chr19	36616566	+	CTCACAGATTTCAAGCCTGGCTACTGGATTGGTGTCCGCTATGATGAGCCACTGGGGAAAAATGATG	0	30	6801878_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GCAG;INSERTION=CTCACAGATTTCAAGCCTGGCTACTGGATTGGTGTCCGCTATGATGAGCCACTGGGGAAAAATGATG;MAPQ=60;MATEID=6801878_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36603001_36628001_63C;SPAN=3944;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:99 GQ:72.2 PL:[72.2, 0.0, 167.9] SR:30 DR:0 LR:-72.21 LO:74.32);ALT=T[chr19:36616566[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36632122	+	chr19	36633553	+	CGAGGCGGCTGCGCAGTACAACCCGGAGCCCCC	5	17	6801436_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CGAGGCGGCTGCGCAGTACAACCCGGAGCCCCC;MAPQ=60;MATEID=6801436_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36627501_36652501_277C;SECONDARY;SPAN=1431;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:90 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:17 DR:5 LR:-38.34 LO:43.57);ALT=G[chr19:36633553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36633644	+	chr19	36637096	+	ACATGGAGGTCAGCGCCACAGAACTCATGAACATTCTCAATAAGGTTGTGACACGACACCCTGATCTGAAGACTGATGGTTTTGGCATTGACACATGTCGCAGCATGGTGGCCGTGATGGATAGCGACACCACAGGCAAGCTGGGCTTTGAGGAATTCAAGTACTTGTGGAACAACATCAAAAGGTGGCAGGCCATATACAAACAGTTCGACACTGACCGATCAGGGACCATTTGCAGTAGTGAACTCCCAGGTGCCTTTGAGGCAGC	0	19	6801444_1	39.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ACATGGAGGTCAGCGCCACAGAACTCATGAACATTCTCAATAAGGTTGTGACACGACACCCTGATCTGAAGACTGATGGTTTTGGCATTGACACATGTCGCAGCATGGTGGCCGTGATGGATAGCGACACCACAGGCAAGCTGGGCTTTGAGGAATTCAAGTACTTGTGGAACAACATCAAAAGGTGGCAGGCCATATACAAACAGTTCGACACTGACCGATCAGGGACCATTTGCAGTAGTGAACTCCCAGGTGCCTTTGAGGCAGC;MAPQ=60;MATEID=6801444_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_19_36627501_36652501_251C;SPAN=3452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:85 GQ:39.8 PL:[39.8, 0.0, 165.2] SR:19 DR:0 LR:-39.69 LO:44.11);ALT=G[chr19:36637096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36637217	+	chr19	36640713	+	CCTTCAAATCTCTTGACAAAGATGGCACTGGACAAATCCAGGTGAACATCCAGG	32	35	6801457_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CCTTCAAATCTCTTGACAAAGATGGCACTGGACAAATCCAGGTGAACATCCAGG;MAPQ=60;MATEID=6801457_2;MATENM=2;NM=0;NUMPARTS=3;SCTG=c_19_36627501_36652501_378C;SPAN=3496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:90 GQ:71.3 PL:[147.2, 0.0, 71.3] SR:35 DR:32 LR:-148.7 LO:148.7);ALT=G[chr19:36640713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	36637217	+	chr19	36640480	+	.	10	11	6801456_1	38.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GTG;MAPQ=60;MATEID=6801456_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_36627501_36652501_378C;SPAN=3263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:91 GQ:38.3 PL:[38.3, 0.0, 180.2] SR:11 DR:10 LR:-38.07 LO:43.46);ALT=G[chr19:36640480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	37064429	+	chr19	37065721	+	.	11	4	6803152_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6803152_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_37044001_37069001_252C;SPAN=1292;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:74 GQ:23 PL:[23.0, 0.0, 155.0] SR:4 DR:11 LR:-22.86 LO:28.64);ALT=T[chr19:37065721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	37065804	+	chr19	37068042	+	.	0	7	6803158_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=6803158_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_19_37044001_37069001_320C;SPAN=2238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:7 DR:0 LR:1.818 LO:12.7);ALT=T[chr19:37068042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	37080653	+	chr19	37096098	+	.	11	0	6803448_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6803448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:37080653(+)-19:37096098(-)__19_37093001_37118001D;SPAN=15445;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:32 GQ:27.8 PL:[27.8, 0.0, 47.6] SR:0 DR:11 LR:-27.64 LO:28.0);ALT=C[chr19:37096098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	37660951	+	chr19	37663531	+	.	20	0	6805813_1	44.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6805813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:37660951(+)-19:37663531(-)__19_37656501_37681501D;SPAN=2580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:81 GQ:44.3 PL:[44.3, 0.0, 149.9] SR:0 DR:20 LR:-44.08 LO:47.43);ALT=A[chr19:37663531[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38343055	-	chr19	38344966	+	.	11	12	6808314_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6808314_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38342501_38367501_259C;SPAN=1911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:73 GQ:39.8 PL:[39.8, 0.0, 135.5] SR:12 DR:11 LR:-39.64 LO:42.67);ALT=[chr19:38344966[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	38755638	+	chr19	38778513	+	ACTTCTGCCTGGTGTCGAAGGTGGTGGGCAGATGCCGGGCCTCCATGCCTAGGTGGTGGTACAATGTCACTGACGGATCCTGCCAGCTGTTTGTGTATGGGGGCTGTGACGGAAACAGCAATAATTACCTGACCAAGGAGGAGTGCCTCAAGAAATGTGCCACTGTCA	2	14	6809869_1	42.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=ACTTCTGCCTGGTGTCGAAGGTGGTGGGCAGATGCCGGGCCTCCATGCCTAGGTGGTGGTACAATGTCACTGACGGATCCTGCCAGCTGTTTGTGTATGGGGGCTGTGACGGAAACAGCAATAATTACCTGACCAAGGAGGAGTGCCTCAAGAAATGTGCCACTGTCA;MAPQ=60;MATEID=6809869_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_38734501_38759501_122C;SPAN=22875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:39 GQ:42.2 PL:[42.2, 0.0, 52.1] SR:14 DR:2 LR:-42.25 LO:42.31);ALT=G[chr19:38778513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38755638	+	chr19	38774266	+	.	17	9	6809868_1	58.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6809868_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_38734501_38759501_122C;SPAN=18628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:39 GQ:35.6 PL:[58.7, 0.0, 35.6] SR:9 DR:17 LR:-59.05 LO:59.05);ALT=G[chr19:38774266[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38800319	+	chr19	38806356	+	.	80	0	6810009_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6810009_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:38800319(+)-19:38806356(-)__19_38783501_38808501D;SPAN=6037;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:97 GQ:3 PL:[240.9, 3.0, 0.0] SR:0 DR:80 LR:-253.2 LO:253.2);ALT=C[chr19:38806356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38865601	+	chr19	38866798	+	.	0	87	6810138_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6810138_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38857001_38882001_57C;SPAN=1197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:89 GQ:24 PL:[264.0, 24.0, 0.0] SR:87 DR:0 LR:-264.1 LO:264.1);ALT=G[chr19:38866798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38867095	+	chr19	38869880	+	.	2	6	6810142_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6810142_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38857001_38882001_204C;SPAN=2785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:6 DR:2 LR:-0.6203 LO:13.03);ALT=G[chr19:38869880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38870045	+	chr19	38871539	+	.	3	4	6810154_1	0	.	DISC_MAPQ=45;EVDNC=ASDIS;MAPQ=60;MATEID=6810154_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38857001_38882001_72C;SPAN=1494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:83 GQ:0.8 PL:[0.8, 0.0, 198.8] SR:4 DR:3 LR:-0.6203 LO:13.03);ALT=A[chr19:38871539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38871640	+	chr19	38872754	+	.	0	12	6810161_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6810161_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38857001_38882001_275C;SPAN=1114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:103 GQ:11.9 PL:[11.9, 0.0, 236.3] SR:12 DR:0 LR:-11.71 LO:24.11);ALT=G[chr19:38872754[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38872868	+	chr19	38873891	+	.	0	32	6810162_1	83.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6810162_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38857001_38882001_248C;SPAN=1023;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:81 GQ:83.9 PL:[83.9, 0.0, 110.3] SR:32 DR:0 LR:-83.69 LO:83.93);ALT=G[chr19:38873891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	38912795	+	chr19	38916708	+	.	17	4	6810288_1	41.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6810288_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_38906001_38931001_206C;SPAN=3913;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:80 GQ:41 PL:[41.0, 0.0, 153.2] SR:4 DR:17 LR:-41.05 LO:44.68);ALT=T[chr19:38916708[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	122804408	+	chr19	39044988	+	.	12	0	6811803_1	30.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6811803_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39044988(-)-23:122804408(+)__19_39028501_39053501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:33 GQ:30.8 PL:[30.8, 0.0, 47.3] SR:0 DR:12 LR:-30.67 LO:30.91);ALT=]chrX:122804408]A;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	39109979	+	chr19	39114716	+	.	81	0	6811129_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6811129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39109979(+)-19:39114716(-)__19_39102001_39127001D;SPAN=4737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:81 DP:125 GQ:68.6 PL:[233.6, 0.0, 68.6] SR:0 DR:81 LR:-238.4 LO:238.4);ALT=G[chr19:39114716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39111078	+	chr19	39114717	+	.	0	191	6811136_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=GTA;MAPQ=60;MATEID=6811136_2;MATENM=0;NM=0;NUMPARTS=6;SCTG=c_19_39102001_39127001_381C;SPAN=3639;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:191 DP:201 GQ:54.1 PL:[594.1, 54.1, 0.0] SR:191 DR:0 LR:-594.1 LO:594.1);ALT=A[chr19:39114717[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39123318	+	chr19	39125632	+	.	3	152	6811178_1	99.0	.	DISC_MAPQ=12;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6811178_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CAGCCAGC;SCTG=c_19_39102001_39127001_62C;SPAN=2314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:155 DP:257 GQ:83.1 PL:[240.7, 0.0, 83.1] SR:152 DR:3 LR:-246.0 LO:246.0);ALT=G[chr19:39125632[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39123318	+	chr19	39127529	+	ACAGCCAGCTAAAGGTGTGGATGAGCAAATACGGCTGGAGTGCCGACGAGTCGGGGCAGATCTTCATCTGTAGCCAAGAAGAGAGCATTAAACCCAAGAACATTGTGGAGAAGATTGACTTTGACA	8	217	6811179_1	99.0	.	DISC_MAPQ=20;EVDNC=TSI_G;HOMSEQ=GTG;INSERTION=ACAGCCAGCTAAAGGTGTGGATGAGCAAATACGGCTGGAGTGCCGACGAGTCGGGGCAGATCTTCATCTGTAGCCAAGAAGAGAGCATTAAACCCAAGAACATTGTGGAGAAGATTGACTTTGACA;MAPQ=60;MATEID=6811179_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_39102001_39127001_62C;SPAN=4211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:219 DP:115 GQ:59.2 PL:[650.2, 59.2, 0.0] SR:217 DR:8 LR:-650.3 LO:650.3);ALT=G[chr19:39127529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39125761	+	chr19	39127529	+	.	6	34	6811187_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GTG;MAPQ=60;MATEID=6811187_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_39102001_39127001_62C;SPAN=1768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:66 GQ:38.3 PL:[120.8, 0.0, 38.3] SR:34 DR:6 LR:-123.0 LO:123.0);ALT=G[chr19:39127529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39138547	+	chr19	39195572	+	ACCTTCACGGCATGGTGCAACTCCCACCTGCGGAAGGCAGGCACACAGATCGAGAACATTGATGAGGACTTCCGAGACGGGCTCAAGCTCATGCTGCTCCTGGAGGTCATATCAGGGGAGCGGTTACCTAAGCCGGAGCGGGGGAAGATGAGAGTGCACAAAATCAACAATGTGAACAAAGCGCTGGACTTTATTGCCAGCAAAGGCGTCAAGCTGGTCTCCATCGGGGCAGA	0	11	6810928_1	25.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ACCTTCACGGCATGGTGCAACTCCCACCTGCGGAAGGCAGGCACACAGATCGAGAACATTGATGAGGACTTCCGAGACGGGCTCAAGCTCATGCTGCTCCTGGAGGTCATATCAGGGGAGCGGTTACCTAAGCCGGAGCGGGGGAAGATGAGAGTGCACAAAATCAACAATGTGAACAAAGCGCTGGACTTTATTGCCAGCAAAGGCGTCAAGCTGGTCTCCATCGGGGCAGA;MAPQ=60;MATEID=6810928_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_39175501_39200501_260C;SPAN=57025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:40 GQ:25.4 PL:[25.4, 0.0, 71.6] SR:11 DR:0 LR:-25.47 LO:26.69);ALT=G[chr19:39195572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39138547	+	chr19	39191238	+	.	9	7	6810927_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6810927_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_19_39175501_39200501_260C;SPAN=52691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:50 GQ:29.3 PL:[29.3, 0.0, 92.0] SR:7 DR:9 LR:-29.37 LO:31.17);ALT=G[chr19:39191238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39308218	+	chr19	39321715	+	.	3	17	6812067_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TACCTG;MAPQ=60;MATEID=6812067_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_39298001_39323001_162C;SPAN=13497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:84 GQ:43.4 PL:[43.4, 0.0, 158.9] SR:17 DR:3 LR:-43.26 LO:47.06);ALT=G[chr19:39321715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39336746	+	chr19	39342934	+	.	14	0	6811979_1	29.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=6811979_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39336746(+)-19:39342934(-)__19_39322501_39347501D;SPAN=6188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:61 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:0 DR:14 LR:-29.69 LO:32.68);ALT=C[chr19:39342934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39338075	+	chr19	39340339	+	.	0	10	6811982_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6811982_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_39322501_39347501_183C;SPAN=2264;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:10 DR:0 LR:-9.44 LO:20.03);ALT=C[chr19:39340339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39380601	+	chr19	39384052	+	ATGTGGAGATTCCAGCTCCCACCAAACAGATGACTCTGCG	0	14	6811874_1	20.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AC;INSERTION=ATGTGGAGATTCCAGCTCCCACCAAACAGATGACTCTGCG;MAPQ=60;MATEID=6811874_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_39371501_39396501_379C;SPAN=3451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:96 GQ:20.3 PL:[20.3, 0.0, 211.7] SR:14 DR:0 LR:-20.21 LO:29.6);ALT=G[chr19:39384052[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39380842	+	chr19	39390144	+	.	9	0	6811876_1	5.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6811876_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39380842(+)-19:39390144(-)__19_39371501_39396501D;SPAN=9302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:91 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.055 LO:17.41);ALT=A[chr19:39390144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39384167	+	chr19	39390145	+	TGTCTGCTTCTCCACCAGCGGCTCCTCCCTCAGAGTCTGAATCTGAGT	16	15	6811888_1	58.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TGTCTGCTTCTCCACCAGCGGCTCCTCCCTCAGAGTCTGAATCTGAGT;MAPQ=60;MATEID=6811888_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_39371501_39396501_110C;SPAN=5978;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:88 GQ:58.7 PL:[58.7, 0.0, 154.4] SR:15 DR:16 LR:-58.68 LO:61.08);ALT=A[chr19:39390145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39384563	+	chr19	39390163	+	.	10	0	6811893_1	9.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6811893_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39384563(+)-19:39390163(-)__19_39371501_39396501D;SPAN=5600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:86 GQ:9.8 PL:[9.8, 0.0, 197.9] SR:0 DR:10 LR:-9.711 LO:20.09);ALT=A[chr19:39390163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39469983	+	chr19	39471117	-	.	8	0	6812399_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6812399_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39469983(+)-19:39471117(+)__19_39445001_39470001D;SPAN=1134;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:0 DR:8 LR:-11.78 LO:16.98);ALT=G]chr19:39471117];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	39819755	+	chr19	39826611	+	.	10	0	6813749_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6813749_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39819755(+)-19:39826611(-)__19_39812501_39837501D;SPAN=6856;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:160 GQ:10.3 PL:[0.0, 10.3, 409.3] SR:0 DR:10 LR:10.34 LO:17.26);ALT=G[chr19:39826611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39820268	+	chr19	39826075	+	GGGCTGTCTCTCCGGCAACTCCATTTTGAGCTCCTCTGGGGAAATGTT	10	45	6813753_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=GGGCTGTCTCTCCGGCAACTCCATTTTGAGCTCCTCTGGGGAAATGTT;MAPQ=60;MATEID=6813753_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_39812501_39837501_145C;SPAN=5807;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:162 GQ:99 PL:[131.3, 0.0, 260.0] SR:45 DR:10 LR:-131.1 LO:133.5);ALT=T[chr19:39826075[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39820312	+	chr19	39826613	+	.	45	0	6813754_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6813754_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39820312(+)-19:39826613(-)__19_39812501_39837501D;SPAN=6301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:176 GQ:99 PL:[101.0, 0.0, 325.4] SR:0 DR:45 LR:-100.9 LO:107.5);ALT=A[chr19:39826613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39824149	+	chr19	39826613	+	.	67	0	6813771_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6813771_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39824149(+)-19:39826613(-)__19_39812501_39837501D;SPAN=2464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:170 GQ:99 PL:[175.1, 0.0, 237.8] SR:0 DR:67 LR:-175.1 LO:175.6);ALT=G[chr19:39826613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39877442	+	chr19	39878978	+	.	4	5	6813840_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6813840_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_39861501_39886501_20C;SPAN=1536;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:5 DR:4 LR:-6.631 LO:15.85);ALT=G[chr19:39878978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39924403	+	chr19	39926247	+	.	0	132	6814129_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6814129_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_39910501_39935501_82C;SPAN=1844;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:132 DP:435 GQ:99 PL:[318.0, 0.0, 737.2] SR:132 DR:0 LR:-317.9 LO:327.1);ALT=T[chr19:39926247[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39924437	+	chr19	39926494	+	.	78	0	6814131_1	99.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=6814131_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:39924437(+)-19:39926494(-)__19_39910501_39935501D;SPAN=2057;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:123 GQ:72.5 PL:[224.3, 0.0, 72.5] SR:0 DR:78 LR:-228.3 LO:228.3);ALT=C[chr19:39926494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39936607	+	chr19	39943994	+	.	6	8	6813974_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6813974_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_39935001_39960001_11C;SPAN=7387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:82 GQ:17.6 PL:[17.6, 0.0, 179.3] SR:8 DR:6 LR:-17.4 LO:25.39);ALT=T[chr19:39943994[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	39979286	+	chr19	39980356	+	.	0	12	6814268_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6814268_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_39959501_39984501_106C;SPAN=1070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:107 GQ:10.7 PL:[10.7, 0.0, 248.3] SR:12 DR:0 LR:-10.62 LO:23.9);ALT=G[chr19:39980356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40325455	+	chr19	40327195	+	.	6	63	6815048_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=6815048_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=AA;SCTG=c_19_40302501_40327501_335C;SPAN=1740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:133 GQ:99 PL:[185.3, 0.0, 135.8] SR:63 DR:6 LR:-185.5 LO:185.5);ALT=T[chr19:40327195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40327309	+	chr19	40328351	+	.	4	21	6815072_1	53.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=6815072_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_40327001_40352001_249C;SPAN=1042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:106 GQ:53.9 PL:[53.9, 0.0, 202.4] SR:21 DR:4 LR:-53.81 LO:58.7);ALT=C[chr19:40328351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40328484	+	chr19	40329674	+	.	8	9	6815073_1	22.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=6815073_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=CC;SCTG=c_19_40327001_40352001_249C;SPAN=1190;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:89 GQ:22.1 PL:[22.1, 0.0, 193.7] SR:9 DR:8 LR:-22.1 LO:30.11);ALT=C[chr19:40329674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40329846	+	chr19	40330872	+	.	11	10	6815082_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6815082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40327001_40352001_160C;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:81 GQ:31.1 PL:[31.1, 0.0, 163.1] SR:10 DR:11 LR:-30.87 LO:36.16);ALT=C[chr19:40330872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40331430	+	chr19	40336930	+	.	186	12	6815089_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6815089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40327001_40352001_248C;SPAN=5500;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:193 DP:91 GQ:52 PL:[571.0, 52.0, 0.0] SR:12 DR:186 LR:-571.0 LO:571.0);ALT=G[chr19:40336930[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40477186	+	chr19	40478273	+	.	23	0	6815847_1	49.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6815847_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:40477186(+)-19:40478273(-)__19_40474001_40499001D;SPAN=1087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:97 GQ:49.7 PL:[49.7, 0.0, 185.0] SR:0 DR:23 LR:-49.64 LO:54.07);ALT=G[chr19:40478273[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40771261	+	chr19	40791088	+	.	8	8	6816593_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6816593_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_40768001_40793001_186C;SPAN=19827;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:86 GQ:19.7 PL:[19.7, 0.0, 188.0] SR:8 DR:8 LR:-19.61 LO:27.71);ALT=G[chr19:40791088[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40854678	+	chr19	40871458	+	.	38	2	6817119_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=6817119_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40841501_40866501_234C;SPAN=16780;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:56 GQ:17.9 PL:[116.9, 0.0, 17.9] SR:2 DR:38 LR:-120.9 LO:120.9);ALT=A[chr19:40871458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40854693	+	chr19	40871784	+	.	9	0	6817120_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6817120_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:40854693(+)-19:40871784(-)__19_40841501_40866501D;SPAN=17091;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:0 DR:9 LR:-14.54 LO:19.45);ALT=G[chr19:40871784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40854693	+	chr19	40872513	+	.	14	0	6817121_1	31.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6817121_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:40854693(+)-19:40872513(-)__19_40841501_40866501D;SPAN=17820;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:56 GQ:31.1 PL:[31.1, 0.0, 103.7] SR:0 DR:14 LR:-31.04 LO:33.29);ALT=G[chr19:40872513[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40877780	+	chr19	40880387	+	.	5	4	6816922_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6816922_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40866001_40891001_333C;SPAN=2607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:98 GQ:3.3 PL:[0.0, 3.3, 244.2] SR:4 DR:5 LR:3.444 LO:12.5);ALT=G[chr19:40880387[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40882681	+	chr19	40883692	+	.	0	6	6816946_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6816946_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40866001_40891001_239C;SPAN=1011;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:84 GQ:2.7 PL:[0.0, 2.7, 207.9] SR:6 DR:0 LR:2.952 LO:10.72);ALT=G[chr19:40883692[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40929455	+	chr19	40931774	+	.	0	10	6817006_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6817006_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_40915001_40940001_59C;SPAN=2319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:10 DR:0 LR:-14.59 LO:21.18);ALT=T[chr19:40931774[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40948021	+	chr19	40950139	+	.	16	0	6817208_1	28.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6817208_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:40948021(+)-19:40950139(-)__19_40939501_40964501D;SPAN=2118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:92 GQ:28.1 PL:[28.1, 0.0, 193.1] SR:0 DR:16 LR:-27.89 LO:35.18);ALT=A[chr19:40950139[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40953958	+	chr19	40957270	+	.	2	37	6817222_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTATG;MAPQ=60;MATEID=6817222_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40939501_40964501_32C;SPAN=3312;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:97 GQ:99 PL:[102.5, 0.0, 132.2] SR:37 DR:2 LR:-102.5 LO:102.7);ALT=G[chr19:40957270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40957400	+	chr19	40964062	+	.	0	9	6817276_1	18.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6817276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40964001_40989001_307C;SPAN=6662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:43 GQ:18.2 PL:[18.2, 0.0, 84.2] SR:9 DR:0 LR:-18.06 LO:20.6);ALT=C[chr19:40964062[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	40964455	+	chr19	40971516	+	.	85	41	6817279_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6817279_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_40964001_40989001_233C;SPAN=7061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:102 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:41 DR:85 LR:-303.7 LO:303.7);ALT=G[chr19:40971516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41086843	+	chr19	41088255	+	.	2	4	6817745_1	0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6817745_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41086501_41111501_274C;SPAN=1412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:95 GQ:9 PL:[0.0, 9.0, 247.5] SR:4 DR:2 LR:9.233 LO:8.25);ALT=G[chr19:41088255[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41257386	+	chr19	41263236	+	.	22	38	6818352_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6818352_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41258001_41283001_153C;SPAN=5850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:45 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:38 DR:22 LR:-132.0 LO:132.0);ALT=G[chr19:41263236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41263409	+	chr19	41265335	+	.	4	3	6818368_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6818368_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41258001_41283001_159C;SPAN=1926;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:78 GQ:1.2 PL:[0.0, 1.2, 191.4] SR:3 DR:4 LR:1.326 LO:10.92);ALT=G[chr19:41265335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41265516	+	chr19	41268805	+	.	6	5	6818373_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6818373_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41258001_41283001_140C;SPAN=3289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:90 GQ:2 PL:[2.0, 0.0, 216.5] SR:5 DR:6 LR:-2.025 LO:15.08);ALT=G[chr19:41268805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41269582	+	chr19	41270913	+	.	3	4	6818383_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=6818383_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41258001_41283001_133C;SPAN=1331;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:92 GQ:1.5 PL:[0.0, 1.5, 224.4] SR:4 DR:3 LR:1.818 LO:12.7);ALT=T[chr19:41270913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41284296	+	chr19	41285923	+	.	6	3	6818439_1	2.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6818439_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41282501_41307501_233C;SPAN=1627;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:78 GQ:2 PL:[2.0, 0.0, 186.8] SR:3 DR:6 LR:-1.975 LO:13.23);ALT=G[chr19:41285923[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41305208	+	chr19	41306242	+	.	20	0	6818505_1	50.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6818505_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41305208(+)-19:41306242(-)__19_41282501_41307501D;SPAN=1034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:58 GQ:50.3 PL:[50.3, 0.0, 89.9] SR:0 DR:20 LR:-50.31 LO:50.93);ALT=A[chr19:41306242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41608725	+	chr19	41610191	+	.	15	11	6819489_1	56.0	.	DISC_MAPQ=39;EVDNC=ASDIS;HOMSEQ=AGAAAACCCCAACATCTC;MAPQ=60;MATEID=6819489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41601001_41626001_271C;SPAN=1466;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:74 GQ:56 PL:[56.0, 0.0, 122.0] SR:11 DR:15 LR:-55.88 LO:57.29);ALT=C[chr19:41610191[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41810166	+	chr19	41811578	+	.	0	5	6820106_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6820106_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41797001_41822001_144C;SPAN=1412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:97 GQ:9.6 PL:[0.0, 9.6, 254.1] SR:5 DR:0 LR:9.775 LO:8.204);ALT=G[chr19:41811578[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41816262	+	chr19	41822288	+	.	10	6	6820230_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6820230_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41821501_41846501_113C;SPAN=6026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:43 GQ:34.7 PL:[34.7, 0.0, 67.7] SR:6 DR:10 LR:-34.56 LO:35.22);ALT=G[chr19:41822288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41837117	+	chr19	41847788	+	TGCTGTACTGCGTGTCCAGGCTCCAAATGTAGGGGCAGGGCCCGAGGCAGAAGTTGGCATGGTAGCCCTTGGGCTCGTGGATCCACTTCCAGCCGAGGTCCTTGCGGAAGTCAATGTACAGCTGCCGCACGCAGCAGTTCTTCTCCGTGGAG	2	53	6820271_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TGCTGTACTGCGTGTCCAGGCTCCAAATGTAGGGGCAGGGCCCGAGGCAGAAGTTGGCATGGTAGCCCTTGGGCTCGTGGATCCACTTCCAGCCGAGGTCCTTGCGGAAGTCAATGTACAGCTGCCGCACGCAGCAGTTCTTCTCCGTGGAG;MAPQ=60;MATEID=6820271_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_41821501_41846501_319C;SPAN=10671;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:51 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:53 DR:2 LR:-155.1 LO:155.1);ALT=T[chr19:41847788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41838189	+	chr19	41847788	+	.	20	12	6820336_1	89.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6820336_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_41846001_41871001_93C;SPAN=9599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:27 DP:31 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:12 DR:20 LR:-87.4 LO:87.4);ALT=G[chr19:41847788[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41848154	+	chr19	41850651	+	.	0	12	6820350_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6820350_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41846001_41871001_7C;SPAN=2497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:100 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:12 DR:0 LR:-12.52 LO:24.28);ALT=T[chr19:41850651[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41848196	+	chr19	41854200	+	.	10	0	6820351_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6820351_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41848196(+)-19:41854200(-)__19_41846001_41871001D;SPAN=6004;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:84 GQ:10.4 PL:[10.4, 0.0, 191.9] SR:0 DR:10 LR:-10.25 LO:20.2);ALT=A[chr19:41854200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41850771	+	chr19	41854200	+	.	15	15	6820365_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6820365_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41846001_41871001_80C;SPAN=3429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:83 GQ:53.6 PL:[53.6, 0.0, 146.0] SR:15 DR:15 LR:-53.44 LO:55.9);ALT=T[chr19:41854200[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41850808	+	chr19	41858594	+	.	8	0	6820366_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6820366_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41850808(+)-19:41858594(-)__19_41846001_41871001D;SPAN=7786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=A[chr19:41858594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41854369	+	chr19	41858594	+	.	8	0	6820380_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6820380_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:41854369(+)-19:41858594(-)__19_41846001_41871001D;SPAN=4225;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:75 GQ:6.2 PL:[6.2, 0.0, 174.5] SR:0 DR:8 LR:-6.089 LO:15.75);ALT=G[chr19:41858594[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41863930	+	chr19	41869862	+	TGTGAATGCCCCACTTGCAGAAGAGGCTACTTTCCGAGAAACCGCTGGCCCCTATGATCTGCCCGATCACGTGCACCTCAGCCATGGC	0	10	6820410_1	10.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TGTGAATGCCCCACTTGCAGAAGAGGCTACTTTCCGAGAAACCGCTGGCCCCTATGATCTGCCCGATCACGTGCACCTCAGCCATGGC;MAPQ=60;MATEID=6820410_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_41846001_41871001_23C;SPAN=5932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:85 GQ:10.1 PL:[10.1, 0.0, 194.9] SR:10 DR:0 LR:-9.982 LO:20.14);ALT=G[chr19:41869862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41870001	+	chr19	41884186	+	.	10	3	6820774_1	22.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6820774_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41870501_41895501_142C;SPAN=14185;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:39 GQ:22.4 PL:[22.4, 0.0, 71.9] SR:3 DR:10 LR:-22.44 LO:23.91);ALT=G[chr19:41884186[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41882760	+	chr19	41884185	+	.	4	4	6820816_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6820816_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_41870501_41895501_103C;SPAN=1425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:69 GQ:4.4 PL:[4.4, 0.0, 162.8] SR:4 DR:4 LR:-4.413 LO:13.62);ALT=G[chr19:41884185[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41884425	+	chr19	41888675	+	.	0	8	6820822_1	4.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6820822_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41870501_41895501_120C;SPAN=4250;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:83 GQ:4.1 PL:[4.1, 0.0, 195.5] SR:8 DR:0 LR:-3.921 LO:15.38);ALT=G[chr19:41888675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41898887	+	chr19	41903084	+	.	0	34	6820640_1	85.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6820640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41895001_41920001_259C;SPAN=4197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:101 GQ:85.1 PL:[85.1, 0.0, 157.7] SR:34 DR:0 LR:-84.87 LO:86.14);ALT=T[chr19:41903084[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41903840	+	chr19	41916550	+	CACCCCCA	37	10	6820662_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CACCCCCA;MAPQ=60;MATEID=6820662_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41895001_41920001_221C;SPAN=12710;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:97 GQ:99 PL:[109.1, 0.0, 125.6] SR:10 DR:37 LR:-109.1 LO:109.1);ALT=T[chr19:41916550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41929078	+	chr19	41930341	+	.	4	3	6820568_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTGA;MAPQ=60;MATEID=6820568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41919501_41944501_246C;SPAN=1263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:98 GQ:3.3 PL:[0.0, 3.3, 244.2] SR:3 DR:4 LR:3.444 LO:12.5);ALT=A[chr19:41930341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	41942378	+	chr19	41944123	+	.	0	8	6820618_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6820618_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_41919501_41944501_21C;SPAN=1745;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:8 DR:0 LR:2.581 LO:14.46);ALT=C[chr19:41944123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42364592	+	chr19	42373099	+	.	29	0	6822031_1	24.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6822031_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:42364592(+)-19:42373099(-)__19_42360501_42385501D;SPAN=8507;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:264 GQ:24.4 PL:[24.4, 0.0, 615.2] SR:0 DR:29 LR:-24.21 LO:57.49);ALT=C[chr19:42373099[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42364949	+	chr19	42373133	+	.	18	0	6822032_1	0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6822032_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:42364949(+)-19:42373133(-)__19_42360501_42385501D;SPAN=8184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:18 DP:1127 GQ:99 PL:[0.0, 245.6, 3228.0] SR:0 DR:18 LR:245.9 LO:20.36);ALT=A[chr19:42373133[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42387390	+	chr19	42392130	+	.	17	0	6821841_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6821841_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:42387390(+)-19:42392130(-)__19_42385001_42410001D;SPAN=4740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:64 GQ:38.9 PL:[38.9, 0.0, 114.8] SR:0 DR:17 LR:-38.78 LO:40.95);ALT=C[chr19:42392130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42387405	+	chr19	42392822	+	.	20	0	6821842_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6821842_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:42387405(+)-19:42392822(-)__19_42385001_42410001D;SPAN=5417;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:87 GQ:42.5 PL:[42.5, 0.0, 167.9] SR:0 DR:20 LR:-42.45 LO:46.71);ALT=G[chr19:42392822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42392936	+	chr19	42396095	+	.	2	3	6821854_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6821854_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_42385001_42410001_304C;SPAN=3159;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:88 GQ:7.2 PL:[0.0, 7.2, 227.7] SR:3 DR:2 LR:7.336 LO:8.42);ALT=G[chr19:42396095[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42461272	+	chr19	42462887	+	AAAGAGCACAAGCTTGGACTCCAAGGTGCGCAGATAGAGAATGTAACAGGCGCCGAAAAAGACAGCCAGAGCCACCAGCAACATAGGGGACGTCAC	2	75	6822312_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AAAGAGCACAAGCTTGGACTCCAAGGTGCGCAGATAGAGAATGTAACAGGCGCCGAAAAAGACAGCCAGAGCCACCAGCAACATAGGGGACGTCAC;MAPQ=60;MATEID=6822312_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_42458501_42483501_314C;SPAN=1615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:76 DP:106 GQ:34.1 PL:[222.2, 0.0, 34.1] SR:75 DR:2 LR:-229.9 LO:229.9);ALT=C[chr19:42462887[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42461272	+	chr19	42462437	+	.	2	16	6822311_1	36.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=6822311_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_19_42458501_42483501_314C;SPAN=1165;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:86 GQ:36.2 PL:[36.2, 0.0, 171.5] SR:16 DR:2 LR:-36.12 LO:41.2);ALT=C[chr19:42462437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42621520	+	chr19	42626663	+	TTGTACTGGGGCCAGTTGGGGACACGGAGAATGGGGAGGTCTTATTTTGGGGGTTCTGATGATTAGTGTCTGGTCCATTTCTTTCGGTGT	0	11	6822725_1	10.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TTGTACTGGGGCCAGTTGGGGACACGGAGAATGGGGAGGTCTTATTTTGGGGGTTCTGATGATTAGTGTCTGGTCCATTTCTTTCGGTGT;MAPQ=60;MATEID=6822725_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_42605501_42630501_47C;SPAN=5143;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:96 GQ:10.4 PL:[10.4, 0.0, 221.6] SR:11 DR:0 LR:-10.3 LO:22.02);ALT=T[chr19:42626663[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42626938	+	chr19	42636535	+	.	9	0	6822835_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6822835_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:42626938(+)-19:42636535(-)__19_42630001_42655001D;SPAN=9597;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=G[chr19:42636535[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	42804441	+	chr19	42806102	+	.	0	10	6823271_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6823271_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_42801501_42826501_346C;SPAN=1661;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:87 GQ:9.5 PL:[9.5, 0.0, 200.9] SR:10 DR:0 LR:-9.44 LO:20.03);ALT=T[chr19:42806102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	43367095	+	chr19	43253495	+	.	17	0	6825144_1	43.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6825144_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:43253495(-)-19:43367095(+)__19_43242501_43267501D;SPAN=113600;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:47 GQ:43.4 PL:[43.4, 0.0, 69.8] SR:0 DR:17 LR:-43.38 LO:43.74);ALT=]chr19:43367095]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	149032062	+	chr19	43993142	+	.	16	17	7552851_1	92.0	.	DISC_MAPQ=1;EVDNC=ASDIS;HOMSEQ=GGGTTTCACCATATTGGCCAGGCTGGTCTCAAATTCCTGACTTCAAGTGATC;MAPQ=44;MATEID=7552851_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_23_149009001_149034001_168C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:6 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:17 DR:16 LR:-92.42 LO:92.42);ALT=]chrX:149032062]G;VARTYPE=BND:TRX-th;JOINTYPE=th
chr19	44011056	+	chr19	44012096	+	.	0	62	6828117_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6828117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_44002001_44027001_383C;SPAN=1040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:105 GQ:77.3 PL:[176.3, 0.0, 77.3] SR:62 DR:0 LR:-178.2 LO:178.2);ALT=T[chr19:44012096[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44013018	+	chr19	44015588	+	.	0	7	6828126_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6828126_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_44002001_44027001_403C;SPAN=2570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:86 GQ:0 PL:[0.0, 0.0, 207.9] SR:7 DR:0 LR:0.1925 LO:12.92);ALT=T[chr19:44015588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44015718	+	chr19	44030667	+	GAAGCGCCCGAAGCGGATGGAGTCTCCATCCTCAATGTGTAAGTCAGCCTGGGCCCCACTAAGGCGGGAGATGACAGACTGGCAGCCAGGGAGGAGGGAACGGAGCAGCCCCGAGCCTGTAATGTGGTCCGCGTGGCAGTGGGTATTCA	0	67	6828134_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GAAGCGCCCGAAGCGGATGGAGTCTCCATCCTCAATGTGTAAGTCAGCCTGGGCCCCACTAAGGCGGGAGATGACAGACTGGCAGCCAGGGAGGAGGGAACGGAGCAGCCCCGAGCCTGTAATGTGGTCCGCGTGGCAGTGGGTATTCA;MAPQ=60;MATEID=6828134_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_44002001_44027001_210C;SPAN=14949;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:67 DP:47 GQ:18 PL:[198.0, 18.0, 0.0] SR:67 DR:0 LR:-198.0 LO:198.0);ALT=C[chr19:44030667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44112263	+	chr19	44118380	+	.	0	46	6827548_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCTGG;MAPQ=60;MATEID=6827548_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_44100001_44125001_160C;SPAN=6117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:110 GQ:99 PL:[122.0, 0.0, 145.1] SR:46 DR:0 LR:-122.0 LO:122.2);ALT=G[chr19:44118380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44112310	+	chr19	44123709	+	.	26	0	6827550_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6827550_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:44112310(+)-19:44123709(-)__19_44100001_44125001D;SPAN=11399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:101 GQ:58.7 PL:[58.7, 0.0, 184.1] SR:0 DR:26 LR:-58.46 LO:62.21);ALT=A[chr19:44123709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44118603	+	chr19	44123709	+	.	87	0	6827570_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6827570_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:44118603(+)-19:44123709(-)__19_44100001_44125001D;SPAN=5106;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:88 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:0 DR:87 LR:-260.8 LO:260.8);ALT=G[chr19:44123709[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44169613	+	chr19	44171733	+	.	0	14	6828447_1	17.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=6828447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_44149001_44174001_454C;SPAN=2120;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:108 GQ:17 PL:[17.0, 0.0, 244.7] SR:14 DR:0 LR:-16.95 LO:28.83);ALT=T[chr19:44171733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44169659	+	chr19	44174239	+	.	8	0	6828448_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6828448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:44169659(+)-19:44174239(-)__19_44149001_44174001D;SPAN=4580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:43 GQ:14.9 PL:[14.9, 0.0, 87.5] SR:0 DR:8 LR:-14.76 LO:17.85);ALT=C[chr19:44174239[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	44171848	+	chr19	44174218	+	.	22	9	6828458_1	64.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTGGG;MAPQ=60;MATEID=6828458_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_44149001_44174001_83C;SPAN=2370;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:55 GQ:64.4 PL:[64.4, 0.0, 67.7] SR:9 DR:22 LR:-64.32 LO:64.33);ALT=G[chr19:44174218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45449371	+	chr19	45451920	+	.	8	0	6831779_1	2.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6831779_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45449371(+)-19:45451920(-)__19_45447501_45472501D;SPAN=2549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:88 GQ:2.6 PL:[2.6, 0.0, 210.5] SR:0 DR:8 LR:-2.567 LO:15.16);ALT=C[chr19:45451920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45458730	+	chr19	45465236	+	.	8	0	6831822_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6831822_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45458730(+)-19:45465236(-)__19_45447501_45472501D;SPAN=6506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:85 GQ:3.5 PL:[3.5, 0.0, 201.5] SR:0 DR:8 LR:-3.379 LO:15.29);ALT=G[chr19:45465236[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45504944	+	chr19	45506205	+	.	0	37	6832116_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6832116_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45496501_45521501_287C;SPAN=1261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:78 GQ:87.8 PL:[101.0, 0.0, 87.8] SR:37 DR:0 LR:-101.0 LO:101.0);ALT=G[chr19:45506205[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45542419	+	chr19	45543438	+	.	14	0	6832315_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6832315_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45542419(+)-19:45543438(-)__19_45521001_45546001D;SPAN=1019;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:83 GQ:23.9 PL:[23.9, 0.0, 175.7] SR:0 DR:14 LR:-23.73 LO:30.57);ALT=G[chr19:45543438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45542419	+	chr19	45555328	+	.	10	0	6832316_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6832316_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45542419(+)-19:45555328(-)__19_45521001_45546001D;SPAN=12909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=G[chr19:45555328[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45543569	+	chr19	45556049	+	AAGAAGGACCCAGCCCAGTTCCTGCAGGTACATGGCCGAGCTTGCAAGGTGCACCTGGATTCTGCAGTCGCCCTGGCCGCTGAGAGCCCTGTTAATAT	0	19	6832319_1	52.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=AAGAAGGACCCAGCCCAGTTCCTGCAGGTACATGGCCGAGCTTGCAAGGTGCACCTGGATTCTGCAGTCGCCCTGGCCGCTGAGAGCCCTGTTAATAT;MAPQ=60;MATEID=6832319_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_45521001_45546001_31C;SPAN=12480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:38 GQ:39.2 PL:[52.4, 0.0, 39.2] SR:19 DR:0 LR:-52.52 LO:52.52);ALT=C[chr19:45556049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45579083	+	chr19	45583163	+	.	6	3	6832370_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTC;MAPQ=60;MATEID=6832370_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45570001_45595001_137C;SPAN=4080;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:82 GQ:1.1 PL:[1.1, 0.0, 195.8] SR:3 DR:6 LR:-0.8912 LO:13.07);ALT=C[chr19:45583163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45583287	+	chr19	45593363	+	.	3	4	6832376_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6832376_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45570001_45595001_285C;SPAN=10076;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:90 GQ:7.8 PL:[0.0, 7.8, 234.3] SR:4 DR:3 LR:7.878 LO:8.37);ALT=G[chr19:45593363[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45667590	+	chr19	45681413	+	.	17	0	6832757_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6832757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45667590(+)-19:45681413(-)__19_45668001_45693001D;SPAN=13823;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:67 GQ:38 PL:[38.0, 0.0, 123.8] SR:0 DR:17 LR:-37.97 LO:40.55);ALT=A[chr19:45681413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45668229	+	chr19	45681392	+	.	77	3	6832621_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6832621_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45643501_45668501_27C;SPAN=13163;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:79 DP:61 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:3 DR:77 LR:-234.4 LO:234.4);ALT=C[chr19:45681392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45668453	+	chr19	45681392	+	.	33	9	6832761_1	81.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6832761_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45668001_45693001_348C;SPAN=12939;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:115 GQ:81.2 PL:[81.2, 0.0, 196.7] SR:9 DR:33 LR:-81.08 LO:83.78);ALT=C[chr19:45681392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45912983	+	chr19	45916934	+	.	3	24	6833671_1	75.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6833671_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45888501_45913501_414C;SPAN=3951;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:37 GQ:13.1 PL:[75.8, 0.0, 13.1] SR:24 DR:3 LR:-78.22 LO:78.22);ALT=C[chr19:45916934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45917003	+	chr19	45918115	+	TCCAAATGTGGTCAGGAGGGTCTGACTGTCCGTTTTGTTGACTGACTTCACGGTGGTCAGACATTCAG	0	51	6833937_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=TCACC;INSERTION=TCCAAATGTGGTCAGGAGGGTCTGACTGTCCGTTTTGTTGACTGACTTCACGGTGGTCAGACATTCAG;MAPQ=60;MATEID=6833937_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_45913001_45938001_359C;SPAN=1112;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:99 GQ:98.6 PL:[141.5, 0.0, 98.6] SR:51 DR:0 LR:-141.9 LO:141.9);ALT=A[chr19:45918115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45918220	+	chr19	45922356	+	CCAGGCGAGGATCAATGTGCAGTCGGCCAGGATACACATCTTAGCCAGCTCCTTGAGGGCCTGCTGGGGATCTTT	0	15	6833945_1	24.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CCAGGCGAGGATCAATGTGCAGTCGGCCAGGATACACATCTTAGCCAGCTCCTTGAGGGCCTGCTGGGGATCTTT;MAPQ=60;MATEID=6833945_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_45913001_45938001_102C;SPAN=4136;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:93 GQ:24.5 PL:[24.5, 0.0, 199.4] SR:15 DR:0 LR:-24.32 LO:32.44);ALT=T[chr19:45922356[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45924652	+	chr19	45926527	+	.	0	42	6833963_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6833963_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45913001_45938001_299C;SPAN=1875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:99 GQ:99 PL:[111.8, 0.0, 128.3] SR:42 DR:0 LR:-111.8 LO:111.9);ALT=C[chr19:45926527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45924696	+	chr19	45927049	+	.	23	0	6833965_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6833965_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45924696(+)-19:45927049(-)__19_45913001_45938001D;SPAN=2353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:81 GQ:54.2 PL:[54.2, 0.0, 140.0] SR:0 DR:23 LR:-53.98 LO:56.19);ALT=A[chr19:45927049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45974560	+	chr19	45975808	+	.	12	5	6834163_1	20.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6834163_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_45962001_45987001_353C;SPAN=1248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:96 GQ:20.3 PL:[20.3, 0.0, 211.7] SR:5 DR:12 LR:-20.21 LO:29.6);ALT=G[chr19:45975808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	45992827	+	chr19	45996417	+	.	9	0	6834055_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6834055_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:45992827(+)-19:45996417(-)__19_45986501_46011501D;SPAN=3590;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:88 GQ:5.9 PL:[5.9, 0.0, 207.2] SR:0 DR:9 LR:-5.868 LO:17.54);ALT=G[chr19:45996417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46010975	+	chr19	46020918	+	.	14	0	6834109_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6834109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46010975(+)-19:46020918(-)__19_45986501_46011501D;SPAN=9943;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:49 GQ:32.9 PL:[32.9, 0.0, 85.7] SR:0 DR:14 LR:-32.94 LO:34.25);ALT=G[chr19:46020918[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46191011	+	chr19	46195142	+	.	32	0	6834934_1	60.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=6834934_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46191011(+)-19:46195142(-)__19_46182501_46207501D;SPAN=4131;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:166 GQ:60.8 PL:[60.8, 0.0, 341.3] SR:0 DR:32 LR:-60.66 LO:71.95);ALT=A[chr19:46195142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46191852	+	chr19	46195141	+	.	139	0	6834939_1	99.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=6834939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46191852(+)-19:46195141(-)__19_46182501_46207501D;SPAN=3289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:139 DP:158 GQ:32.8 PL:[448.9, 32.8, 0.0] SR:0 DR:139 LR:-452.2 LO:452.2);ALT=G[chr19:46195141[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46658318	-	chr19	46749040	+	.	16	0	6836618_1	44.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6836618_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46658318(-)-19:46749040(-)__19_46746001_46771001D;SPAN=90722;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:29 GQ:25.1 PL:[44.9, 0.0, 25.1] SR:0 DR:16 LR:-45.25 LO:45.25);ALT=[chr19:46749040[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	46658486	+	chr19	46748743	-	.	19	0	6836619_1	52.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6836619_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:46658486(+)-19:46748743(+)__19_46746001_46771001D;SPAN=90257;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:37 GQ:36.2 PL:[52.7, 0.0, 36.2] SR:0 DR:19 LR:-52.84 LO:52.84);ALT=A]chr19:46748743];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	46850474	+	chr19	46857003	+	.	23	5	6836941_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6836941_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_46844001_46869001_189C;SPAN=6529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:78 GQ:61.4 PL:[61.4, 0.0, 127.4] SR:5 DR:23 LR:-61.39 LO:62.68);ALT=G[chr19:46857003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	46857249	+	chr19	46878860	+	.	3	8	6837202_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6837202_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_46868501_46893501_206C;SPAN=21611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:8 DR:3 LR:-20.5 LO:21.66);ALT=G[chr19:46878860[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47104695	+	chr19	47111451	+	CTGACCAGCTGACTGAGGAGCAGATTG	95	58	6837877_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CTGACCAGCTGACTGAGGAGCAGATTG;MAPQ=60;MATEID=6837877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47089001_47114001_115C;SPAN=6756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:117 DP:78 GQ:31.5 PL:[346.5, 31.5, 0.0] SR:58 DR:95 LR:-346.6 LO:346.6);ALT=G[chr19:47111451[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47342105	+	chr19	47354020	+	.	9	0	6839003_1	6.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=6839003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:47342105(+)-19:47354020(-)__19_47334001_47359001D;SPAN=11915;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:85 GQ:6.8 PL:[6.8, 0.0, 198.2] SR:0 DR:9 LR:-6.68 LO:17.69);ALT=C[chr19:47354020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47342837	+	chr19	47349250	+	.	3	99	6839006_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6839006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47334001_47359001_317C;SPAN=6413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:140 GQ:47.9 PL:[292.1, 0.0, 47.9] SR:99 DR:3 LR:-302.2 LO:302.2);ALT=T[chr19:47349250[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47342909	+	chr19	47354019	+	.	87	0	6839008_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6839008_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:47342909(+)-19:47354019(-)__19_47334001_47359001D;SPAN=11110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:87 DP:91 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:0 DR:87 LR:-267.4 LO:267.4);ALT=T[chr19:47354019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47349400	+	chr19	47354021	+	.	108	18	6839035_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6839035_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47334001_47359001_269C;SPAN=4621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:104 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:18 DR:108 LR:-340.0 LO:340.0);ALT=C[chr19:47354021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47549946	+	chr19	47551665	+	.	0	61	6839730_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6839730_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47530001_47555001_232C;SPAN=1719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:109 GQ:92.6 PL:[171.8, 0.0, 92.6] SR:61 DR:0 LR:-173.1 LO:173.1);ALT=G[chr19:47551665[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47634286	+	chr19	47646750	+	.	17	7	6839803_1	41.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6839803_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47628001_47653001_147C;SPAN=12464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:93 GQ:41 PL:[41.0, 0.0, 182.9] SR:7 DR:17 LR:-40.82 LO:46.04);ALT=G[chr19:47646750[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47646864	+	chr19	47653457	+	.	4	12	6839851_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=7;MATEID=6839851_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47628001_47653001_139C;SPAN=6593;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:34 GQ:37.1 PL:[43.7, 0.0, 37.1] SR:12 DR:4 LR:-43.62 LO:43.62);ALT=T[chr19:47653457[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47962798	+	chr19	47961550	+	.	27	0	6841074_1	64.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6841074_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:47961550(-)-19:47962798(+)__19_47946501_47971501D;SPAN=1248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:92 GQ:64.4 PL:[64.4, 0.0, 156.8] SR:0 DR:27 LR:-64.2 LO:66.43);ALT=]chr19:47962798]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	47987781	+	chr19	47996704	+	.	5	4	6841238_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6841238_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47971001_47996001_293C;SPAN=8923;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:34 GQ:10.7 PL:[10.7, 0.0, 70.1] SR:4 DR:5 LR:-10.59 LO:13.23);ALT=T[chr19:47996704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	47996859	+	chr19	47998283	+	.	0	4	6841118_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6841118_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47995501_48020501_303C;SPAN=1424;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:65 GQ:4.2 PL:[0.0, 4.2, 165.0] SR:4 DR:0 LR:4.406 LO:6.878);ALT=G[chr19:47998283[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48004007	+	chr19	48006680	+	.	0	21	6841138_1	42.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6841138_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47995501_48020501_129C;SPAN=2673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:98 GQ:42.8 PL:[42.8, 0.0, 194.6] SR:21 DR:0 LR:-42.77 LO:48.31);ALT=C[chr19:48006680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48004042	+	chr19	48018098	+	.	10	0	6841139_1	10.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6841139_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48004042(+)-19:48018098(-)__19_47995501_48020501D;SPAN=14056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:83 GQ:10.7 PL:[10.7, 0.0, 188.9] SR:0 DR:10 LR:-10.52 LO:20.25);ALT=G[chr19:48018098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48006760	+	chr19	48018100	+	.	0	33	6841147_1	80.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6841147_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_47995501_48020501_70C;SPAN=11340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:104 GQ:80.9 PL:[80.9, 0.0, 170.0] SR:33 DR:0 LR:-80.76 LO:82.56);ALT=C[chr19:48018100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48282049	+	chr19	48284544	+	.	16	0	6842461_1	23.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6842461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48282049(+)-19:48284544(-)__19_48265001_48290001D;SPAN=2495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:111 GQ:23 PL:[23.0, 0.0, 244.1] SR:0 DR:16 LR:-22.74 LO:33.74);ALT=C[chr19:48284544[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48282049	+	chr19	48284118	+	.	18	0	6842460_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6842460_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48282049(+)-19:48284118(-)__19_48265001_48290001D;SPAN=2069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:112 GQ:29.3 PL:[29.3, 0.0, 240.5] SR:0 DR:18 LR:-29.07 LO:38.89);ALT=C[chr19:48284118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48284645	+	chr19	48287545	+	.	5	21	6842475_1	60.0	.	DISC_MAPQ=46;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6842475_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48265001_48290001_300C;SPAN=2900;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:94 GQ:60.5 PL:[60.5, 0.0, 166.1] SR:21 DR:5 LR:-60.36 LO:63.17);ALT=G[chr19:48287545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48657227	+	chr19	48660271	+	.	3	10	6843571_1	11.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6843571_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48657001_48682001_99C;SPAN=3044;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:90 GQ:11.9 PL:[11.9, 0.0, 206.6] SR:10 DR:3 LR:-11.93 LO:22.35);ALT=G[chr19:48660271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48660401	+	chr19	48664629	+	.	2	7	6843580_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=6843580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48657001_48682001_42C;SPAN=4228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:7 DR:2 LR:-4.192 LO:15.42);ALT=G[chr19:48664629[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48665608	+	chr19	48673497	+	ATGATACTTCGCTGCATGTTGGCGTCAGAATTCTCCCTTCCTGTCCAGCACTTTTCTTCGTCTGTCAGCTGCT	9	14	6843601_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=ATGATACTTCGCTGCATGTTGGCGTCAGAATTCTCCCTTCCTGTCCAGCACTTTTCTTCGTCTGTCAGCTGCT;MAPQ=60;MATEID=6843601_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_48657001_48682001_211C;SPAN=7889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:60 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:14 DR:9 LR:-43.16 LO:44.49);ALT=C[chr19:48673497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48668882	+	chr19	48673497	+	.	6	5	6843611_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCT;MAPQ=60;MATEID=6843611_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_48657001_48682001_211C;SPAN=4615;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:62 GQ:6.5 PL:[6.5, 0.0, 141.8] SR:5 DR:6 LR:-6.31 LO:13.96);ALT=T[chr19:48673497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48741790	+	chr19	48744218	+	.	0	18	6843847_1	36.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6843847_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48730501_48755501_11C;SPAN=2428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:84 GQ:36.8 PL:[36.8, 0.0, 165.5] SR:18 DR:0 LR:-36.66 LO:41.41);ALT=C[chr19:48744218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48741835	+	chr19	48753006	+	.	8	0	6843848_1	2.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6843848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48741835(+)-19:48753006(-)__19_48730501_48755501D;SPAN=11171;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:89 GQ:2.3 PL:[2.3, 0.0, 213.5] SR:0 DR:8 LR:-2.296 LO:15.12);ALT=C[chr19:48753006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48744320	+	chr19	48752779	+	.	0	8	6843857_1	5.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6843857_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48730501_48755501_42C;SPAN=8459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:77 GQ:5.6 PL:[5.6, 0.0, 180.5] SR:8 DR:0 LR:-5.547 LO:15.65);ALT=C[chr19:48752779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48744363	+	chr19	48753009	+	.	8	0	6843858_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6843858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48744363(+)-19:48753009(-)__19_48730501_48755501D;SPAN=8646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=A[chr19:48753009[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48828867	+	chr19	48830777	+	.	26	13	6844667_1	63.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6844667_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48828501_48853501_16C;SPAN=1910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:194 GQ:63.1 PL:[63.1, 0.0, 406.4] SR:13 DR:26 LR:-62.98 LO:77.57);ALT=G[chr19:48830777[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48828868	+	chr19	48830086	+	.	43	72	6844163_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6844163_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48804001_48829001_26C;SPAN=1218;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:115 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:72 DR:43 LR:-340.0 LO:340.0);ALT=G[chr19:48830086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48828868	+	chr19	48832608	+	.	7	3	6844670_1	0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6844670_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48828501_48853501_118C;SPAN=3740;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:191 GQ:18.4 PL:[0.0, 18.4, 498.4] SR:3 DR:7 LR:18.74 LO:16.48);ALT=G[chr19:48832608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48830881	+	chr19	48832608	+	.	12	67	6844677_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6844677_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48828501_48853501_356C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:76 DP:138 GQ:99 PL:[213.5, 0.0, 121.1] SR:67 DR:12 LR:-214.8 LO:214.8);ALT=G[chr19:48832608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48830924	+	chr19	48833556	+	.	8	0	6844678_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6844678_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:48830924(+)-19:48833556(-)__19_48828501_48853501D;SPAN=2632;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:138 GQ:10.8 PL:[0.0, 10.8, 356.4] SR:0 DR:8 LR:10.98 LO:13.54);ALT=A[chr19:48833556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	48887741	+	chr19	48892810	+	.	3	3	6845190_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6845190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_48877501_48902501_278C;SPAN=5069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:85 GQ:3 PL:[0.0, 3.0, 211.2] SR:3 DR:3 LR:3.223 LO:10.69);ALT=T[chr19:48892810[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49120720	+	chr19	49122396	+	.	26	0	6846698_1	49.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6846698_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49120720(+)-19:49122396(-)__19_49098001_49123001D;SPAN=1676;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:134 GQ:49.7 PL:[49.7, 0.0, 274.1] SR:0 DR:26 LR:-49.52 LO:58.54);ALT=G[chr19:49122396[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49121135	+	chr19	49122397	+	.	8	40	6846699_1	97.0	.	DISC_MAPQ=24;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6846699_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49098001_49123001_370C;SPAN=1262;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:200 GQ:97.6 PL:[97.6, 0.0, 388.1] SR:40 DR:8 LR:-97.66 LO:107.4);ALT=C[chr19:49122397[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49310010	+	chr19	49314240	+	.	15	0	6846432_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6846432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49310010(+)-19:49314240(-)__19_49294001_49319001D;SPAN=4230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:89 GQ:25.4 PL:[25.4, 0.0, 190.4] SR:0 DR:15 LR:-25.4 LO:32.75);ALT=C[chr19:49314240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49404124	+	chr19	49407602	+	.	44	0	6847145_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847145_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49404124(+)-19:49407602(-)__19_49392001_49417001D;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:130 GQ:99 PL:[110.0, 0.0, 205.7] SR:0 DR:44 LR:-110.0 LO:111.6);ALT=T[chr19:49407602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49404124	+	chr19	49409006	+	.	20	0	6847146_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847146_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49404124(+)-19:49409006(-)__19_49392001_49417001D;SPAN=4882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:111 GQ:36.2 PL:[36.2, 0.0, 230.9] SR:0 DR:20 LR:-35.95 LO:44.31);ALT=T[chr19:49409006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49407711	+	chr19	49409008	+	.	3	23	6847157_1	56.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6847157_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49392001_49417001_132C;SPAN=1297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:107 GQ:56.9 PL:[56.9, 0.0, 202.1] SR:23 DR:3 LR:-56.84 LO:61.44);ALT=G[chr19:49409008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49414510	+	chr19	49416267	+	.	6	8	6847182_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6847182_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49392001_49417001_181C;SPAN=1757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:8 DR:6 LR:-16.31 LO:25.12);ALT=G[chr19:49416267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49416474	+	chr19	49421981	+	.	10	0	6847209_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49416474(+)-19:49421981(-)__19_49416501_49441501D;SPAN=5507;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:0 DR:10 LR:-17.3 LO:21.94);ALT=C[chr19:49421981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49416821	+	chr19	49422285	+	ATATCAACAGTGATGGTGTCCTGGATGAGCAGGAGCTGGAGGCACTCTTCACCAAGG	0	19	6847212_1	43.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATATCAACAGTGATGGTGTCCTGGATGAGCAGGAGCTGGAGGCACTCTTCACCAAGG;MAPQ=60;MATEID=6847212_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_49416501_49441501_259C;SPAN=5464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:73 GQ:43.1 PL:[43.1, 0.0, 132.2] SR:19 DR:0 LR:-42.94 LO:45.56);ALT=G[chr19:49422285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49459091	+	chr19	49464065	+	ATGATTGCCGCCGTGGACACAGACTCCCCCCGAGAGGTCTTTTTCCGAGTGGCAGCTGACATGTTTTCTGACGGCAACTTCAACTGGGGCCGGGTTGTCGCCCTTTTCTACTTTGCCAGCAAACTGGTGCTCA	0	90	6847387_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATGATTGCCGCCGTGGACACAGACTCCCCCCGAGAGGTCTTTTTCCGAGTGGCAGCTGACATGTTTTCTGACGGCAACTTCAACTGGGGCCGGGTTGTCGCCCTTTTCTACTTTGCCAGCAAACTGGTGCTCA;MAPQ=60;MATEID=6847387_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_49441001_49466001_377C;SPAN=4974;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:113 GQ:5.9 PL:[266.6, 0.0, 5.9] SR:90 DR:0 LR:-281.3 LO:281.3);ALT=G[chr19:49464065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49497233	+	chr19	49507530	+	.	24	0	6847852_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847852_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49497233(+)-19:49507530(-)__19_49490001_49515001D;SPAN=10297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:79 GQ:57.8 PL:[57.8, 0.0, 133.7] SR:0 DR:24 LR:-57.82 LO:59.49);ALT=G[chr19:49507530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49502659	+	chr19	49507530	+	.	18	0	6847878_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6847878_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49502659(+)-19:49507530(-)__19_49490001_49515001D;SPAN=4871;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:88 GQ:35.6 PL:[35.6, 0.0, 177.5] SR:0 DR:18 LR:-35.58 LO:40.99);ALT=T[chr19:49507530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49507676	+	chr19	49510274	+	.	5	17	6847895_1	42.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6847895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49490001_49515001_317C;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:88 GQ:42.2 PL:[42.2, 0.0, 170.9] SR:17 DR:5 LR:-42.18 LO:46.59);ALT=G[chr19:49510274[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49514567	+	chr19	49517740	+	.	3	3	6847918_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6847918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49490001_49515001_98C;SPAN=3173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:30 GQ:11.6 PL:[11.6, 0.0, 61.1] SR:3 DR:3 LR:-11.68 LO:13.6);ALT=G[chr19:49517740[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49607993	+	chr19	49610880	+	.	5	13	6848092_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6848092_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_49588001_49613001_250C;SPAN=2887;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:105 GQ:24.5 PL:[24.5, 0.0, 229.1] SR:13 DR:5 LR:-24.37 LO:34.16);ALT=G[chr19:49610880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49670800	+	chr19	49669732	+	.	27	0	6848644_1	68.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=6848644_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49669732(-)-19:49670800(+)__19_49661501_49686501D;SPAN=1068;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:77 GQ:68.3 PL:[68.3, 0.0, 117.8] SR:0 DR:27 LR:-68.27 LO:69.01);ALT=]chr19:49670800]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	49839044	+	chr19	49840165	+	.	46	113	6849161_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6849161_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_49833001_49858001_283C;SPAN=1121;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:129 DP:184 GQ:69.1 PL:[376.1, 0.0, 69.1] SR:113 DR:46 LR:-387.8 LO:387.8);ALT=G[chr19:49840165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49841286	+	chr19	49843506	+	CTGCGCTGCTGCGGCTGGCACTACCCGCAGGACTGGTTCCAAGTCCTCATCCTGAGAGGTAACGGGTCGGAGGCGCACCGCGTGCCCTGCTCCTGCTACAACTTGTCGGCGACCAACGACTCCACAATCCTAGATAAGGTGATCTTGCCCCAGCTCAGCAGGCTTGGACACCTGGCGCGGTCCAGACACAGTGCAGACATCTGCGCTGTCCCTGCAGAGAGCCACATCTACCGCGAGGGCTGCGCGCAGGGCCTCCAGAAGTGGCTGCACAACAACCTTATTTCCATAGTGGGCATTTGCCTGGGCGTCGGCCTACTCG	0	36	6849172_1	89.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTGCGCTGCTGCGGCTGGCACTACCCGCAGGACTGGTTCCAAGTCCTCATCCTGAGAGGTAACGGGTCGGAGGCGCACCGCGTGCCCTGCTCCTGCTACAACTTGTCGGCGACCAACGACTCCACAATCCTAGATAAGGTGATCTTGCCCCAGCTCAGCAGGCTTGGACACCTGGCGCGGTCCAGACACAGTGCAGACATCTGCGCTGTCCCTGCAGAGAGCCACATCTACCGCGAGGGCTGCGCGCAGGGCCTCCAGAAGTGGCTGCACAACAACCTTATTTCCATAGTGGGCATTTGCCTGGGCGTCGGCCTACTCG;MAPQ=60;MATEID=6849172_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_19_49833001_49858001_15C;SPAN=2220;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:108 GQ:89.6 PL:[89.6, 0.0, 172.1] SR:36 DR:0 LR:-89.58 LO:91.02);ALT=G[chr19:49843506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49956679	+	chr19	49961742	+	.	13	7	6849250_1	8.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6849250_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CTGGCTGG;SCTG=c_19_49955501_49980501_240C;SPAN=5063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:80 GQ:8.5 PL:[8.5, 0.0, 92.3] SR:7 DR:13 LR:-8.326 LO:14.18);ALT=G[chr19:49961742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49956679	+	chr19	49962214	+	CCTGGCTGGACACCCAGGACCGGTGCTTGGGCCACTATGTGAATGGGAAGTGGTTAAAGCCTGAACACAGAAATTCAGTGCCTTGCCAGGATCCCATCA	5	18	6849251_1	39.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CCTGGCTGGACACCCAGGACCGGTGCTTGGGCCACTATGTGAATGGGAAGTGGTTAAAGCCTGAACACAGAAATTCAGTGCCTTGCCAGGATCCCATCA;MAPQ=60;MATEID=6849251_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_49955501_49980501_240C;SPAN=5535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:87 GQ:39.2 PL:[39.2, 0.0, 171.2] SR:18 DR:5 LR:-39.15 LO:43.89);ALT=G[chr19:49962214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	49999773	+	chr19	50001172	+	.	18	0	6849514_1	7.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6849514_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:49999773(+)-19:50001172(-)__19_49980001_50005001D;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:190 GQ:7.9 PL:[7.9, 0.0, 453.5] SR:0 DR:18 LR:-7.942 LO:34.46);ALT=C[chr19:50001172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50000886	+	chr19	50002765	+	.	29	0	6849518_1	18.0	.	DISC_MAPQ=23;EVDNC=DSCRD;IMPRECISE;MAPQ=23;MATEID=6849518_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50000886(+)-19:50002765(-)__19_49980001_50005001D;SPAN=1879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:286 GQ:18.4 PL:[18.4, 0.0, 675.2] SR:0 DR:29 LR:-18.24 LO:56.42);ALT=A[chr19:50002765[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50060508	+	chr19	50062153	+	.	0	15	6849757_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6849757_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50053501_50078501_167C;SPAN=1645;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:82 GQ:27.5 PL:[27.5, 0.0, 169.4] SR:15 DR:0 LR:-27.3 LO:33.34);ALT=T[chr19:50062153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50060542	+	chr19	50083770	+	.	10	0	6849758_1	24.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6849758_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50060542(+)-19:50083770(-)__19_50053501_50078501D;SPAN=23228;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:33 GQ:24.2 PL:[24.2, 0.0, 53.9] SR:0 DR:10 LR:-24.07 LO:24.77);ALT=G[chr19:50083770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50062283	+	chr19	50083770	+	.	24	0	6849766_1	68.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6849766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50062283(+)-19:50083770(-)__19_50053501_50078501D;SPAN=21487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:41 GQ:28.7 PL:[68.3, 0.0, 28.7] SR:0 DR:24 LR:-68.85 LO:68.85);ALT=C[chr19:50083770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50063331	+	chr19	50083770	+	.	24	0	6849775_1	68.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6849775_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50063331(+)-19:50083770(-)__19_50053501_50078501D;SPAN=20439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:41 GQ:28.7 PL:[68.3, 0.0, 28.7] SR:0 DR:24 LR:-68.85 LO:68.85);ALT=G[chr19:50083770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50063988	+	chr19	50083770	+	.	10	0	6849778_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6849778_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50063988(+)-19:50083770(-)__19_50053501_50078501D;SPAN=19782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.19 LO:22.57);ALT=G[chr19:50083770[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50173746	+	chr19	50176954	+	.	0	10	6850000_1	20.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6850000_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50151501_50176501_139C;SPAN=3208;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:10 DR:0 LR:-20.55 LO:23.07);ALT=G[chr19:50176954[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50180576	+	chr19	50183742	+	.	30	5	6850108_1	77.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=20;MATEID=6850108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50176001_50201001_75C;SPAN=3166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:116 GQ:77.6 PL:[77.6, 0.0, 203.0] SR:5 DR:30 LR:-77.51 LO:80.66);ALT=G[chr19:50183742[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50180613	+	chr19	50185162	+	.	53	0	6850109_1	99.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6850109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50180613(+)-19:50185162(-)__19_50176001_50201001D;SPAN=4549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:69 GQ:11 PL:[156.2, 0.0, 11.0] SR:0 DR:53 LR:-163.7 LO:163.7);ALT=T[chr19:50185162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50183846	+	chr19	50185165	+	.	0	37	6850120_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6850120_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50176001_50201001_109C;SPAN=1319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:84 GQ:99 PL:[99.5, 0.0, 102.8] SR:37 DR:0 LR:-99.38 LO:99.39);ALT=G[chr19:50185165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50189983	+	chr19	50191419	+	.	2	28	6850145_1	75.0	.	DISC_MAPQ=12;EVDNC=ASDIS;MAPQ=31;MATEID=6850145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50176001_50201001_248C;SPAN=1436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:88 GQ:75.2 PL:[75.2, 0.0, 137.9] SR:28 DR:2 LR:-75.19 LO:76.21);ALT=C[chr19:50191419[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50197790	+	chr19	50198936	-	.	10	0	6850168_1	8.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=6850168_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50197790(+)-19:50198936(+)__19_50176001_50201001D;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:89 GQ:8.9 PL:[8.9, 0.0, 206.9] SR:0 DR:10 LR:-8.898 LO:19.93);ALT=G]chr19:50198936];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	50432659	+	chr19	50433989	+	.	0	8	6851478_1	3.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=6851478_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50421001_50446001_69C;SPAN=1330;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:86 GQ:3.2 PL:[3.2, 0.0, 204.5] SR:8 DR:0 LR:-3.109 LO:15.25);ALT=T[chr19:50433989[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50511085	+	chr19	50512492	+	.	0	5	6851110_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6851110_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50494501_50519501_145C;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:80 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:5 DR:0 LR:5.169 LO:8.632);ALT=T[chr19:50512492[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50512644	+	chr19	50523842	+	TGGAAGGATGACACATGTGGATTGACAAAGGTCTGGGACCCTACATGCTCCTCTACAGGCAAAGAATTTCCACAGTAGGGGCAGAATTTGAATGCCGCTTGGATACTTTTGCCACAGTCTGGACAGAAGGAGATCATG	9	12	6851349_1	47.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TGGAAGGATGACACATGTGGATTGACAAAGGTCTGGGACCCTACATGCTCCTCTACAGGCAAAGAATTTCCACAGTAGGGGCAGAATTTGAATGCCGCTTGGATACTTTTGCCACAGTCTGGACAGAAGGAGATCATG;MAPQ=60;MATEID=6851349_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_50519001_50544001_7C;SPAN=11198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:33 GQ:30.8 PL:[47.3, 0.0, 30.8] SR:12 DR:9 LR:-47.31 LO:47.31);ALT=T[chr19:50523842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50519422	+	chr19	50523842	+	.	4	5	6851351_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6851351_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_50519001_50544001_7C;SPAN=4420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:5 DR:4 LR:-10.2 LO:18.38);ALT=T[chr19:50523842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50519461	+	chr19	50528599	+	.	8	0	6851352_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6851352_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50519461(+)-19:50528599(-)__19_50519001_50544001D;SPAN=9138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:73 GQ:6.8 PL:[6.8, 0.0, 168.5] SR:0 DR:8 LR:-6.631 LO:15.85);ALT=G[chr19:50528599[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50840933	+	chr19	50847929	+	.	124	15	6852589_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6852589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_50837501_50862501_102C;SPAN=6996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:99 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:15 DR:124 LR:-382.9 LO:382.9);ALT=C[chr19:50847929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50879834	+	chr19	50880842	+	GCAACAGGAGTAGTTCACTCCGCGAGAGGCCGTCCACGAGACCCCCGCGCGCAGCCATGAGCCCCGCCCCCCGCTGTTGCTTGGAGAGGGGCGGGACCTGGAGAG	24	32	6852527_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=GCAACAGGAGTAGTTCACTCCGCGAGAGGCCGTCCACGAGACCCCCGCGCGCAGCCATGAGCCCCGCCCCCCGCTGTTGCTTGGAGAGGGGCGGGACCTGGAGAG;MAPQ=60;MATEID=6852527_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_50862001_50887001_260C;SPAN=1008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:98 GQ:99 PL:[115.4, 0.0, 122.0] SR:32 DR:24 LR:-115.4 LO:115.4);ALT=G[chr19:50880842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50887689	+	chr19	50902104	+	.	10	0	6852747_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6852747_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:50887689(+)-19:50902104(-)__19_50886501_50911501D;SPAN=14415;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:98 GQ:6.5 PL:[6.5, 0.0, 230.9] SR:0 DR:10 LR:-6.459 LO:19.48);ALT=G[chr19:50902104[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	50979916	+	chr19	50982213	+	CTGGGGCGGAAGGTCGAGAGGGCGAGGCCTGTGGCACGGTGGGGCTGCTGCTGGAGCACTCATTTGAGATC	41	67	6852878_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTGGGGCGGAAGGTCGAGAGGGCGAGGCCTGTGGCACGGTGGGGCTGCTGCTGGAGCACTCATTTGAGATC;MAPQ=60;MATEID=6852878_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_50960001_50985001_164C;SPAN=2297;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:102 GQ:17.4 PL:[280.5, 17.4, 0.0] SR:67 DR:41 LR:-283.6 LO:283.6);ALT=G[chr19:50982213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51009831	+	chr19	51013542	+	.	0	7	6852987_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6852987_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51009001_51034001_193C;SPAN=3711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:94 GQ:2.1 PL:[0.0, 2.1, 231.0] SR:7 DR:0 LR:2.36 LO:12.64);ALT=T[chr19:51013542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51010958	+	chr19	51013541	+	.	0	23	6852990_1	51.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6852990_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51009001_51034001_307C;SPAN=2583;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:91 GQ:51.5 PL:[51.5, 0.0, 167.0] SR:23 DR:0 LR:-51.27 LO:54.81);ALT=T[chr19:51013541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51011004	+	chr19	51014347	+	.	21	0	6852991_1	49.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6852991_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51011004(+)-19:51014347(-)__19_51009001_51034001D;SPAN=3343;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:75 GQ:49.1 PL:[49.1, 0.0, 131.6] SR:0 DR:21 LR:-49.0 LO:51.15);ALT=C[chr19:51014347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51302230	+	chr19	51307824	+	.	9	0	6855160_1	18.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6855160_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51302230(+)-19:51307824(-)__19_51278501_51303501D;SPAN=5594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:40 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:0 DR:9 LR:-18.87 LO:20.92);ALT=A[chr19:51307824[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51302260	+	chr19	51305475	+	.	54	0	6855161_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6855161_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51302260(+)-19:51305475(-)__19_51278501_51303501D;SPAN=3215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:41 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:54 LR:-158.4 LO:158.4);ALT=C[chr19:51305475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51406777	+	chr19	51408332	+	.	24	11	6855780_1	94.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=GAGTAGCTGGGATTACAGGCAC;MAPQ=60;MATEID=6855780_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_51401001_51426001_5C;SPAN=1555;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:55 GQ:38 PL:[94.1, 0.0, 38.0] SR:11 DR:24 LR:-95.25 LO:95.25);ALT=C[chr19:51408332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51848636	+	chr19	51850154	+	.	6	75	6857069_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6857069_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51842001_51867001_218C;SPAN=1518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:119 GQ:60.2 PL:[228.5, 0.0, 60.2] SR:75 DR:6 LR:-234.0 LO:234.0);ALT=C[chr19:51850154[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51853648	+	chr19	51856385	+	.	5	13	6857089_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=6857089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51842001_51867001_159C;SPAN=2737;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:93 GQ:31.1 PL:[31.1, 0.0, 192.8] SR:13 DR:5 LR:-30.92 LO:37.78);ALT=G[chr19:51856385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51856597	+	chr19	51869525	+	.	54	0	6857157_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6857157_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:51856597(+)-19:51869525(-)__19_51866501_51891501D;SPAN=12928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:54 DP:56 GQ:15 PL:[165.0, 15.0, 0.0] SR:0 DR:54 LR:-165.0 LO:165.0);ALT=A[chr19:51869525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	51857564	+	chr19	51869524	+	.	143	30	6857158_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6857158_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_51866501_51891501_197C;SPAN=11960;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:145 DP:55 GQ:39.1 PL:[429.1, 39.1, 0.0] SR:30 DR:143 LR:-429.1 LO:429.1);ALT=T[chr19:51869524[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52175937	+	chr19	52177514	+	.	60	30	6857843_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=TAATTTTC;MAPQ=60;MATEID=6857843_2;MATENM=5;NM=0;NUMPARTS=2;SCTG=c_19_52160501_52185501_270C;SPAN=1577;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:83 DP:31 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:30 DR:60 LR:-244.3 LO:244.3);ALT=C[chr19:52177514[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52693413	+	chr19	52714509	+	.	8	0	6859281_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6859281_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52693413(+)-19:52714509(-)__19_52699501_52724501D;SPAN=21096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:0 DR:8 LR:-7.985 LO:16.11);ALT=A[chr19:52714509[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52693419	+	chr19	52709211	+	.	50	0	6859425_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6859425_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52693419(+)-19:52709211(-)__19_52675001_52700001D;SPAN=15792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:43 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:0 DR:50 LR:-148.5 LO:148.5);ALT=G[chr19:52709211[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52693427	+	chr19	52705195	+	.	48	32	6859426_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6859426_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52675001_52700001_321C;SPAN=11768;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:39 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:32 DR:48 LR:-181.5 LO:181.5);ALT=G[chr19:52705195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52705287	+	chr19	52709212	+	.	0	60	6859298_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACAG;MAPQ=60;MATEID=6859298_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52699501_52724501_142C;SPAN=3925;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:123 GQ:99 PL:[164.9, 0.0, 131.9] SR:60 DR:0 LR:-164.9 LO:164.9);ALT=G[chr19:52709212[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52709316	+	chr19	52714512	+	.	3	24	6859306_1	54.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6859306_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_52699501_52724501_335C;SPAN=5196;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:128 GQ:54.5 PL:[54.5, 0.0, 255.8] SR:24 DR:3 LR:-54.45 LO:61.9);ALT=G[chr19:52714512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52725494	+	chr19	52728967	+	.	2	5	6859205_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6859205_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52724001_52749001_106C;SPAN=3473;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:84 GQ:0.5 PL:[0.5, 0.0, 201.8] SR:5 DR:2 LR:-0.3493 LO:12.99);ALT=G[chr19:52728967[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52800521	+	chr19	52817403	+	.	17	0	6859686_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6859686_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52800521(+)-19:52817403(-)__19_52797501_52822501D;SPAN=16882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:51 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.3 LO:42.98);ALT=C[chr19:52817403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52803738	+	chr19	52817404	+	.	0	8	6859693_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6859693_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52797501_52822501_172C;SPAN=13666;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:8 DR:0 LR:-7.443 LO:16.0);ALT=G[chr19:52817404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52860681	+	chr19	52861707	-	.	9	0	6859797_1	6.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6859797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52860681(+)-19:52861707(+)__19_52846501_52871501D;SPAN=1026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:86 GQ:6.5 PL:[6.5, 0.0, 201.2] SR:0 DR:9 LR:-6.41 LO:17.64);ALT=G]chr19:52861707];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	52873281	+	chr19	52877550	+	.	10	0	6860433_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6860433_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:52873281(+)-19:52877550(-)__19_52871001_52896001D;SPAN=4269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:106 GQ:4.4 PL:[4.4, 0.0, 251.9] SR:0 DR:10 LR:-4.292 LO:19.12);ALT=C[chr19:52877550[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	52876491	+	chr19	52877551	+	.	0	10	6860446_1	11.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6860446_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_52871001_52896001_142C;SPAN=1060;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:80 GQ:11.3 PL:[11.3, 0.0, 182.9] SR:10 DR:0 LR:-11.34 LO:20.42);ALT=G[chr19:52877551[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53096022	+	chr19	53097609	+	.	94	28	6860645_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CTAATTTTGTATTTTT;MAPQ=60;MATEID=6860645_2;MATENM=2;NM=5;NUMPARTS=2;SCTG=c_19_53091501_53116501_68C;SPAN=1587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:25 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:28 DR:94 LR:-320.2 LO:320.2);ALT=T[chr19:53097609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53418276	+	chr19	53391273	+	.	11	0	6862106_1	25.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=6862106_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53391273(-)-19:53418276(+)__19_53410001_53435001D;SPAN=27003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:39 GQ:25.7 PL:[25.7, 0.0, 68.6] SR:0 DR:11 LR:-25.75 LO:26.84);ALT=]chr19:53418276]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	53422211	+	chr19	53424207	+	.	66	20	6862139_1	84.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AAAAAAAAAAAAAA;MAPQ=60;MATEID=6862139_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_19_53410001_53435001_234C;SPAN=1996;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:78 DP:640 GQ:84.1 PL:[84.1, 0.0, 1470.0] SR:20 DR:66 LR:-84.09 LO:158.4);ALT=A[chr19:53424207[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	53788594	+	chr19	53801879	-	.	12	0	6862513_1	21.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=6862513_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53788594(+)-19:53801879(+)__19_53777501_53802501D;SPAN=13285;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:68 GQ:21.2 PL:[21.2, 0.0, 143.3] SR:0 DR:12 LR:-21.19 LO:26.47);ALT=G]chr19:53801879];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr19	53983536	+	chr19	53946077	+	.	9	0	6863475_1	17.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6863475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:53946077(-)-19:53983536(+)__19_53924501_53949501D;SPAN=37459;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=]chr19:53983536]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54263915	+	chr19	54232687	+	GCAGGATAGACCACAGACTAGGATGTAAAAGCTCCTCAATAAAATTTGAATCTAAATACACAAGTACAGG	12	84	6864913_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;INSERTION=GCAGGATAGACCACAGACTAGGATGTAAAAGCTCCTCAATAAAATTTGAATCTAAATACACAAGTACAGG;MAPQ=60;MATEID=6864913_2;MATENM=9;NM=0;NUMPARTS=2;SCTG=c_19_54243001_54268001_203C;SPAN=31228;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:55 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:84 DR:12 LR:-267.4 LO:267.4);ALT=]chr19:54263915]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54251538	+	chr19	54232719	+	.	12	0	6864914_1	28.0	.	DISC_MAPQ=41;EVDNC=DSCRD;IMPRECISE;MAPQ=41;MATEID=6864914_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54232719(-)-19:54251538(+)__19_54243001_54268001D;SPAN=18819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:43 GQ:28.1 PL:[28.1, 0.0, 74.3] SR:0 DR:12 LR:-27.96 LO:29.21);ALT=]chr19:54251538]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54371200	+	chr19	54373006	+	.	8	4	6865217_1	3.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AGGTG;MAPQ=60;MATEID=6865217_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54365501_54390501_220C;SPAN=1806;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:122 GQ:3.5 PL:[3.5, 0.0, 290.6] SR:4 DR:8 LR:-3.258 LO:20.81);ALT=G[chr19:54373006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54371200	+	chr19	54376781	+	CTCTTACAGCCTGTTCCAAGTGTGGCTTAATCCGTCTCCACCACCAGATCTTTCTCCGTGGATTCCTCTGCTAAGACCGCT	114	46	6865218_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CTCTTACAGCCTGTTCCAAGTGTGGCTTAATCCGTCTCCACCACCAGATCTTTCTCCGTGGATTCCTCTGCTAAGACCGCT;MAPQ=60;MATEID=6865218_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54365501_54390501_220C;SPAN=5581;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:138 DP:157 GQ:32.5 PL:[445.6, 32.5, 0.0] SR:46 DR:114 LR:-448.7 LO:448.7);ALT=G[chr19:54376781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54373092	+	chr19	54376781	+	.	44	41	6865225_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6865225_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54365501_54390501_220C;SPAN=3689;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:105 GQ:11.3 PL:[242.3, 0.0, 11.3] SR:41 DR:44 LR:-254.6 LO:254.6);ALT=G[chr19:54376781[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54428719	+	chr19	54426619	+	.	41	0	6865939_1	99.0	.	DISC_MAPQ=20;EVDNC=DSCRD;IMPRECISE;MAPQ=20;MATEID=6865939_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54426619(-)-19:54428719(+)__19_54414501_54439501D;SPAN=2100;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:130 GQ:99 PL:[100.1, 0.0, 215.6] SR:0 DR:41 LR:-100.1 LO:102.4);ALT=]chr19:54428719]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr19	54600512	+	chr19	54604044	+	.	24	0	6866500_1	57.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6866500_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54600512(+)-19:54604044(-)__19_54586001_54611001D;SPAN=3532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:79 GQ:57.8 PL:[57.8, 0.0, 133.7] SR:0 DR:24 LR:-57.82 LO:59.49);ALT=A[chr19:54604044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54602972	+	chr19	54604045	+	.	9	0	6866506_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6866506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54602972(+)-19:54604045(-)__19_54586001_54611001D;SPAN=1073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:80 GQ:8 PL:[8.0, 0.0, 186.2] SR:0 DR:9 LR:-8.035 LO:17.94);ALT=A[chr19:54604045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54606496	+	chr19	54609240	+	.	37	49	6866525_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6866525_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54586001_54611001_271C;SPAN=2744;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:75 DP:132 GQ:99 PL:[212.0, 0.0, 106.4] SR:49 DR:37 LR:-213.6 LO:213.6);ALT=G[chr19:54609240[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54606545	+	chr19	54610112	+	.	64	0	6866526_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6866526_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54606545(+)-19:54610112(-)__19_54586001_54611001D;SPAN=3567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:134 GQ:99 PL:[175.1, 0.0, 148.7] SR:0 DR:64 LR:-175.1 LO:175.1);ALT=C[chr19:54610112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54611704	+	chr19	54613432	+	.	0	12	6866166_1	14.0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6866166_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54610501_54635501_257C;SPAN=1728;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:92 GQ:14.9 PL:[14.9, 0.0, 206.3] SR:12 DR:0 LR:-14.69 LO:24.74);ALT=T[chr19:54613432[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54611752	+	chr19	54617846	+	.	14	0	6866167_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6866167_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54611752(+)-19:54617846(-)__19_54610501_54635501D;SPAN=6094;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:90 GQ:21.8 PL:[21.8, 0.0, 196.7] SR:0 DR:14 LR:-21.83 LO:30.03);ALT=G[chr19:54617846[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54613506	+	chr19	54617820	+	.	0	7	6866176_1	0	.	EVDNC=ASSMB;HOMSEQ=ACCT;MAPQ=60;MATEID=6866176_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54610501_54635501_383C;SPAN=4314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:96 GQ:2.7 PL:[0.0, 2.7, 237.6] SR:7 DR:0 LR:2.902 LO:12.57);ALT=T[chr19:54617820[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54621835	+	chr19	54625237	+	TTTGCTGAGATTATGATGAAGATTGAGGAGTATATCAGCAAGCAAGCCAAAGCTTCAGA	0	18	6866213_1	36.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTTGCTGAGATTATGATGAAGATTGAGGAGTATATCAGCAAGCAAGCCAAAGCTTCAGA;MAPQ=60;MATEID=6866213_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54610501_54635501_295C;SPAN=3402;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:86 GQ:36.2 PL:[36.2, 0.0, 171.5] SR:18 DR:0 LR:-36.12 LO:41.2);ALT=G[chr19:54625237[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54629995	+	chr19	54631446	+	.	0	6	6866249_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGTG;MAPQ=60;MATEID=6866249_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54610501_54635501_207C;SPAN=1451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:75 GQ:0.3 PL:[0.0, 0.3, 181.5] SR:6 DR:0 LR:0.5133 LO:11.02);ALT=G[chr19:54631446[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54678126	+	chr19	54682481	+	.	6	8	6866416_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6866416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54659501_54684501_113C;SPAN=4355;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:84 GQ:13.7 PL:[13.7, 0.0, 188.6] SR:8 DR:6 LR:-13.55 LO:22.7);ALT=C[chr19:54682481[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54682661	+	chr19	54684490	+	.	8	4	6866620_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6866620_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54684001_54709001_321C;SPAN=1829;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:34 GQ:27.2 PL:[27.2, 0.0, 53.6] SR:4 DR:8 LR:-27.1 LO:27.63);ALT=G[chr19:54684490[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54684854	+	chr19	54691043	+	CATGATTCCCACGTAGCAGTAGCTGTAGCTGAGTGTCTCCATCAGGGAGGGCACGTCGGGCAGCAGCCCCAGGGTGGGCCCCTTGCTGAAGCCTGAGGCCATTTCCTTCCTCTGGGCCAGATGCAGGTCCTGGACTTCACTGGCCAGGCTCACCAG	2	20	6866625_1	43.0	.	DISC_MAPQ=45;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CATGATTCCCACGTAGCAGTAGCTGTAGCTGAGTGTCTCCATCAGGGAGGGCACGTCGGGCAGCAGCCCCAGGGTGGGCCCCTTGCTGAAGCCTGAGGCCATTTCCTTCCTCTGGGCCAGATGCAGGTCCTGGACTTCACTGGCCAGGCTCACCAG;MAPQ=60;MATEID=6866625_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54684001_54709001_179C;SPAN=6189;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:96 GQ:43.4 PL:[43.4, 0.0, 188.6] SR:20 DR:2 LR:-43.31 LO:48.52);ALT=T[chr19:54691043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54684854	+	chr19	54687403	+	.	4	6	6866624_1	6.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CCTGT;MAPQ=60;MATEID=6866624_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54684001_54709001_179C;SPAN=2549;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:86 GQ:6.5 PL:[6.5, 0.0, 201.2] SR:6 DR:4 LR:-6.41 LO:17.64);ALT=T[chr19:54687403[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54687565	+	chr19	54691043	+	.	4	15	6866634_1	25.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6866634_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_54684001_54709001_179C;SPAN=3478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:100 GQ:25.7 PL:[25.7, 0.0, 217.1] SR:15 DR:4 LR:-25.72 LO:34.54);ALT=T[chr19:54691043[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54691217	+	chr19	54693152	+	.	10	0	6866649_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6866649_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54691217(+)-19:54693152(-)__19_54684001_54709001D;SPAN=1935;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:79 GQ:11.6 PL:[11.6, 0.0, 179.9] SR:0 DR:10 LR:-11.61 LO:20.48);ALT=C[chr19:54693152[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54715185	+	chr19	54719888	+	.	6	3	6866892_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6866892_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54708501_54733501_128C;SPAN=4703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:77 GQ:2.3 PL:[2.3, 0.0, 183.8] SR:3 DR:6 LR:-2.246 LO:13.27);ALT=G[chr19:54719888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54800856	+	chr19	54807621	+	AGATG	22	33	6866846_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;INSERTION=AGATG;MAPQ=0;MATEID=6866846_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_19_54782001_54807001_21C;SPAN=6765;SUBN=9;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:18 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:33 DR:22 LR:-148.5 LO:148.5);ALT=G[chr19:54807621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54819037	+	chr19	54822683	+	.	4	2	6867017_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTGA;MAPQ=60;MATEID=6867017_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_54806501_54831501_212C;SPAN=3646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:81 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:2 DR:4 LR:5.44 LO:8.605);ALT=A[chr19:54822683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54872898	+	chr19	54876380	+	.	46	0	6867202_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6867202_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54872898(+)-19:54876380(-)__19_54855501_54880501D;SPAN=3482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:103 GQ:99 PL:[124.1, 0.0, 124.1] SR:0 DR:46 LR:-123.9 LO:123.9);ALT=A[chr19:54876380[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54960480	+	chr19	54963267	+	.	9	0	6867502_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6867502_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54960480(+)-19:54963267(-)__19_54953501_54978501D;SPAN=2787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:0 DR:9 LR:-8.306 LO:17.99);ALT=T[chr19:54963267[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	54960483	+	chr19	54962465	+	.	9	0	6867503_1	10.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6867503_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:54960483(+)-19:54962465(-)__19_54953501_54978501D;SPAN=1982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:73 GQ:10.1 PL:[10.1, 0.0, 165.2] SR:0 DR:9 LR:-9.932 LO:18.32);ALT=T[chr19:54962465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	55407697	-	chr19	55638661	+	.	10	0	6869596_1	23.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=6869596_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:55407697(-)-19:55638661(-)__19_55615001_55640001D;SPAN=230964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:37 GQ:23 PL:[23.0, 0.0, 65.9] SR:0 DR:10 LR:-22.99 LO:24.18);ALT=[chr19:55638661[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr19	55758445	+	chr19	55767071	+	.	10	0	6870209_1	19.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6870209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:55758445(+)-19:55767071(-)__19_55762001_55787001D;SPAN=8626;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:50 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:0 DR:10 LR:-19.46 LO:22.66);ALT=T[chr19:55767071[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	55897385	+	chr19	55899304	+	.	12	0	6870679_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6870679_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:55897385(+)-19:55899304(-)__19_55884501_55909501D;SPAN=1919;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:12 DP:1168 GQ:99 PL:[0.0, 276.5, 3390.0] SR:0 DR:12 LR:276.8 LO:11.34);ALT=C[chr19:55899304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	55898062	+	chr19	55899297	+	.	0	89	6870685_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6870685_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_55884501_55909501_250C;SPAN=1235;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:89 DP:1211 GQ:33.8 PL:[0.0, 33.8, 3007.0] SR:89 DR:0 LR:34.3 LO:160.1);ALT=G[chr19:55899297[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	55967857	+	chr19	55972879	+	.	41	19	6871088_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6871088_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_55958001_55983001_289C;SPAN=5022;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:106 GQ:99 PL:[123.2, 0.0, 133.1] SR:19 DR:41 LR:-123.1 LO:123.2);ALT=C[chr19:55972879[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56111826	+	chr19	56113436	+	.	33	0	6871337_1	89.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6871337_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:56111826(+)-19:56113436(-)__19_56105001_56130001D;SPAN=1610;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:72 GQ:83 PL:[89.6, 0.0, 83.0] SR:0 DR:33 LR:-89.43 LO:89.43);ALT=A[chr19:56113436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56152549	+	chr19	56153869	+	CTGCCA	30	5	6871804_1	92.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CTGCCA;MAPQ=60;MATEID=6871804_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_56154001_56179001_17C;SPAN=1320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:0 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:5 DR:30 LR:-92.42 LO:92.42);ALT=G[chr19:56153869[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56166531	+	chr19	56170571	+	.	23	0	6871842_1	53.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6871842_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:56166531(+)-19:56170571(-)__19_56154001_56179001D;SPAN=4040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:85 GQ:53 PL:[53.0, 0.0, 152.0] SR:0 DR:23 LR:-52.89 LO:55.62);ALT=G[chr19:56170571[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	56186801	+	chr19	56189891	+	.	36	33	6871691_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6871691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_56178501_56203501_40C;SPAN=3090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:93 GQ:80.6 PL:[143.3, 0.0, 80.6] SR:33 DR:36 LR:-144.0 LO:144.0);ALT=G[chr19:56189891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	57875072	+	chr19	57876181	+	.	12	7	6876953_1	28.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6876953_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_57869001_57894001_238C;SPAN=1109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:79 GQ:28.1 PL:[28.1, 0.0, 163.4] SR:7 DR:12 LR:-28.11 LO:33.61);ALT=G[chr19:57876181[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	57946962	+	chr19	57949468	+	.	0	11	6877182_1	13.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6877182_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_57942501_57967501_139C;SPAN=2506;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:86 GQ:13.1 PL:[13.1, 0.0, 194.6] SR:11 DR:0 LR:-13.01 LO:22.58);ALT=G[chr19:57949468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58816860	+	chr19	58823383	+	.	18	0	6880137_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6880137_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:58816860(+)-19:58823383(-)__19_58800001_58825001D;SPAN=6523;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:113 GQ:29 PL:[29.0, 0.0, 243.5] SR:0 DR:18 LR:-28.8 LO:38.82);ALT=G[chr19:58823383[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58817583	+	chr19	58823530	+	.	0	10	6880139_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6880139_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_58800001_58825001_98C;SPAN=5947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:88 GQ:9.2 PL:[9.2, 0.0, 203.9] SR:10 DR:0 LR:-9.169 LO:19.98);ALT=G[chr19:58823530[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58826404	+	chr19	58838189	+	CCATAAAGGCAGGCCATGCTTATCATCATTGCAGTATCCAATCTGCAGTGGTGCTGGCTGCCTGTTGTGGGTGCTCAGTATTTAT	28	23	6880336_1	99.0	.	DISC_MAPQ=55;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CCATAAAGGCAGGCCATGCTTATCATCATTGCAGTATCCAATCTGCAGTGGTGCTGGCTGCCTGTTGTGGGTGCTCAGTATTTAT;MAPQ=60;MATEID=6880336_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_58824501_58849501_295C;SPAN=11785;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:91 GQ:99 PL:[114.2, 0.0, 104.3] SR:23 DR:28 LR:-114.0 LO:114.0);ALT=T[chr19:58838189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58836729	+	chr19	58838189	+	.	9	5	6880355_1	19.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6880355_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_19_58824501_58849501_295C;SPAN=1460;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:5 DR:9 LR:-19.34 LO:27.64);ALT=T[chr19:58838189[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58898735	+	chr19	58904339	+	.	57	0	6880845_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6880845_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:58898735(+)-19:58904339(-)__19_58898001_58923001D;SPAN=5604;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:149 GQ:99 PL:[147.8, 0.0, 213.8] SR:0 DR:57 LR:-147.8 LO:148.5);ALT=A[chr19:58904339[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58899613	+	chr19	58905862	+	.	0	10	6880850_1	0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6880850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_58898001_58923001_139C;SPAN=6249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:384 GQ:70.7 PL:[0.0, 70.7, 1073.0] SR:10 DR:0 LR:71.03 LO:13.42);ALT=G[chr19:58905862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	58899613	+	chr19	58904350	+	GGTAAT	9	479	6880849_1	99.0	.	DISC_MAPQ=35;EVDNC=ASDIS;HOMSEQ=CCTGCACTGTGAGGCAGGTACTTGGCATACTTCTCCTTCACTGCAA;INSERTION=GGTAAT;MAPQ=0;MATEID=6880849_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_19_58898001_58923001_318C;SECONDARY;SPAN=4737;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:487 DP:299 GQ:99 PL:[1446.0, 131.7, 0.0] SR:479 DR:9 LR:-1446.0 LO:1446.0);ALT=G[chr19:58904350[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	59063806	+	chr19	59065411	+	.	45	58	6880793_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6880793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_59045001_59070001_254C;SPAN=1605;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:85 DP:110 GQ:16.4 PL:[250.7, 0.0, 16.4] SR:58 DR:45 LR:-263.1 LO:263.1);ALT=C[chr19:59065411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	59063850	+	chr19	59066304	+	.	16	0	6880794_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6880794_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=19:59063850(+)-19:59066304(-)__19_59045001_59070001D;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:96 GQ:26.9 PL:[26.9, 0.0, 205.1] SR:0 DR:16 LR:-26.81 LO:34.85);ALT=C[chr19:59066304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr19	59086955	+	chr19	59092610	+	.	19	5	6880999_1	53.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6880999_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_19_59069501_59094501_71C;SPAN=5655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:70 GQ:53.6 PL:[53.6, 0.0, 116.3] SR:5 DR:19 LR:-53.66 LO:54.93);ALT=G[chr19:59092610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	814594	+	chr20	825348	+	.	3	2	6884052_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6884052_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_808501_833501_158C;SPAN=10754;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:103 GQ:14.4 PL:[0.0, 14.4, 277.2] SR:2 DR:3 LR:14.7 LO:6.063);ALT=G[chr20:825348[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1099545	+	chr20	1106137	+	.	0	41	6885460_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=6885460_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_1078001_1103001_5C;SPAN=6592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:90 GQ:99 PL:[110.9, 0.0, 107.6] SR:41 DR:0 LR:-111.0 LO:111.0);ALT=G[chr20:1106137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1106294	+	chr20	1108068	+	.	0	7	6885491_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6885491_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_1102501_1127501_272C;SPAN=1774;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:95 GQ:2.4 PL:[0.0, 2.4, 234.3] SR:7 DR:0 LR:2.631 LO:12.6);ALT=G[chr20:1108068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1389146	+	chr20	1390815	+	.	67	38	6886506_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACA;MAPQ=60;MATEID=6886506_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_20_1372001_1397001_298C;SPAN=1669;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:93 DP:94 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:38 DR:67 LR:-277.3 LO:277.3);ALT=A[chr20:1390815[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1438923	+	chr20	1447365	+	GGGCTGTGCCTCTGGACACTGAACTGGGGGTTGCCTGCGAAATGGTCACAATGTCTTCATCCCCTCCGTCCTCATAAAAGCTCGCTAGCGCGAT	0	27	6886723_1	74.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=GGGCTGTGCCTCTGGACACTGAACTGGGGGTTGCCTGCGAAATGGTCACAATGTCTTCATCCCCTCCGTCCTCATAAAAGCTCGCTAGCGCGAT;MAPQ=60;MATEID=6886723_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_1445501_1470501_177C;SPAN=8442;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:54 GQ:54.8 PL:[74.6, 0.0, 54.8] SR:27 DR:0 LR:-74.63 LO:74.63);ALT=G[chr20:1447365[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1445117	+	chr20	1447416	+	.	16	0	6886726_1	39.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=6886726_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:1445117(+)-20:1447416(-)__20_1445501_1470501D;SPAN=2299;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:48 GQ:39.8 PL:[39.8, 0.0, 76.1] SR:0 DR:16 LR:-39.81 LO:40.45);ALT=C[chr20:1447416[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	1561036	+	chr20	1594065	+	.	9	0	6887035_1	19.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6887035_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:1561036(+)-20:1594065(-)__20_1592501_1617501D;SPAN=33029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:39 GQ:19.1 PL:[19.1, 0.0, 75.2] SR:0 DR:9 LR:-19.14 LO:21.04);ALT=A[chr20:1594065[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2444545	+	chr20	2446354	+	.	3	17	6890165_1	26.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6890165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2425501_2450501_132C;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:147 GQ:26.3 PL:[26.3, 0.0, 329.9] SR:17 DR:3 LR:-26.19 LO:41.64);ALT=T[chr20:2446354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2446465	+	chr20	2448252	+	.	0	67	6890176_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6890176_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2425501_2450501_364C;SPAN=1787;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:67 DP:147 GQ:99 PL:[181.4, 0.0, 174.8] SR:67 DR:0 LR:-181.3 LO:181.3);ALT=C[chr20:2448252[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2446514	+	chr20	2451333	+	.	49	0	6890323_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6890323_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:2446514(+)-20:2451333(-)__20_2450001_2475001D;SPAN=4819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:58 GQ:5.7 PL:[151.8, 5.7, 0.0] SR:0 DR:49 LR:-156.5 LO:156.5);ALT=G[chr20:2451333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2448405	+	chr20	2451334	+	.	118	27	6890324_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6890324_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2450001_2475001_216C;SPAN=2929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:126 DP:59 GQ:33.9 PL:[372.9, 33.9, 0.0] SR:27 DR:118 LR:-373.0 LO:373.0);ALT=C[chr20:2451334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2633570	+	chr20	2635057	+	.	8	0	6890827_1	0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6890827_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:2633570(+)-20:2635057(-)__20_2621501_2646501D;SPAN=1487;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:122 GQ:6.3 PL:[0.0, 6.3, 306.9] SR:0 DR:8 LR:6.645 LO:13.98);ALT=A[chr20:2635057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2634040	+	chr20	2635058	+	.	0	12	6890831_1	9.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6890831_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2621501_2646501_270C;SPAN=1018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:111 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:12 DR:0 LR:-9.539 LO:23.7);ALT=G[chr20:2635058[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2641616	+	chr20	2644091	+	.	8	6	6890869_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6890869_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2621501_2646501_178C;SPAN=2475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:113 GQ:9.2 PL:[9.2, 0.0, 263.3] SR:6 DR:8 LR:-8.998 LO:23.6);ALT=C[chr20:2644091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2779540	+	chr20	2781046	+	.	0	10	6891934_1	0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=6891934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2768501_2793501_353C;SPAN=1506;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:147 GQ:6.6 PL:[0.0, 6.6, 369.6] SR:10 DR:0 LR:6.816 LO:17.64);ALT=C[chr20:2781046[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	2803162	+	chr20	2806410	+	.	49	34	6891520_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAAGAACTTGATTT;MAPQ=60;MATEID=6891520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_2793001_2818001_85C;SPAN=3248;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:70 DP:87 GQ:2.9 PL:[207.5, 0.0, 2.9] SR:34 DR:49 LR:-219.6 LO:219.6);ALT=T[chr20:2806410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3016587	+	chr20	3017795	+	.	0	4	6892501_1	0	.	EVDNC=ASSMB;HOMSEQ=TGCAG;MAPQ=60;MATEID=6892501_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3013501_3038501_307C;SPAN=1208;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:105 GQ:15 PL:[0.0, 15.0, 283.8] SR:4 DR:0 LR:15.24 LO:6.029);ALT=G[chr20:3017795[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3180750	+	chr20	3183859	+	CACGCTGGGCCTTTCGCGCTTGTTTCTCCTCCAGCTTCCGCAGTTTCTTAGCTCCAATTTTCCCCGACAGGTGAGTTTCCGCTGGCTTCTCGACACCTTCCTCCTCCTGGG	2	17	6893206_1	27.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=CACGCTGGGCCTTTCGCGCTTGTTTCTCCTCCAGCTTCCGCAGTTTCTTAGCTCCAATTTTCCCCGACAGGTGAGTTTCCGCTGGCTTCTCGACACCTTCCTCCTCCTGGG;MAPQ=60;MATEID=6893206_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_3160501_3185501_261C;SPAN=3109;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:107 GQ:27.2 PL:[27.2, 0.0, 231.8] SR:17 DR:2 LR:-27.13 LO:36.64);ALT=T[chr20:3183859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3181102	+	chr20	3183859	+	.	0	9	6893207_1	1.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6893207_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_20_3160501_3185501_261C;SPAN=2757;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:9 DR:0 LR:-1.262 LO:16.82);ALT=T[chr20:3183859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3184065	+	chr20	3185183	+	.	37	17	6893221_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=6893221_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3160501_3185501_215C;SPAN=1118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:125 GQ:99 PL:[118.1, 0.0, 184.1] SR:17 DR:37 LR:-118.0 LO:118.8);ALT=G[chr20:3185183[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3190265	+	chr20	3193813	+	.	40	12	6893356_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AGGT;MAPQ=60;MATEID=6893356_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_3185001_3210001_191C;SPAN=3548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:113 GQ:99 PL:[108.2, 0.0, 164.3] SR:12 DR:40 LR:-108.0 LO:108.7);ALT=T[chr20:3193813[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3190265	+	chr20	3194628	+	CGTTCAGATTCTAGGAGATAAGTTTCCATGCACTTTGGTGGCACAGAAAATTGACCTGCCGGAGTACCAGGGGGAGCCGGATGAGATTTCCATACAGAAATGTCAGGAGGCAGTTCGC	28	37	6893357_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAGGT;INSERTION=CGTTCAGATTCTAGGAGATAAGTTTCCATGCACTTTGGTGGCACAGAAAATTGACCTGCCGGAGTACCAGGGGGAGCCGGATGAGATTTCCATACAGAAATGTCAGGAGGCAGTTCGC;MAPQ=60;MATEID=6893357_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_3185001_3210001_191C;SPAN=4363;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:64 DP:117 GQ:99 PL:[179.6, 0.0, 103.7] SR:37 DR:28 LR:-180.6 LO:180.6);ALT=T[chr20:3194628[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3190271	+	chr20	3199160	+	.	15	0	6893358_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6893358_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:3190271(+)-20:3199160(-)__20_3185001_3210001D;SPAN=8889;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:109 GQ:20 PL:[20.0, 0.0, 244.4] SR:0 DR:15 LR:-19.98 LO:31.31);ALT=G[chr20:3199160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3194704	+	chr20	3199161	+	AAAGTGGTTTCTGGAGAAGTTAAAGCCTGA	2	33	6893378_1	74.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAAGTGGTTTCTGGAGAAGTTAAAGCCTGA;MAPQ=60;MATEID=6893378_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3185001_3210001_288C;SPAN=4457;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:128 GQ:74.3 PL:[74.3, 0.0, 236.0] SR:33 DR:2 LR:-74.26 LO:78.98);ALT=T[chr20:3199161[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3363156	+	chr20	3388122	+	.	5	6	6894122_1	12.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=6894122_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_3356501_3381501_359C;SPAN=24966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:6 DR:5 LR:-12.59 LO:17.19);ALT=G[chr20:3388122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3736256	+	chr20	3740728	+	TGACCAGAAAGCTGCTGTCACTCTCCTGGGTGACCATGACCACCGAGTCATGCAGCTTCTCATCAAAGTGGACGTGGCTGTGGGATCCTTCTGCATCGTGGCCTGCCGCAAAGCGGATACTCCGGACTCTGGGCTTGTTG	0	47	6895351_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGACCAGAAAGCTGCTGTCACTCTCCTGGGTGACCATGACCACCGAGTCATGCAGCTTCTCATCAAAGTGGACGTGGCTGTGGGATCCTTCTGCATCGTGGCCTGCCGCAAAGCGGATACTCCGGACTCTGGGCTTGTTG;MAPQ=60;MATEID=6895351_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_3724001_3749001_364C;SPAN=4472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:98 GQ:99 PL:[128.6, 0.0, 108.8] SR:47 DR:0 LR:-128.7 LO:128.7);ALT=T[chr20:3740728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3739374	+	chr20	3748330	+	.	25	0	6895367_1	55.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6895367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:3739374(+)-20:3748330(-)__20_3724001_3749001D;SPAN=8956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:99 GQ:55.7 PL:[55.7, 0.0, 184.4] SR:0 DR:25 LR:-55.7 LO:59.57);ALT=A[chr20:3748330[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3740835	+	chr20	3748309	+	.	32	11	6895379_1	82.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6895379_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3724001_3749001_394C;SPAN=7474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:99 GQ:82.1 PL:[82.1, 0.0, 158.0] SR:11 DR:32 LR:-82.11 LO:83.43);ALT=T[chr20:3748309[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3870579	+	chr20	3888572	+	.	6	2	6896604_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6896604_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_3846501_3871501_443C;SPAN=17993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:49 GQ:9.8 PL:[9.8, 0.0, 108.8] SR:2 DR:6 LR:-9.832 LO:14.73);ALT=G[chr20:3888572[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3944713	+	chr20	3996112	+	.	19	0	6896765_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6896765_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:3944713(+)-20:3996112(-)__20_3993501_4018501D;SPAN=51399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:28 GQ:12.2 PL:[55.1, 0.0, 12.2] SR:0 DR:19 LR:-56.61 LO:56.61);ALT=T[chr20:3996112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	3970516	+	chr20	3995974	+	.	23	0	6896768_1	66.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6896768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:3970516(+)-20:3995974(-)__20_3993501_4018501D;SPAN=25458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:23 DP:23 GQ:6 PL:[66.0, 6.0, 0.0] SR:0 DR:23 LR:-66.02 LO:66.02);ALT=T[chr20:3995974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	4129626	+	chr20	4155675	+	.	7	4	6897208_1	17.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=6897208_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_4116001_4141001_348C;SPAN=26049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:22 GQ:17.3 PL:[17.3, 0.0, 33.8] SR:4 DR:7 LR:-17.15 LO:17.52);ALT=T[chr20:4155675[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	4667195	+	chr20	4679859	+	.	13	0	6899369_1	30.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6899369_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:4667195(+)-20:4679859(-)__20_4679501_4704501D;SPAN=12664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:0 DR:13 LR:-30.18 LO:31.58);ALT=A[chr20:4679859[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	4781708	+	chr20	4802974	+	.	0	7	6899890_1	10.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6899890_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_4802001_4827001_173C;SPAN=21266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:46 GQ:10.7 PL:[10.7, 0.0, 99.8] SR:7 DR:0 LR:-10.64 LO:14.94);ALT=C[chr20:4802974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5090140	+	chr20	5093480	+	.	11	0	6900932_1	7.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=6900932_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:5090140(+)-20:5093480(-)__20_5071501_5096501D;SPAN=3340;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:106 GQ:7.7 PL:[7.7, 0.0, 248.6] SR:0 DR:11 LR:-7.593 LO:21.52);ALT=T[chr20:5093480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5092252	+	chr20	5093607	+	.	6	3	6900947_1	0	.	DISC_MAPQ=49;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6900947_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_5071501_5096501_425C;SECONDARY;SPAN=1355;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:111 GQ:9.9 PL:[0.0, 9.9, 287.1] SR:3 DR:6 LR:10.27 LO:9.971);ALT=C[chr20:5093607[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5096239	+	chr20	5098111	+	.	9	0	6901237_1	8.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=6901237_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:5096239(+)-20:5098111(-)__20_5096001_5121001D;SPAN=1872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:79 GQ:8.3 PL:[8.3, 0.0, 183.2] SR:0 DR:9 LR:-8.306 LO:17.99);ALT=C[chr20:5098111[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5107796	+	chr20	5154167	+	.	13	4	6901334_1	31.0	.	DISC_MAPQ=57;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=6901334_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_20_5145001_5170001_36C;SPAN=46371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:44 GQ:31.1 PL:[31.1, 0.0, 74.0] SR:4 DR:13 LR:-30.99 LO:32.03);ALT=G[chr20:5154167[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5731166	+	chr20	5753775	+	.	8	0	6904133_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6904133_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:5731166(+)-20:5753775(-)__20_5708501_5733501D;SPAN=22609;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.3 LO:18.03);ALT=G[chr20:5753775[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	5731177	+	chr20	5753505	+	.	20	0	6904134_1	53.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6904134_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:5731177(+)-20:5753505(-)__20_5708501_5733501D;SPAN=22328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:47 GQ:53.3 PL:[53.3, 0.0, 59.9] SR:0 DR:20 LR:-53.29 LO:53.31);ALT=C[chr20:5753505[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16710805	+	chr20	16712805	+	.	38	0	6938933_1	94.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6938933_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:16710805(+)-20:16712805(-)__20_16709001_16734001D;SPAN=2000;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:38 DP:114 GQ:94.7 PL:[94.7, 0.0, 180.5] SR:0 DR:38 LR:-94.55 LO:96.07);ALT=C[chr20:16712805[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16710809	+	chr20	16712312	+	.	19	23	6938934_1	73.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6938934_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_16709001_16734001_12C;SPAN=1503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:120 GQ:73.1 PL:[73.1, 0.0, 218.3] SR:23 DR:19 LR:-73.12 LO:77.14);ALT=G[chr20:16712312[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	16712981	+	chr20	16717905	+	.	4	18	6938942_1	44.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=C;MAPQ=7;MATEID=6938942_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_16709001_16734001_14C;SPAN=4924;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:106 GQ:44 PL:[44.0, 0.0, 212.3] SR:18 DR:4 LR:-43.9 LO:50.26);ALT=G[chr20:16717905[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	17550857	+	chr20	17581382	+	.	38	14	6941437_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6941437_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=GG;SCTG=c_20_17542001_17567001_402C;SECONDARY;SPAN=30525;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:45 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:14 DR:38 LR:-151.8 LO:151.8);ALT=G[chr20:17581382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	17641176	+	chr20	17662671	+	.	9	7	6941853_1	32.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ACCTG;MAPQ=60;MATEID=6941853_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_17640001_17665001_234C;SPAN=21495;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:7 DR:9 LR:-31.91 LO:35.06);ALT=G[chr20:17662671[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	17937683	+	chr20	17949018	+	.	4	20	6942909_1	44.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=37;MATEID=6942909_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_17934001_17959001_351C;SPAN=11335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:118 GQ:44 PL:[44.0, 0.0, 242.0] SR:20 DR:4 LR:-43.95 LO:51.84);ALT=T[chr20:17949018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	18191155	+	chr20	18189739	+	.	34	0	6944072_1	90.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6944072_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:18189739(-)-20:18191155(+)__20_18179001_18204001D;SPAN=1416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:80 GQ:90.5 PL:[90.5, 0.0, 103.7] SR:0 DR:34 LR:-90.56 LO:90.61);ALT=]chr20:18191155]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	18548240	+	chr20	18549881	+	.	78	50	6945633_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6945633_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_18546501_18571501_261C;SPAN=1641;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:151 GQ:74.9 PL:[289.4, 0.0, 74.9] SR:50 DR:78 LR:-296.0 LO:296.0);ALT=G[chr20:18549881[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	18568759	+	chr20	18574373	+	.	23	15	6945730_1	74.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=6945730_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_18571001_18596001_345C;SPAN=5614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:68 GQ:74 PL:[74.0, 0.0, 90.5] SR:15 DR:23 LR:-74.01 LO:74.1);ALT=G[chr20:18574373[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	18568781	+	chr20	18576649	+	.	25	0	6945731_1	66.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=6945731_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:18568781(+)-20:18576649(-)__20_18571001_18596001D;SPAN=7868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:61 GQ:66.2 PL:[66.2, 0.0, 79.4] SR:0 DR:25 LR:-66.0 LO:66.1);ALT=C[chr20:18576649[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	18574466	+	chr20	18576650	+	.	3	28	6945746_1	67.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6945746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_18571001_18596001_379C;SPAN=2184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:129 GQ:67.4 PL:[67.4, 0.0, 245.6] SR:28 DR:3 LR:-67.38 LO:73.09);ALT=G[chr20:18576650[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	19998089	+	chr20	20007427	+	.	18	0	6950194_1	31.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6950194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:19998089(+)-20:20007427(-)__20_19992001_20017001D;SPAN=9338;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:104 GQ:31.4 PL:[31.4, 0.0, 219.5] SR:0 DR:18 LR:-31.24 LO:39.53);ALT=A[chr20:20007427[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	19998089	+	chr20	20006320	+	.	19	0	6950193_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6950193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:19998089(+)-20:20006320(-)__20_19992001_20017001D;SPAN=8231;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:89 GQ:38.6 PL:[38.6, 0.0, 177.2] SR:0 DR:19 LR:-38.61 LO:43.67);ALT=A[chr20:20006320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	20006411	+	chr20	20007428	+	.	0	19	6950218_1	31.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6950218_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_19992001_20017001_96C;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:116 GQ:31.4 PL:[31.4, 0.0, 249.2] SR:19 DR:0 LR:-31.29 LO:41.22);ALT=A[chr20:20007428[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	20007563	+	chr20	20013148	+	.	2	6	6950225_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAAG;MAPQ=60;MATEID=6950225_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_19992001_20017001_99C;SPAN=5585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:102 GQ:4.2 PL:[0.0, 4.2, 254.1] SR:6 DR:2 LR:4.527 LO:12.38);ALT=G[chr20:20013148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	20031269	+	chr20	20032934	+	.	11	6	6950300_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTT;MAPQ=60;MATEID=6950300_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_20016501_20041501_288C;SPAN=1665;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:98 GQ:13.1 PL:[13.1, 0.0, 224.3] SR:6 DR:11 LR:-13.06 LO:24.39);ALT=T[chr20:20032934[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	20336634	+	chr20	20335485	+	.	32	0	6951625_1	75.0	.	DISC_MAPQ=28;EVDNC=DSCRD;IMPRECISE;MAPQ=28;MATEID=6951625_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:20335485(-)-20:20336634(+)__20_20335001_20360001D;SPAN=1149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:112 GQ:75.5 PL:[75.5, 0.0, 194.3] SR:0 DR:32 LR:-75.29 LO:78.28);ALT=]chr20:20336634]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	21284111	+	chr20	21306915	+	.	87	22	6954551_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6954551_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_21290501_21315501_193C;SPAN=22804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:57 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:22 DR:87 LR:-270.7 LO:270.7);ALT=G[chr20:21306915[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	21286127	+	chr20	21288773	+	.	98	40	6954360_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CCATGTTGGCCAGGCTGGTCTCGAACTCCTGACCTCA;MAPQ=60;MATEID=6954360_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_20_21266001_21291001_41C;SPAN=2646;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:29 GQ:34.8 PL:[382.8, 34.8, 0.0] SR:40 DR:98 LR:-382.9 LO:382.9);ALT=A[chr20:21288773[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	21307240	+	chr20	21309196	+	.	2	8	6954624_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6954624_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_21290501_21315501_102C;SPAN=1956;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:8 DR:2 LR:3.394 LO:14.36);ALT=G[chr20:21309196[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	21313078	+	chr20	21314180	+	.	4	4	6954649_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6954649_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_21290501_21315501_389C;SPAN=1102;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:94 GQ:1.1 PL:[1.1, 0.0, 225.5] SR:4 DR:4 LR:-0.9411 LO:14.92);ALT=G[chr20:21314180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	21321490	+	chr20	21324728	+	.	0	7	6954494_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6954494_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_21315001_21340001_166C;SPAN=3238;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:93 GQ:1.8 PL:[0.0, 1.8, 227.7] SR:7 DR:0 LR:2.089 LO:12.67);ALT=T[chr20:21324728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	23331698	+	chr20	23334614	+	.	0	18	6960817_1	27.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=6960817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_23324001_23349001_174C;SPAN=2916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:118 GQ:27.5 PL:[27.5, 0.0, 258.5] SR:18 DR:0 LR:-27.45 LO:38.44);ALT=G[chr20:23334614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	23614637	+	chr20	23615891	+	.	0	32	6961793_1	46.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6961793_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_23593501_23618501_247C;SPAN=1254;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:218 GQ:46.6 PL:[46.6, 0.0, 482.3] SR:32 DR:0 LR:-46.57 LO:67.76);ALT=C[chr20:23615891[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	23616006	+	chr20	23618257	+	.	24	66	6961839_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6961839_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_23618001_23643001_3C;SPAN=2251;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:90 DP:187 GQ:99 PL:[246.5, 0.0, 206.9] SR:66 DR:24 LR:-246.6 LO:246.6);ALT=T[chr20:23618257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	24930211	+	chr20	24937920	+	.	0	9	6965810_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=6965810_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_24916501_24941501_385C;SPAN=7709;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:9 DR:0 LR:-3.971 LO:17.23);ALT=G[chr20:24937920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	24959521	+	chr20	24964539	+	.	0	17	6966077_1	26.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6966077_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_24941001_24966001_76C;SPAN=5018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:109 GQ:26.6 PL:[26.6, 0.0, 237.8] SR:17 DR:0 LR:-26.59 LO:36.49);ALT=G[chr20:24964539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	24959565	+	chr20	24973276	+	.	9	0	6966178_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6966178_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:24959565(+)-20:24973276(-)__20_24965501_24990501D;SPAN=13711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=G[chr20:24973276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	24964660	+	chr20	24973230	+	.	23	5	6966179_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGCC;MAPQ=60;MATEID=6966179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_24965501_24990501_339C;SPAN=8570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:59 GQ:63.2 PL:[63.2, 0.0, 79.7] SR:5 DR:23 LR:-63.24 LO:63.35);ALT=C[chr20:24973230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	25319991	+	chr20	25371148	+	.	0	7	6967809_1	7.0	.	EVDNC=ASSMB;HOMSEQ=CCTGC;MAPQ=60;MATEID=6967809_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_25308501_25333501_160C;SPAN=51157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:57 GQ:7.7 PL:[7.7, 0.0, 129.8] SR:7 DR:0 LR:-7.664 LO:14.24);ALT=C[chr20:25371148[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	26299409	+	chr20	26300542	+	.	30	0	6971378_1	84.0	.	DISC_MAPQ=43;EVDNC=DSCRD;IMPRECISE;MAPQ=43;MATEID=6971378_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:26299409(+)-20:26300542(-)__20_26288501_26313501D;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:55 GQ:47.9 PL:[84.2, 0.0, 47.9] SR:0 DR:30 LR:-84.61 LO:84.61);ALT=A[chr20:26300542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30102537	+	chr20	30115285	+	.	0	37	6973999_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=6973999_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30110501_30135501_252C;SPAN=12748;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:63 GQ:45.8 PL:[105.2, 0.0, 45.8] SR:37 DR:0 LR:-106.2 LO:106.2);ALT=G[chr20:30115285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30154098	+	chr20	30156919	+	.	2	2	6974277_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=60;MATEID=6974277_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30135001_30160001_171C;SPAN=2821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:108 GQ:15.9 PL:[0.0, 15.9, 293.7] SR:2 DR:2 LR:16.06 LO:5.98);ALT=G[chr20:30156919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30536686	+	chr20	30538115	+	.	0	12	6975873_1	17.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6975873_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30527001_30552001_62C;SPAN=1429;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:84 GQ:17 PL:[17.0, 0.0, 185.3] SR:12 DR:0 LR:-16.85 LO:25.26);ALT=C[chr20:30538115[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30538193	+	chr20	30539678	+	.	0	12	6975881_1	9.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6975881_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30527001_30552001_146C;SPAN=1485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:111 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:12 DR:0 LR:-9.539 LO:23.7);ALT=G[chr20:30539678[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30640290	+	chr20	30659462	+	.	0	13	6976539_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6976539_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30649501_30674501_258C;SPAN=19172;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:78 GQ:21.8 PL:[21.8, 0.0, 167.0] SR:13 DR:0 LR:-21.78 LO:28.31);ALT=G[chr20:30659462[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30686939	+	chr20	30689117	+	.	7	3	6976473_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=6976473_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30674001_30699001_90C;SPAN=2178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:123 GQ:6.6 PL:[0.0, 6.6, 310.2] SR:3 DR:7 LR:6.916 LO:13.95);ALT=G[chr20:30689117[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	30723977	+	chr20	30729299	+	.	0	7	6976640_1	0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=6976640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_30723001_30748001_230C;SPAN=5322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:112 GQ:6.9 PL:[0.0, 6.9, 283.8] SR:7 DR:0 LR:7.237 LO:12.09);ALT=G[chr20:30729299[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31292708	+	chr20	31294385	+	.	3	8	6979463_1	9.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=6979463_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TT;SCTG=c_20_31286501_31311501_469C;SPAN=1677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:101 GQ:9.2 PL:[9.2, 0.0, 233.6] SR:8 DR:3 LR:-8.948 LO:21.76);ALT=T[chr20:31294385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31292708	+	chr20	31315697	+	TTTCAGAAAAGTAAGTGGCTTTCTCCTCACTAAGACCCAGAGTTATGAAATCCGCCTGGACCTGCTTGGCTGTGAGACTCTTCTTCAAAG	2	25	6979464_1	75.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CACC;INSERTION=TTTCAGAAAAGTAAGTGGCTTTCTCCTCACTAAGACCCAGAGTTATGAAATCCGCCTGGACCTGCTTGGCTGTGAGACTCTTCTTCAAAG;MAPQ=60;MATEID=6979464_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_31286501_31311501_469C;SPAN=22989;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:52 GQ:48.8 PL:[75.2, 0.0, 48.8] SR:25 DR:2 LR:-75.28 LO:75.28);ALT=T[chr20:31315697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31294610	+	chr20	31331180	+	.	22	0	6979275_1	45.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6979275_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31294610(+)-20:31331180(-)__20_31311001_31336001D;SPAN=36570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:99 GQ:45.8 PL:[45.8, 0.0, 194.3] SR:0 DR:22 LR:-45.8 LO:51.0);ALT=G[chr20:31331180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31310872	+	chr20	31312779	+	TAAT	23	20	6979567_1	99.0	.	DISC_MAPQ=31;EVDNC=ASDIS;INSERTION=TAAT;MAPQ=60;MATEID=6979567_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_31286501_31311501_242C;SPAN=1907;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:35 DP:23 GQ:9.3 PL:[102.3, 9.3, 0.0] SR:20 DR:23 LR:-102.3 LO:102.3);ALT=A[chr20:31312779[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31316016	+	chr20	31331112	+	.	130	0	6979298_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6979298_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31316016(+)-20:31331112(-)__20_31311001_31336001D;SPAN=15096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:130 DP:126 GQ:35.1 PL:[386.1, 35.1, 0.0] SR:0 DR:130 LR:-386.2 LO:386.2);ALT=G[chr20:31331112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31407870	+	chr20	31413729	+	.	22	0	6979687_1	56.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6979687_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31407870(+)-20:31413729(-)__20_31384501_31409501D;SPAN=5859;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:61 GQ:56.3 PL:[56.3, 0.0, 89.3] SR:0 DR:22 LR:-56.1 LO:56.57);ALT=G[chr20:31413729[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31407876	+	chr20	31421518	+	.	22	0	6979688_1	56.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6979688_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31407876(+)-20:31421518(-)__20_31384501_31409501D;SPAN=13642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:62 GQ:56 PL:[56.0, 0.0, 92.3] SR:0 DR:22 LR:-55.83 LO:56.37);ALT=G[chr20:31421518[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31413855	+	chr20	31421519	+	.	0	20	6979724_1	38.0	.	DISC_MAPQ=255;EVDNC=TSI_L;HOMSEQ=TCAGG;MAPQ=60;MATEID=6979724_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_20_31409001_31434001_231C;SPAN=7664;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:102 GQ:38.6 PL:[38.6, 0.0, 206.9] SR:20 DR:0 LR:-38.39 LO:45.13);ALT=G[chr20:31421519[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	31984844	+	chr20	31989258	+	.	16	0	6981925_1	16.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6981925_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:31984844(+)-20:31989258(-)__20_31972501_31997501D;SPAN=4414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:134 GQ:16.7 PL:[16.7, 0.0, 307.1] SR:0 DR:16 LR:-16.51 LO:32.33);ALT=T[chr20:31989258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32399464	+	chr20	32436272	+	.	3	15	6983916_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6983916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32389001_32414001_323C;SPAN=36808;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:75 GQ:39.2 PL:[39.2, 0.0, 141.5] SR:15 DR:3 LR:-39.1 LO:42.43);ALT=G[chr20:32436272[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32581940	+	chr20	32659871	+	.	34	4	6985114_1	97.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6985114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32658501_32683501_315C;SPAN=77931;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:79 GQ:94.1 PL:[97.4, 0.0, 94.1] SR:4 DR:34 LR:-97.44 LO:97.44);ALT=G[chr20:32659871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32581942	+	chr20	32619327	+	.	40	53	6984726_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGAG;MAPQ=60;MATEID=6984726_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32560501_32585501_62C;SPAN=37385;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:60 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:53 DR:40 LR:-208.0 LO:208.0);ALT=G[chr20:32619327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32619413	+	chr20	32659871	+	.	18	30	6985115_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTG;MAPQ=60;MATEID=6985115_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32658501_32683501_102C;SPAN=40458;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:79 GQ:57.8 PL:[133.7, 0.0, 57.8] SR:30 DR:18 LR:-135.4 LO:135.4);ALT=G[chr20:32659871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32660136	+	chr20	32661368	+	.	0	10	6985122_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=6985122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32658501_32683501_373C;SPAN=1232;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:143 GQ:5.4 PL:[0.0, 5.4, 356.4] SR:10 DR:0 LR:5.732 LO:17.77);ALT=G[chr20:32661368[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32665052	+	chr20	32667713	+	AACACAGCCAGGACACAGACGCGGATGATGGGGCCTTGCAGTAAG	7	26	6985150_1	70.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=AACACAGCCAGGACACAGACGCGGATGATGGGGCCTTGCAGTAAG;MAPQ=60;MATEID=6985150_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_32658501_32683501_139C;SPAN=2661;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:131 GQ:70.4 PL:[70.4, 0.0, 245.3] SR:26 DR:7 LR:-70.14 LO:75.71);ALT=G[chr20:32667713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32666359	+	chr20	32667713	+	.	10	22	6985152_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=6985152_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_32658501_32683501_139C;SPAN=1354;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:129 GQ:60.8 PL:[60.8, 0.0, 252.2] SR:22 DR:10 LR:-60.78 LO:67.4);ALT=G[chr20:32667713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32693371	+	chr20	32699909	+	.	12	0	6984915_1	15.0	.	DISC_MAPQ=12;EVDNC=DSCRD;IMPRECISE;MAPQ=12;MATEID=6984915_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:32693371(+)-20:32699909(-)__20_32683001_32708001D;SPAN=6538;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:91 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:0 DR:12 LR:-14.96 LO:24.81);ALT=C[chr20:32699909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32815938	+	chr20	32819226	+	.	78	25	6985680_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAGAACTTTC;MAPQ=60;MATEID=6985680_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32805501_32830501_34C;SPAN=3288;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:109 DP:610 GQ:99 PL:[194.6, 0.0, 1287.0] SR:25 DR:78 LR:-194.5 LO:241.1);ALT=C[chr20:32819226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32881964	+	chr20	32883198	+	.	0	29	6985735_1	61.0	.	EVDNC=ASSMB;HOMSEQ=CACCT;MAPQ=60;MATEID=6985735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32879001_32904001_241C;SPAN=1234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:126 GQ:61.7 PL:[61.7, 0.0, 243.2] SR:29 DR:0 LR:-61.59 LO:67.74);ALT=T[chr20:32883198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32882001	+	chr20	32891051	+	.	9	0	6985736_1	4.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=6985736_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:32882001(+)-20:32891051(-)__20_32879001_32904001D;SPAN=9050;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:95 GQ:4.1 PL:[4.1, 0.0, 225.2] SR:0 DR:9 LR:-3.971 LO:17.23);ALT=G[chr20:32891051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32883392	+	chr20	32891049	+	.	91	15	6985741_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6985741_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_32879001_32904001_160C;SPAN=7657;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:95 DP:109 GQ:19.5 PL:[303.6, 19.5, 0.0] SR:15 DR:91 LR:-307.6 LO:307.6);ALT=C[chr20:32891049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	32951201	+	chr20	32957198	+	.	20	0	6986707_1	51.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6986707_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:32951201(+)-20:32957198(-)__20_32928001_32953001D;SPAN=5997;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:53 GQ:51.8 PL:[51.8, 0.0, 74.9] SR:0 DR:20 LR:-51.66 LO:51.93);ALT=G[chr20:32957198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33104318	+	chr20	33128381	+	.	8	0	6987148_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6987148_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33104318(+)-20:33128381(-)__20_33099501_33124501D;SPAN=24063;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:48 GQ:13.4 PL:[13.4, 0.0, 102.5] SR:0 DR:8 LR:-13.4 LO:17.42);ALT=A[chr20:33128381[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33104318	+	chr20	33122429	+	.	61	0	6987147_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6987147_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33104318(+)-20:33122429(-)__20_33099501_33124501D;SPAN=18111;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:113 GQ:99 PL:[170.9, 0.0, 101.6] SR:0 DR:61 LR:-171.6 LO:171.6);ALT=A[chr20:33122429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33114149	+	chr20	33122430	+	.	4	17	6987179_1	34.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6987179_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33099501_33124501_108C;SPAN=8281;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:128 GQ:34.7 PL:[34.7, 0.0, 275.6] SR:17 DR:4 LR:-34.64 LO:45.58);ALT=G[chr20:33122430[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33122599	+	chr20	33128382	+	.	6	23	6987203_1	83.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=6987203_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33099501_33124501_363C;SPAN=5783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:44 GQ:21.2 PL:[83.9, 0.0, 21.2] SR:23 DR:6 LR:-85.73 LO:85.73);ALT=G[chr20:33128382[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33464626	+	chr20	33470596	+	.	8	13	6988919_1	43.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6988919_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33467001_33492001_100C;SPAN=5970;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:61 GQ:43.1 PL:[43.1, 0.0, 102.5] SR:13 DR:8 LR:-42.89 LO:44.34);ALT=G[chr20:33470596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33530814	+	chr20	33539525	+	AAGAGTTTGCTCCAGGAAGGCAGCGTTCTGGCTGACAGCATCCACTAGCAGGTTGAAGTCCATCTGCACAGCATAGGCTTGCTCCAGCAGGGCACTGGGGACCAGTGAGGGGAAGAGCGTGAATGGGGCATAGCTCACC	2	41	6988674_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=AAGAGTTTGCTCCAGGAAGGCAGCGTTCTGGCTGACAGCATCCACTAGCAGGTTGAAGTCCATCTGCACAGCATAGGCTTGCTCCAGCAGGGCACTGGGGACCAGTGAGGGGAAGAGCGTGAATGGGGCATAGCTCACC;MAPQ=60;MATEID=6988674_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_33516001_33541001_28C;SPAN=8711;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:125 GQ:99 PL:[101.6, 0.0, 200.6] SR:41 DR:2 LR:-101.5 LO:103.3);ALT=A[chr20:33539525[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33533954	+	chr20	33543526	+	.	20	0	6988742_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6988742_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33533954(+)-20:33543526(-)__20_33540501_33565501D;SPAN=9572;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:51 GQ:52.4 PL:[52.4, 0.0, 68.9] SR:0 DR:20 LR:-52.2 LO:52.37);ALT=G[chr20:33543526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33539663	+	chr20	33543528	+	.	28	5	6988743_1	84.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=6988743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33540501_33565501_158C;SPAN=3865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:53 GQ:41.9 PL:[84.8, 0.0, 41.9] SR:5 DR:28 LR:-85.37 LO:85.37);ALT=C[chr20:33543528[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33665980	+	chr20	33680417	+	.	0	11	6989583_1	5.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=6989583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33663001_33688001_286C;SPAN=14437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:113 GQ:5.9 PL:[5.9, 0.0, 266.6] SR:11 DR:0 LR:-5.697 LO:21.19);ALT=G[chr20:33680417[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33859950	+	chr20	33865849	+	.	8	2	6990246_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=6990246_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33859001_33884001_104C;SPAN=5899;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:135 GQ:6.6 PL:[0.0, 6.6, 339.9] SR:2 DR:8 LR:6.866 LO:15.8);ALT=T[chr20:33865849[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33867922	+	chr20	33871978	+	.	3	8	6990276_1	3.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6990276_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33859001_33884001_322C;SPAN=4056;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:120 GQ:3.8 PL:[3.8, 0.0, 287.6] SR:8 DR:3 LR:-3.8 LO:20.89);ALT=C[chr20:33871978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33868633	+	chr20	33871978	+	.	2	42	6990279_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=6990279_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_33859001_33884001_15C;SPAN=3345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:150 GQ:99 PL:[104.6, 0.0, 259.7] SR:42 DR:2 LR:-104.6 LO:108.2);ALT=C[chr20:33871978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33868676	+	chr20	33872230	+	.	10	0	6990280_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=6990280_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33868676(+)-20:33872230(-)__20_33859001_33884001D;SPAN=3554;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:132 GQ:2.4 PL:[0.0, 2.4, 323.4] SR:0 DR:10 LR:2.752 LO:18.13);ALT=T[chr20:33872230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	33868678	+	chr20	33872526	+	.	25	0	6990281_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6990281_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:33868678(+)-20:33872526(-)__20_33859001_33884001D;SPAN=3848;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:132 GQ:47 PL:[47.0, 0.0, 271.4] SR:0 DR:25 LR:-46.76 LO:55.99);ALT=A[chr20:33872526[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34064551	+	chr20	34078713	+	.	13	0	6991003_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6991003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:34064551(+)-20:34078713(-)__20_34055001_34080001D;SPAN=14162;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:110 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:0 DR:13 LR:-13.11 LO:26.21);ALT=A[chr20:34078713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34130690	+	chr20	34135162	+	.	2	10	6991420_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6991420_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34128501_34153501_117C;SPAN=4472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:110 GQ:9.8 PL:[9.8, 0.0, 257.3] SR:10 DR:2 LR:-9.81 LO:23.75);ALT=G[chr20:34135162[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34135259	+	chr20	34136262	+	.	0	11	6991434_1	3.0	.	EVDNC=ASSMB;HOMSEQ=GTG;MAPQ=60;MATEID=6991434_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34128501_34153501_159C;SPAN=1003;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:120 GQ:3.8 PL:[3.8, 0.0, 287.6] SR:11 DR:0 LR:-3.8 LO:20.89);ALT=G[chr20:34136262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34220846	+	chr20	34252682	+	.	72	17	6991850_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6991850_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34202001_34227001_425C;SPAN=31836;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:76 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:17 DR:72 LR:-227.8 LO:227.8);ALT=C[chr20:34252682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34287686	+	chr20	34288715	+	.	0	125	6992185_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CTCAGG;MAPQ=60;MATEID=6992185_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34275501_34300501_255C;SPAN=1029;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:125 DP:208 GQ:99 PL:[356.3, 0.0, 148.3] SR:125 DR:0 LR:-360.9 LO:360.9);ALT=G[chr20:34288715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34320057	+	chr20	34326889	+	.	3	13	6992405_1	40.0	.	DISC_MAPQ=36;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=6992405_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_34324501_34349501_38C;SPAN=6832;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:46 GQ:40.4 PL:[40.4, 0.0, 70.1] SR:13 DR:3 LR:-40.35 LO:40.82);ALT=C[chr20:34326889[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34360037	+	chr20	34389410	+	.	17	0	6992717_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6992717_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:34360037(+)-20:34389410(-)__20_34373501_34398501D;SPAN=29373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:67 GQ:38 PL:[38.0, 0.0, 123.8] SR:0 DR:17 LR:-37.97 LO:40.55);ALT=C[chr20:34389410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34360042	+	chr20	34430493	+	.	21	0	6992855_1	52.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6992855_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:34360042(+)-20:34430493(-)__20_34422501_34447501D;SPAN=70451;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:64 GQ:52.1 PL:[52.1, 0.0, 101.6] SR:0 DR:21 LR:-51.98 LO:52.91);ALT=T[chr20:34430493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34360045	+	chr20	34362410	+	.	30	0	6992611_1	69.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6992611_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:34360045(+)-20:34362410(-)__20_34349001_34374001D;SPAN=2365;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:109 GQ:69.5 PL:[69.5, 0.0, 194.9] SR:0 DR:30 LR:-69.5 LO:72.81);ALT=G[chr20:34362410[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	34430667	+	chr20	34446223	+	AATTTCAAATAAATGAGCAGGTCCTTGCTTGCTGGTCTGATTGTCGTTTTTACCCGGCCAAAGTCACTGCTGTTAACAAGGAT	0	12	6992898_1	12.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=GGTA;INSERTION=AATTTCAAATAAATGAGCAGGTCCTTGCTTGCTGGTCTGATTGTCGTTTTTACCCGGCCAAAGTCACTGCTGTTAACAAGGAT;MAPQ=60;MATEID=6992898_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_34422501_34447501_435C;SPAN=15556;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:100 GQ:12.5 PL:[12.5, 0.0, 230.3] SR:12 DR:0 LR:-12.52 LO:24.28);ALT=G[chr20:34446223[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35089954	+	chr20	35125129	+	.	9	0	6995656_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6995656_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35089954(+)-20:35125129(-)__20_35084001_35109001D;SPAN=35175;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:14 GQ:6.2 PL:[26.0, 0.0, 6.2] SR:0 DR:9 LR:-26.43 LO:26.43);ALT=G[chr20:35125129[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35170015	+	chr20	35173268	+	.	16	0	6996003_1	26.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6996003_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35170015(+)-20:35173268(-)__20_35157501_35182501D;SPAN=3253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:99 GQ:26 PL:[26.0, 0.0, 214.1] SR:0 DR:16 LR:-25.99 LO:34.61);ALT=C[chr20:35173268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35234469	+	chr20	35236116	+	.	0	47	6996206_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=6996206_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35231001_35256001_271C;SPAN=1647;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:123 GQ:99 PL:[122.0, 0.0, 174.8] SR:47 DR:0 LR:-121.8 LO:122.4);ALT=G[chr20:35236116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35236221	+	chr20	35238003	+	.	3	14	6996213_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=6996213_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35231001_35256001_166C;SPAN=1782;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:119 GQ:17.3 PL:[17.3, 0.0, 271.4] SR:14 DR:3 LR:-17.28 LO:30.69);ALT=G[chr20:35238003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35521471	+	chr20	35526224	+	.	2	4	6997504_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=6997504_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35500501_35525501_373C;SPAN=4753;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:62 GQ:0 PL:[0.0, 0.0, 148.5] SR:4 DR:2 LR:0.2923 LO:9.206);ALT=T[chr20:35526224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35533951	+	chr20	35540862	+	.	13	0	6997603_1	19.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6997603_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35533951(+)-20:35540862(-)__20_35525001_35550001D;SPAN=6911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:87 GQ:19.4 PL:[19.4, 0.0, 191.0] SR:0 DR:13 LR:-19.34 LO:27.64);ALT=G[chr20:35540862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35539736	+	chr20	35540863	+	.	0	15	6997640_1	24.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=6997640_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35525001_35550001_199C;SPAN=1127;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:94 GQ:24.2 PL:[24.2, 0.0, 202.4] SR:15 DR:0 LR:-24.05 LO:32.36);ALT=C[chr20:35540863[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35540957	+	chr20	35545124	+	.	0	9	6997644_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=6997644_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35525001_35550001_384C;SPAN=4167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:101 GQ:2.6 PL:[2.6, 0.0, 240.2] SR:9 DR:0 LR:-2.346 LO:16.98);ALT=T[chr20:35545124[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35559279	+	chr20	35563431	+	.	2	3	6997996_1	0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=6997996_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_20_35549501_35574501_167C;SPAN=4152;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:104 GQ:14.7 PL:[0.0, 14.7, 280.5] SR:3 DR:2 LR:14.97 LO:6.046);ALT=C[chr20:35563431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35569516	+	chr20	35579839	+	TACTCCAAGATTTTCAAAACGAGACTCATCAAGACAAGGCAGTAATGCGCCTGTGATTTCATTTT	0	37	6998043_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TACTCCAAGATTTTCAAAACGAGACTCATCAAGACAAGGCAGTAATGCGCCTGTGATTTCATTTT;MAPQ=60;MATEID=6998043_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_35549501_35574501_72C;SPAN=10323;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:37 DP:44 GQ:5.1 PL:[115.5, 5.1, 0.0] SR:37 DR:0 LR:-118.0 LO:118.0);ALT=T[chr20:35579839[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35575257	+	chr20	35579919	+	.	11	0	6997709_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6997709_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35575257(+)-20:35579919(-)__20_35574001_35599001D;SPAN=4662;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:113 GQ:5.9 PL:[5.9, 0.0, 266.6] SR:0 DR:11 LR:-5.697 LO:21.19);ALT=T[chr20:35579919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35807826	+	chr20	35826797	+	.	16	0	6999173_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=6999173_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35807826(+)-20:35826797(-)__20_35819001_35844001D;SPAN=18971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:51 GQ:39.2 PL:[39.2, 0.0, 82.1] SR:0 DR:16 LR:-39.0 LO:39.93);ALT=T[chr20:35826797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35807826	+	chr20	35812581	+	.	28	0	6998997_1	56.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6998997_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35807826(+)-20:35812581(-)__20_35794501_35819501D;SPAN=4755;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:133 GQ:56.6 PL:[56.6, 0.0, 264.5] SR:0 DR:28 LR:-56.4 LO:64.16);ALT=T[chr20:35812581[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35812665	+	chr20	35826797	+	.	17	0	6999175_1	42.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6999175_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:35812665(+)-20:35826797(-)__20_35819001_35844001D;SPAN=14132;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:51 GQ:42.5 PL:[42.5, 0.0, 78.8] SR:0 DR:17 LR:-42.3 LO:42.98);ALT=T[chr20:35826797[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35833305	+	chr20	35835674	+	.	3	2	6999247_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=6999247_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35819001_35844001_402C;SPAN=2369;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:112 GQ:16.8 PL:[0.0, 16.8, 303.6] SR:2 DR:3 LR:17.14 LO:5.916);ALT=G[chr20:35835674[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35852373	+	chr20	35854090	+	.	2	4	6999089_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=6999089_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35843501_35868501_112C;SPAN=1717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:125 GQ:17.1 PL:[0.0, 17.1, 336.6] SR:4 DR:2 LR:17.36 LO:7.644);ALT=G[chr20:35854090[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35854205	+	chr20	35856951	+	.	3	5	6999095_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6999095_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_35843501_35868501_285C;SPAN=2746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:114 GQ:4.2 PL:[0.0, 4.2, 283.8] SR:5 DR:3 LR:4.477 LO:14.23);ALT=G[chr20:35856951[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35857148	+	chr20	35860696	+	CTGATGTGGTCATCAAGTTCCCTGAGGAAGAAGCTCCCTCGACTGTCTTGTCCCAGAACCTTTTCACTCCAAAACAGGAAATT	5	21	6999105_1	35.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=CTGATGTGGTCATCAAGTTCCCTGAGGAAGAAGCTCCCTCGACTGTCTTGTCCCAGAACCTTTTCACTCCAAAACAGGAAATT;MAPQ=60;MATEID=6999105_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_35843501_35868501_363C;SPAN=3548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:151 GQ:35.3 PL:[35.3, 0.0, 329.0] SR:21 DR:5 LR:-35.01 LO:49.11);ALT=G[chr20:35860696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35857148	+	chr20	35858375	+	.	8	11	6999104_1	17.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=6999104_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_20_35843501_35868501_363C;SPAN=1227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:121 GQ:17 PL:[17.0, 0.0, 274.4] SR:11 DR:8 LR:-16.73 LO:30.57);ALT=G[chr20:35858375[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35858462	+	chr20	35860696	+	.	2	10	6999116_1	2.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAG;MAPQ=60;MATEID=6999116_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_35843501_35868501_363C;SPAN=2234;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:138 GQ:2.3 PL:[2.3, 0.0, 332.3] SR:10 DR:2 LR:-2.224 LO:22.5);ALT=G[chr20:35860696[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35860794	+	chr20	35862422	+	.	6	17	6999126_1	29.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=6999126_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_20_35843501_35868501_36C;SPAN=1628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:136 GQ:29.3 PL:[29.3, 0.0, 299.9] SR:17 DR:6 LR:-29.17 LO:42.37);ALT=G[chr20:35862422[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35860794	+	chr20	35864982	+	TGGATCCGGATTGGTGCCAATGTCTCCAACTTCACTTTTGCTCCTAGCACGATTATATTTCACCTGGGACATGCT	9	48	6999127_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=TGGATCCGGATTGGTGCCAATGTCTCCAACTTCACTTTTGCTCCTAGCACGATTATATTTCACCTGGGACATGCT;MAPQ=60;MATEID=6999127_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_20_35843501_35868501_36C;SPAN=4188;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:128 GQ:99 PL:[133.7, 0.0, 176.6] SR:48 DR:9 LR:-133.7 LO:134.0);ALT=G[chr20:35864982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	35865112	+	chr20	35869704	+	.	10	20	6999307_1	80.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=6999307_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_20_35868001_35893001_287C;SPAN=4592;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:55 GQ:51.2 PL:[80.9, 0.0, 51.2] SR:20 DR:10 LR:-81.15 LO:81.15);ALT=G[chr20:35869704[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	36147755	+	chr20	36156194	+	.	23	1	7000363_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=7000363_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_20_36137501_36162501_360C;SPAN=8439;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:134 GQ:39.8 PL:[39.8, 0.0, 284.0] SR:1 DR:23 LR:-39.62 LO:50.42);ALT=G[chr20:36156194[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	36322554	+	chr20	36361278	+	.	19	4	7001178_1	51.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7001178_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_36358001_36383001_172C;SPAN=38724;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:66 GQ:51.5 PL:[51.5, 0.0, 107.6] SR:4 DR:19 LR:-51.44 LO:52.57);ALT=G[chr20:36361278[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	36488746	+	chr20	36500326	+	.	0	14	7001542_1	18.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7001542_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_36480501_36505501_342C;SPAN=11580;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:103 GQ:18.5 PL:[18.5, 0.0, 229.7] SR:14 DR:0 LR:-18.31 LO:29.14);ALT=G[chr20:36500326[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	37055149	+	chr20	37059683	+	.	0	13	7003735_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=7003735_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_37044001_37069001_423C;SPAN=4534;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:134 GQ:6.8 PL:[6.8, 0.0, 317.0] SR:13 DR:0 LR:-6.609 LO:25.03);ALT=G[chr20:37059683[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	37059756	+	chr20	37063146	+	.	0	29	7003751_1	66.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=7003751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_37044001_37069001_258C;SPAN=3390;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:108 GQ:66.5 PL:[66.5, 0.0, 195.2] SR:29 DR:0 LR:-66.47 LO:70.01);ALT=C[chr20:37063146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	37059807	+	chr20	37063880	+	.	20	0	7003752_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7003752_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:37059807(+)-20:37063880(-)__20_37044001_37069001D;SPAN=4073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:103 GQ:38.3 PL:[38.3, 0.0, 209.9] SR:0 DR:20 LR:-38.12 LO:45.04);ALT=G[chr20:37063880[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	46130764	+	chr20	46211925	+	.	8	5	7036791_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7036791_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_46207001_46232001_248C;SPAN=81161;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:61 GQ:13.4 PL:[13.4, 0.0, 132.2] SR:5 DR:8 LR:-13.18 LO:19.08);ALT=G[chr20:46211925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	46131192	+	chr20	46250970	+	.	9	0	7036283_1	16.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=7036283_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:46131192(+)-20:46250970(-)__20_46231501_46256501D;SPAN=119778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:48 GQ:16.7 PL:[16.7, 0.0, 99.2] SR:0 DR:9 LR:-16.7 LO:20.11);ALT=G[chr20:46250970[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47643305	-	chr20	47644438	+	.	8	0	7041416_1	0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7041416_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:47643305(-)-20:47644438(-)__20_47628001_47653001D;SPAN=1133;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:105 GQ:1.8 PL:[0.0, 1.8, 257.4] SR:0 DR:8 LR:2.039 LO:14.52);ALT=[chr20:47644438[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	47770611	+	chr20	47804653	+	.	3	2	7042830_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7042830_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47799501_47824501_5C;SPAN=34042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:43 GQ:5 PL:[5.0, 0.0, 97.4] SR:2 DR:3 LR:-4.855 LO:10.04);ALT=G[chr20:47804653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47836079	+	chr20	47837987	+	.	48	17	7042751_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7042751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47824001_47849001_305C;SPAN=1908;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:127 GQ:99 PL:[143.9, 0.0, 163.7] SR:17 DR:48 LR:-143.8 LO:143.9);ALT=G[chr20:47837987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47853047	+	chr20	47855484	+	.	3	9	7042443_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7042443_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47848501_47873501_201C;SPAN=2437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:116 GQ:1.5 PL:[0.0, 1.5, 283.8] SR:9 DR:3 LR:1.718 LO:16.41);ALT=G[chr20:47855484[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47888289	+	chr20	47892315	+	.	4	2	7043022_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7043022_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47873001_47898001_387C;SPAN=4026;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:107 GQ:12.3 PL:[0.0, 12.3, 283.8] SR:2 DR:4 LR:12.48 LO:7.986);ALT=T[chr20:47892315[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47895263	+	chr20	47897021	+	.	43	0	7043046_1	87.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7043046_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:47895263(+)-20:47897021(-)__20_47873001_47898001D;SPAN=1758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:203 GQ:87.1 PL:[87.1, 0.0, 404.0] SR:0 DR:43 LR:-86.95 LO:98.67);ALT=C[chr20:47897021[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47895263	+	chr20	47897436	+	.	11	0	7043047_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7043047_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:47895263(+)-20:47897436(-)__20_47873001_47898001D;SPAN=2173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:11 DP:151 GQ:4.3 PL:[0.0, 4.3, 372.9] SR:0 DR:11 LR:4.599 LO:19.75);ALT=C[chr20:47897436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47895747	+	chr20	47897022	+	.	0	138	7043050_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GT;MAPQ=60;MATEID=7043050_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_47873001_47898001_86C;SPAN=1275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:138 DP:322 GQ:99 PL:[368.5, 0.0, 411.4] SR:138 DR:0 LR:-368.3 LO:368.4);ALT=T[chr20:47897022[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47897501	+	chr20	47905582	+	ATACAGGGTATGATACAGCATCCTACAAGAATGAGCAAACCTATTCTGATGGCAGGAGATTGAGGAC	5	13	7043061_1	32.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CAG;INSERTION=ATACAGGGTATGATACAGCATCCTACAAGAATGAGCAAACCTATTCTGATGGCAGGAGATTGAGGAC;MAPQ=60;MATEID=7043061_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_47873001_47898001_48C;SPAN=8081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:102 GQ:32 PL:[32.0, 0.0, 213.5] SR:13 DR:5 LR:-31.78 LO:39.7);ALT=G[chr20:47905582[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	47897501	+	chr20	47905580	+	.	5	57	7043060_1	99.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=7043060_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AA;SCTG=c_20_47873001_47898001_256C;SPAN=8079;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:102 GQ:68.3 PL:[177.2, 0.0, 68.3] SR:57 DR:5 LR:-179.5 LO:179.5);ALT=G[chr20:47905580[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48429486	+	chr20	48431545	+	.	10	9	7045348_1	17.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7045348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_48412001_48437001_382C;SPAN=2059;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:129 GQ:17.9 PL:[17.9, 0.0, 295.1] SR:9 DR:10 LR:-17.87 LO:32.62);ALT=G[chr20:48431545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48553089	+	chr20	48558098	+	.	0	28	7045902_1	60.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7045902_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_48534501_48559501_292C;SPAN=5009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:118 GQ:60.5 PL:[60.5, 0.0, 225.5] SR:28 DR:0 LR:-60.46 LO:65.83);ALT=T[chr20:48558098[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48562789	+	chr20	48565784	+	.	0	13	7045976_1	13.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7045976_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_48559001_48584001_293C;SPAN=2995;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:111 GQ:13.1 PL:[13.1, 0.0, 254.0] SR:13 DR:0 LR:-12.84 LO:26.15);ALT=T[chr20:48565784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48565893	+	chr20	48568612	+	.	0	15	7045991_1	18.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=7045991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_48559001_48584001_257C;SPAN=2719;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:115 GQ:18.5 PL:[18.5, 0.0, 259.4] SR:15 DR:0 LR:-18.36 LO:30.93);ALT=G[chr20:48568612[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48760199	+	chr20	48770144	+	.	13	0	7047090_1	16.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7047090_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:48760199(+)-20:48770144(-)__20_48755001_48780001D;SPAN=9945;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:99 GQ:16.1 PL:[16.1, 0.0, 224.0] SR:0 DR:13 LR:-16.09 LO:26.85);ALT=A[chr20:48770144[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48892927	+	chr20	48894026	+	.	10	4	7047197_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7047197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_48877501_48902501_127C;SPAN=1099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:114 GQ:2.3 PL:[2.3, 0.0, 272.9] SR:4 DR:10 LR:-2.125 LO:18.79);ALT=G[chr20:48894026[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	48892956	+	chr20	48894712	+	.	22	0	7047199_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7047199_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:48892956(+)-20:48894712(-)__20_48877501_48902501D;SPAN=1756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:111 GQ:42.8 PL:[42.8, 0.0, 224.3] SR:0 DR:22 LR:-42.55 LO:49.76);ALT=T[chr20:48894712[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	49127071	+	chr20	49177897	+	.	11	0	7048522_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7048522_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:49127071(+)-20:49177897(-)__20_49171501_49196501D;SPAN=50826;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:59 GQ:20.3 PL:[20.3, 0.0, 122.6] SR:0 DR:11 LR:-20.33 LO:24.55);ALT=A[chr20:49177897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	49127128	+	chr20	49184914	+	ATATCCGACATGAAGCCAGTGACTTCCCATGTAGAGTGGCCAAGCTTCCTAAGAACAAAAACCGAAATAGGTACAGAGACGTCAGTCCCTTTGACCATAGTCGGATTAAACTACATCAAGAAGATAATGACTATATCAACGCTAGTTTGATAAAAATGGAAGAAGCCCAAAGGAGTTACATTCTTACC	0	22	7048524_1	58.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=ATATCCGACATGAAGCCAGTGACTTCCCATGTAGAGTGGCCAAGCTTCCTAAGAACAAAAACCGAAATAGGTACAGAGACGTCAGTCCCTTTGACCATAGTCGGATTAAACTACATCAAGAAGATAATGACTATATCAACGCTAGTTTGATAAAAATGGAAGAAGCCCAAAGGAGTTACATTCTTACC;MAPQ=60;MATEID=7048524_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_49171501_49196501_369C;SPAN=57786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:52 GQ:58.7 PL:[58.7, 0.0, 65.3] SR:22 DR:0 LR:-58.53 LO:58.57);ALT=G[chr20:49184914[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	49127128	+	chr20	49181506	+	ATATCCGACATGAAGCCAGTGACTTCCCATGTAGAGTGGCCAAGCTTCCTAAGAACAAAAACCGAAATAGGTACAGAGACGTCAGTCCCT	0	25	7048208_1	60.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=ATATCCGACATGAAGCCAGTGACTTCCCATGTAGAGTGGCCAAGCTTCCTAAGAACAAAAACCGAAATAGGTACAGAGACGTCAGTCCCT;MAPQ=60;MATEID=7048208_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_49122501_49147501_211C;SPAN=54378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:81 GQ:60.8 PL:[60.8, 0.0, 133.4] SR:25 DR:0 LR:-60.58 LO:62.17);ALT=G[chr20:49181506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	49571871	+	chr20	49575008	+	.	10	0	7050115_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7050115_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:49571871(+)-20:49575008(-)__20_49563501_49588501D;SPAN=3137;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:101 GQ:5.9 PL:[5.9, 0.0, 236.9] SR:0 DR:10 LR:-5.647 LO:19.35);ALT=T[chr20:49575008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	52233413	-	chr20	52234937	+	.	8	0	7060239_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7060239_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:52233413(-)-20:52234937(-)__20_52209501_52234501D;SPAN=1524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:50 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:0 DR:8 LR:-12.86 LO:17.27);ALT=[chr20:52234937[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	52689060	+	chr20	52687447	+	.	2	4	7062355_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7062355_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_52675001_52700001_262C;SPAN=1613;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:113 GQ:17.1 PL:[0.0, 17.1, 306.9] SR:4 DR:2 LR:17.41 LO:5.901);ALT=]chr20:52689060]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	52830997	+	chr20	52835556	+	AAACAACTCCAAAACCTAGAAGATGCTTGTGATGACATCATGCTTGCAGATGATGATTGCTTAATGATACCTTATCAAATTGGTGATGTCTTCATTAGCCATTCTCAAGAAGAAACGCAAGAAATGTTAGAAGAAGCAA	3	39	7062915_1	99.0	.	DISC_MAPQ=32;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AAACAACTCCAAAACCTAGAAGATGCTTGTGATGACATCATGCTTGCAGATGATGATTGCTTAATGATACCTTATCAAATTGGTGATGTCTTCATTAGCCATTCTCAAGAAGAAACGCAAGAAATGTTAGAAGAAGCAA;MAPQ=60;MATEID=7062915_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_52822001_52847001_5C;SPAN=4559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:75 GQ:68.9 PL:[111.8, 0.0, 68.9] SR:39 DR:3 LR:-112.2 LO:112.2);ALT=G[chr20:52835556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	52831979	+	chr20	52835556	+	.	3	20	7062917_1	52.0	.	DISC_MAPQ=40;EVDNC=TSI_L;HOMSEQ=AG;MAPQ=60;MATEID=7062917_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=AAAA;SCTG=c_20_52822001_52847001_5C;SPAN=3577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:87 GQ:52.4 PL:[52.4, 0.0, 158.0] SR:20 DR:3 LR:-52.35 LO:55.34);ALT=G[chr20:52835556[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	53699589	-	chr20	53700625	+	.	9	0	7065825_1	2.0	.	DISC_MAPQ=35;EVDNC=DSCRD;IMPRECISE;MAPQ=35;MATEID=7065825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:53699589(-)-20:53700625(-)__20_53679501_53704501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:99 GQ:2.9 PL:[2.9, 0.0, 237.2] SR:0 DR:9 LR:-2.887 LO:17.06);ALT=[chr20:53700625[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr20	54434623	+	chr20	54440617	+	.	66	46	7068164_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AATAAATTTGTGG;MAPQ=60;MATEID=7068164_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_20_54439001_54464001_8C;SPAN=5994;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:66 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:46 DR:66 LR:-260.8 LO:260.8);ALT=G[chr20:54440617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	54934248	+	chr20	54940140	+	.	0	24	7069404_1	51.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=7069404_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_54929001_54954001_300C;SPAN=5892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:104 GQ:51.2 PL:[51.2, 0.0, 199.7] SR:24 DR:0 LR:-51.05 LO:56.09);ALT=G[chr20:54940140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55043823	+	chr20	55045653	+	.	4	2	7069982_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=7069982_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_55027001_55052001_310C;SPAN=1830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:130 GQ:15.3 PL:[0.0, 15.3, 346.5] SR:2 DR:4 LR:15.41 LO:9.551);ALT=G[chr20:55045653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55043825	+	chr20	55048355	+	.	27	6	7069983_1	67.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AGGTC;MAPQ=60;MATEID=7069983_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_55027001_55052001_333C;SPAN=4530;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:130 GQ:67.1 PL:[67.1, 0.0, 248.6] SR:6 DR:27 LR:-67.11 LO:72.97);ALT=C[chr20:55048355[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55043829	+	chr20	55049727	+	.	53	0	7069985_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7069985_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:55043829(+)-20:55049727(-)__20_55027001_55052001D;SPAN=5898;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:132 GQ:99 PL:[139.4, 0.0, 179.0] SR:0 DR:53 LR:-139.2 LO:139.5);ALT=G[chr20:55049727[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55043831	+	chr20	55052038	+	.	12	0	7070107_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7070107_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:55043831(+)-20:55052038(-)__20_55051501_55076501D;SPAN=8207;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:66 GQ:21.8 PL:[21.8, 0.0, 137.3] SR:0 DR:12 LR:-21.73 LO:26.64);ALT=T[chr20:55052038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55048451	+	chr20	55049730	+	.	0	50	7070001_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=7070001_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_55027001_55052001_114C;SPAN=1279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:123 GQ:99 PL:[131.9, 0.0, 164.9] SR:50 DR:0 LR:-131.7 LO:132.0);ALT=G[chr20:55049730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55049827	+	chr20	55052039	+	.	2	35	7070108_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7070108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_55051501_55076501_150C;SPAN=2212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:66 GQ:54.8 PL:[104.3, 0.0, 54.8] SR:35 DR:2 LR:-105.0 LO:105.0);ALT=G[chr20:55052039[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	55052183	+	chr20	55059164	+	.	0	14	7070114_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CAGGTT;MAPQ=60;MATEID=7070114_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_55051501_55076501_220C;SPAN=6981;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:127 GQ:11.9 PL:[11.9, 0.0, 295.7] SR:14 DR:0 LR:-11.81 LO:27.77);ALT=T[chr20:55059164[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	23852644	+	chr20	55239234	+	.	21	58	7236357_1	99.0	.	DISC_MAPQ=20;EVDNC=ASDIS;HOMSEQ=TGGTGCAATCTCGGCTCACTGCAACCTCTG;MAPQ=33;MATEID=7236357_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_23838501_23863501_229C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:75 DP:43 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:58 DR:21 LR:-221.2 LO:221.2);ALT=]chr22:23852644]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr20	60712007	+	chr20	60714130	+	TGAGGGATTGATCTCGCCTCATGACAGCAAGTTCAATGTTTTTGCCACCTGACTGAACCACTTCCAGGAGTGCCTTGATCACCAGCTTAATGGTCAGATCATCTGTTTCAATGGCTTCGTCAGTATAGTTCTTCTCCAGGAACTCACGCACTGACTTGGCACCCCGGCCTATGGCATTGG	0	190	7089926_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CCT;INSERTION=TGAGGGATTGATCTCGCCTCATGACAGCAAGTTCAATGTTTTTGCCACCTGACTGAACCACTTCCAGGAGTGCCTTGATCACCAGCTTAATGGTCAGATCATCTGTTTCAATGGCTTCGTCAGTATAGTTCTTCTCCAGGAACTCACGCACTGACTTGGCACCCCGGCCTATGGCATTGG;MAPQ=60;MATEID=7089926_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_20_60711001_60736001_54C;SPAN=2123;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:190 DP:185 GQ:51.4 PL:[564.4, 51.4, 0.0] SR:190 DR:0 LR:-564.4 LO:564.4);ALT=T[chr20:60714130[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	60712050	+	chr20	60713224	+	.	10	0	7089927_1	0	.	DISC_MAPQ=36;EVDNC=DSCRD;IMPRECISE;MAPQ=36;MATEID=7089927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:60712050(+)-20:60713224(-)__20_60711001_60736001D;SPAN=1174;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:158 GQ:9.7 PL:[0.0, 9.7, 402.6] SR:0 DR:10 LR:9.796 LO:17.32);ALT=A[chr20:60713224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	60714967	+	chr20	60718262	+	AGGCCATGCAGACGTTGTCATCCAAAGCACAGATCTTCCGCACTGTTCTTTCATCCTGCAGTTTGGCCACTGACTTCTTCTCCACACCAAGAACAACAATGTCTCTTCCTCGAACACCA	91	133	7089945_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=ACC;INSERTION=AGGCCATGCAGACGTTGTCATCCAAAGCACAGATCTTCCGCACTGTTCTTTCATCCTGCAGTTTGGCCACTGACTTCTTCTCCACACCAAGAACAACAATGTCTCTTCCTCGAACACCA;MAPQ=60;MATEID=7089945_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_20_60711001_60736001_226C;SPAN=3295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:179 DP:153 GQ:48.4 PL:[531.4, 48.4, 0.0] SR:133 DR:91 LR:-531.4 LO:531.4);ALT=A[chr20:60718262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	60716001	+	chr20	60718262	+	.	118	39	7089949_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=ACC;MAPQ=60;MATEID=7089949_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_20_60711001_60736001_226C;SPAN=2261;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:129 DP:142 GQ:38.2 PL:[419.2, 38.2, 0.0] SR:39 DR:118 LR:-419.2 LO:419.2);ALT=C[chr20:60718262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	61177144	+	chr20	61176057	+	.	29	0	7091746_1	77.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7091746_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:61176057(-)-20:61177144(+)__20_61176501_61201501D;SPAN=1087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:67 GQ:77.6 PL:[77.6, 0.0, 84.2] SR:0 DR:29 LR:-77.58 LO:77.6);ALT=]chr20:61177144]C;VARTYPE=BND:DUP-th;JOINTYPE=th
chr20	61436382	+	chr20	61438885	+	.	0	7	7092292_1	0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=7092292_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_61421501_61446501_369C;SPAN=2503;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:91 GQ:1.2 PL:[0.0, 1.2, 221.1] SR:7 DR:0 LR:1.547 LO:12.74);ALT=G[chr20:61438885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	61569605	+	chr20	61572842	+	.	13	10	7092810_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7092810_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_61568501_61593501_179C;SPAN=3237;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:73 GQ:39.8 PL:[39.8, 0.0, 135.5] SR:10 DR:13 LR:-39.64 LO:42.67);ALT=G[chr20:61572842[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	61572972	+	chr20	61574336	+	.	0	5	7092821_1	0	.	EVDNC=ASSMB;HOMSEQ=CAG;MAPQ=60;MATEID=7092821_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_61568501_61593501_332C;SPAN=1364;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:88 GQ:7.2 PL:[0.0, 7.2, 227.7] SR:5 DR:0 LR:7.336 LO:8.42);ALT=G[chr20:61574336[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	61584242	+	chr20	61588114	+	.	13	9	7092849_1	38.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=7092849_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_61568501_61593501_162C;SPAN=3872;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:77 GQ:38.6 PL:[38.6, 0.0, 147.5] SR:9 DR:13 LR:-38.56 LO:42.19);ALT=G[chr20:61588114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62275331	+	chr20	62284682	+	.	14	0	7095429_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7095429_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62275331(+)-20:62284682(-)__20_62279001_62304001D;SPAN=9351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:21 GQ:7.7 PL:[40.7, 0.0, 7.7] SR:0 DR:14 LR:-41.52 LO:41.52);ALT=T[chr20:62284682[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62275663	+	chr20	62284680	+	.	9	3	7095430_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7095430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62279001_62304001_16C;SPAN=9017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:21 GQ:20.9 PL:[27.5, 0.0, 20.9] SR:3 DR:9 LR:-27.33 LO:27.33);ALT=C[chr20:62284680[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62368115	+	chr20	62369170	+	.	25	0	7095633_1	58.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7095633_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62368115(+)-20:62369170(-)__20_62352501_62377501D;SPAN=1055;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:90 GQ:58.1 PL:[58.1, 0.0, 160.4] SR:0 DR:25 LR:-58.14 LO:60.79);ALT=G[chr20:62369170[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62496737	+	chr20	62500647	+	.	13	2	7096223_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7096223_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62499501_62524501_292C;SPAN=3910;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:51 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:2 DR:13 LR:-32.4 LO:33.96);ALT=G[chr20:62500647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62496765	+	chr20	62505018	+	.	12	0	7096224_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7096224_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62496765(+)-20:62505018(-)__20_62499501_62524501D;SPAN=8253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:55 GQ:24.8 PL:[24.8, 0.0, 107.3] SR:0 DR:12 LR:-24.71 LO:27.71);ALT=G[chr20:62505018[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62500797	+	chr20	62505019	+	.	2	10	7096231_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTG;MAPQ=60;MATEID=7096231_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62499501_62524501_21C;SPAN=4222;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:10 DR:2 LR:-7.051 LO:21.42);ALT=G[chr20:62505019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62577997	+	chr20	62587613	+	.	0	12	7096078_1	15.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7096078_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62573001_62598001_350C;SPAN=9616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:91 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:12 DR:0 LR:-14.96 LO:24.81);ALT=C[chr20:62587613[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62596231	+	chr20	62597441	+	.	41	0	7096127_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7096127_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62596231(+)-20:62597441(-)__20_62573001_62598001D;SPAN=1210;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:59 GQ:23.6 PL:[119.3, 0.0, 23.6] SR:0 DR:41 LR:-123.0 LO:123.0);ALT=G[chr20:62597441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62612669	+	chr20	62614399	+	.	42	36	7096555_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7096555_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62597501_62622501_283C;SPAN=1730;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:60 DP:113 GQ:99 PL:[167.6, 0.0, 104.9] SR:36 DR:42 LR:-168.2 LO:168.2);ALT=G[chr20:62614399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62614568	+	chr20	62616258	+	.	2	15	7096566_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7096566_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62597501_62622501_388C;SPAN=1690;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:94 GQ:27.5 PL:[27.5, 0.0, 199.1] SR:15 DR:2 LR:-27.35 LO:35.01);ALT=G[chr20:62616258[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62701991	+	chr20	62703218	+	.	0	4	7096707_1	0	.	EVDNC=ASSMB;HOMSEQ=CACAGGTG;MAPQ=60;MATEID=7096707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62695501_62720501_115C;SPAN=1227;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:76 GQ:7.2 PL:[0.0, 7.2, 198.0] SR:4 DR:0 LR:7.386 LO:6.6);ALT=G[chr20:62703218[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62705895	+	chr20	62707877	+	.	5	11	7096722_1	14.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=7096722_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CC;SCTG=c_20_62695501_62720501_108C;SPAN=1982;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:119 GQ:14 PL:[14.0, 0.0, 274.7] SR:11 DR:5 LR:-13.97 LO:28.2);ALT=C[chr20:62707877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62705947	+	chr20	62711224	+	.	9	0	7096723_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7096723_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62705947(+)-20:62711224(-)__20_62695501_62720501D;SPAN=5277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:0 DR:9 LR:-12.1 LO:18.81);ALT=A[chr20:62711224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62708042	+	chr20	62711225	+	.	11	0	7096732_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7096732_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=20:62708042(+)-20:62711225(-)__20_62695501_62720501D;SPAN=3183;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=A[chr20:62711225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr20	62708308	+	chr20	62710647	+	.	0	14	7096736_1	26.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7096736_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_20_62695501_62720501_233C;SPAN=2339;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:73 GQ:26.6 PL:[26.6, 0.0, 148.7] SR:14 DR:0 LR:-26.44 LO:31.44);ALT=C[chr20:62710647[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30397103	+	chr21	30400190	+	.	16	0	7151843_1	33.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7151843_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:30397103(+)-21:30400190(-)__21_30380001_30405001D;SPAN=3087;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:72 GQ:33.5 PL:[33.5, 0.0, 139.1] SR:0 DR:16 LR:-33.31 LO:37.09);ALT=G[chr21:30400190[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30397120	+	chr21	30402912	+	.	9	0	7151844_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7151844_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:30397120(+)-21:30402912(-)__21_30380001_30405001D;SPAN=5792;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:64 GQ:12.5 PL:[12.5, 0.0, 141.2] SR:0 DR:9 LR:-12.37 LO:18.88);ALT=T[chr21:30402912[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30400295	+	chr21	30402913	+	.	0	12	7151851_1	21.0	.	EVDNC=ASSMB;HOMSEQ=TAG;MAPQ=60;MATEID=7151851_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_30380001_30405001_163C;SPAN=2618;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:67 GQ:21.5 PL:[21.5, 0.0, 140.3] SR:12 DR:0 LR:-21.46 LO:26.55);ALT=G[chr21:30402913[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30440031	+	chr21	30445871	+	.	17	0	7151205_1	37.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7151205_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:30440031(+)-21:30445871(-)__21_30429001_30454001D;SPAN=5840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:69 GQ:37.4 PL:[37.4, 0.0, 129.8] SR:0 DR:17 LR:-37.42 LO:40.29);ALT=T[chr21:30445871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30441881	+	chr21	30445874	+	.	27	0	7151207_1	72.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7151207_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:30441881(+)-21:30445874(-)__21_30429001_30454001D;SPAN=3993;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:63 GQ:72.2 PL:[72.2, 0.0, 78.8] SR:0 DR:27 LR:-72.06 LO:72.09);ALT=C[chr21:30445874[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30671330	+	chr21	30693541	+	.	13	0	7151916_1	26.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7151916_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:30671330(+)-21:30693541(-)__21_30674001_30699001D;SPAN=22211;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:60 GQ:26.6 PL:[26.6, 0.0, 119.0] SR:0 DR:13 LR:-26.66 LO:29.98);ALT=G[chr21:30693541[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	30677645	+	chr21	30693542	+	.	5	9	7151923_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GT;MAPQ=60;MATEID=7151923_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_30674001_30699001_328C;SPAN=15897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:9 DR:5 LR:-11.39 LO:22.24);ALT=T[chr21:30693542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	39817576	+	chr21	39870302	+	.	19	0	7176812_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7176812_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:39817576(+)-21:39870302(-)__21_39861501_39886501D;SPAN=52726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:27 GQ:9.2 PL:[55.4, 0.0, 9.2] SR:0 DR:19 LR:-57.18 LO:57.18);ALT=C[chr21:39870302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40178044	+	chr21	40181958	+	.	0	18	7177472_1	48.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7177472_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40180001_40205001_3C;SPAN=3914;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:41 GQ:48.5 PL:[48.5, 0.0, 48.5] SR:18 DR:0 LR:-48.31 LO:48.32);ALT=G[chr21:40181958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40178051	+	chr21	40184924	+	.	16	0	7177473_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7177473_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:40178051(+)-21:40184924(-)__21_40180001_40205001D;SPAN=6873;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:45 GQ:40.7 PL:[40.7, 0.0, 67.1] SR:0 DR:16 LR:-40.62 LO:41.02);ALT=G[chr21:40184924[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40182030	+	chr21	40184925	+	.	0	20	7177483_1	42.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7177483_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40180001_40205001_303C;SPAN=2895;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:88 GQ:42.2 PL:[42.2, 0.0, 170.9] SR:20 DR:0 LR:-42.18 LO:46.59);ALT=G[chr21:40184925[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40185038	+	chr21	40186705	+	ACTCCGCCAACTGTGAATTGCCTTTGTTAACCCCGTGCAGCAAGGCTGTGATGAGTCAAGCCTTAAAAGCTACCTTCAGTGGCTTCAAAAAGGAACAGCGGCGCCTGGGCATTCCAAAGA	0	23	7177492_1	54.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ACTCCGCCAACTGTGAATTGCCTTTGTTAACCCCGTGCAGCAAGGCTGTGATGAGTCAAGCCTTAAAAGCTACCTTCAGTGGCTTCAAAAAGGAACAGCGGCGCCTGGGCATTCCAAAGA;MAPQ=60;MATEID=7177492_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_21_40180001_40205001_82C;SPAN=1667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:79 GQ:54.5 PL:[54.5, 0.0, 137.0] SR:23 DR:0 LR:-54.52 LO:56.49);ALT=G[chr21:40186705[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40383249	+	chr21	40386577	+	.	35	2	7178258_1	95.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=7178258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40376001_40401001_274C;SPAN=3328;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:88 GQ:95 PL:[95.0, 0.0, 118.1] SR:2 DR:35 LR:-95.0 LO:95.14);ALT=G[chr21:40386577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40547592	+	chr21	40549361	+	.	0	23	7178586_1	59.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7178586_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_21_40523001_40548001_101C;SPAN=1769;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:60 GQ:59.6 PL:[59.6, 0.0, 86.0] SR:23 DR:0 LR:-59.67 LO:59.93);ALT=T[chr21:40549361[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40552391	+	chr21	40555282	+	.	8	0	7178477_1	3.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7178477_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:40552391(+)-21:40555282(-)__21_40547501_40572501D;SPAN=2891;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:84 GQ:3.8 PL:[3.8, 0.0, 198.5] SR:0 DR:8 LR:-3.65 LO:15.33);ALT=G[chr21:40555282[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40553806	+	chr21	40555177	+	.	0	17	7178486_1	27.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7178486_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_21_40547501_40572501_315C;SPAN=1371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:107 GQ:27.2 PL:[27.2, 0.0, 231.8] SR:17 DR:0 LR:-27.13 LO:36.64);ALT=T[chr21:40555177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40717204	+	chr21	40720902	+	.	19	0	7179002_1	43.0	.	DISC_MAPQ=26;EVDNC=DSCRD;IMPRECISE;MAPQ=26;MATEID=7179002_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:40717204(+)-21:40720902(-)__21_40719001_40744001D;SPAN=3698;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:73 GQ:43.1 PL:[43.1, 0.0, 132.2] SR:0 DR:19 LR:-42.94 LO:45.56);ALT=T[chr21:40720902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr21	40752475	+	chr21	40762623	+	.	16	0	7179101_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7179101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=21:40752475(+)-21:40762623(-)__21_40743501_40768501D;SPAN=10148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:102 GQ:25.4 PL:[25.4, 0.0, 220.1] SR:0 DR:16 LR:-25.18 LO:34.39);ALT=T[chr21:40762623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	16862336	+	chr22	16855969	+	.	9	0	7205179_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7205179_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:16855969(-)-22:16862336(+)__22_16856001_16881001D;SPAN=6367;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:175 GQ:17.5 PL:[0.0, 17.5, 458.8] SR:0 DR:9 LR:17.7 LO:14.76);ALT=]chr22:16862336]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	17004009	+	chr22	17033723	+	TTTTT	15	16	7207082_1	66.0	.	DISC_MAPQ=17;EVDNC=ASDIS;INSERTION=TTTTT;MAPQ=0;MATEID=7207082_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_17027501_17052501_304C;SPAN=29714;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:34 GQ:14 PL:[66.8, 0.0, 14.0] SR:16 DR:15 LR:-68.47 LO:68.47);ALT=A[chr22:17033723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	17630662	+	chr22	17640082	+	.	10	0	7208145_1	20.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7208145_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:17630662(+)-22:17640082(-)__22_17640001_17665001D;SPAN=9420;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:45 GQ:20.9 PL:[20.9, 0.0, 86.9] SR:0 DR:10 LR:-20.82 LO:23.18);ALT=G[chr22:17640082[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	17770350	+	chr22	17779109	+	C	88	83	7208307_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=C;MAPQ=60;MATEID=7208307_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_17762501_17787501_215C;SPAN=8759;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:144 DP:32 GQ:38.8 PL:[425.8, 38.8, 0.0] SR:83 DR:88 LR:-425.8 LO:425.8);ALT=C[chr22:17779109[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18057770	+	chr22	18060458	+	.	91	18	7210196_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=ATTCTCCTGCCTCAGCCTCC;MAPQ=60;MATEID=7210196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18032001_18057001_398C;SPAN=2688;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:105 DP:0 GQ:28.2 PL:[310.2, 28.2, 0.0] SR:18 DR:91 LR:-310.3 LO:310.3);ALT=C[chr22:18060458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18075505	+	chr22	18077295	+	.	3	3	7209962_1	0	.	DISC_MAPQ=45;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=0;MATEID=7209962_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18056501_18081501_328C;SECONDARY;SPAN=1790;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:108 GQ:9.3 PL:[0.0, 9.3, 280.5] SR:3 DR:3 LR:9.454 LO:10.04);ALT=G[chr22:18077295[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18121654	+	chr22	18138426	+	.	29	6	7210606_1	86.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=7210606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18130001_18155001_149C;SPAN=16772;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:45 GQ:20.9 PL:[86.9, 0.0, 20.9] SR:6 DR:29 LR:-88.96 LO:88.96);ALT=T[chr22:18138426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18178976	+	chr22	18185006	+	.	0	9	7210744_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AAG;MAPQ=60;MATEID=7210744_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18179001_18204001_67C;SPAN=6030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:83 GQ:7.4 PL:[7.4, 0.0, 192.2] SR:9 DR:0 LR:-7.222 LO:17.79);ALT=G[chr22:18185006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18218357	+	chr22	18220782	+	.	2	35	7210991_1	89.0	.	DISC_MAPQ=37;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7210991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18203501_18228501_327C;SPAN=2425;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:119 GQ:89.9 PL:[89.9, 0.0, 198.8] SR:35 DR:2 LR:-89.9 LO:92.16);ALT=C[chr22:18220782[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18220997	+	chr22	18222114	+	.	3	6	7211009_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7211009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18203501_18228501_229C;SPAN=1117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:122 GQ:3 PL:[0.0, 3.0, 300.3] SR:6 DR:3 LR:3.344 LO:16.21);ALT=T[chr22:18222114[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18221041	+	chr22	18257146	+	.	9	0	7211010_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7211010_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:18221041(+)-22:18257146(-)__22_18203501_18228501D;SPAN=36105;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:44 GQ:17.9 PL:[17.9, 0.0, 87.2] SR:0 DR:9 LR:-17.79 LO:20.5);ALT=T[chr22:18257146[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18226781	+	chr22	18232867	+	.	0	20	7211226_1	49.0	.	EVDNC=ASSMB;HOMSEQ=TGACCT;MAPQ=60;MATEID=7211226_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18228001_18253001_382C;SPAN=6086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:60 GQ:49.7 PL:[49.7, 0.0, 95.9] SR:20 DR:0 LR:-49.76 LO:50.57);ALT=T[chr22:18232867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18226825	+	chr22	18257142	+	.	55	0	7211033_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7211033_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:18226825(+)-22:18257142(-)__22_18203501_18228501D;SPAN=30317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:55 DP:66 GQ:4.5 PL:[168.3, 4.5, 0.0] SR:0 DR:55 LR:-174.7 LO:174.7);ALT=G[chr22:18257142[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18232941	+	chr22	18257145	+	.	8	6	7211249_1	20.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=7211249_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18228001_18253001_109C;SPAN=24204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:58 GQ:20.6 PL:[20.6, 0.0, 119.6] SR:6 DR:8 LR:-20.6 LO:24.64);ALT=C[chr22:18257145[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	18918714	+	chr22	18923528	+	.	0	9	7214317_1	3.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7214317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_18914001_18939001_240C;SPAN=4814;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:97 GQ:3.5 PL:[3.5, 0.0, 231.2] SR:9 DR:0 LR:-3.429 LO:17.14);ALT=G[chr22:18923528[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19420131	+	chr22	19422257	+	CTTCTGGGAACTTGGCAGACGCAGCTTAGAGAGACTCACCAGCGAGCGTCATTGTTGTCTTTCTGGGAACTCATTCCCATG	33	28	7216473_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CTTCTGGGAACTTGGCAGACGCAGCTTAGAGAGACTCACCAGCGAGCGTCATTGTTGTCTTTCTGGGAACTCATTCCCATG;MAPQ=60;MATEID=7216473_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_19404001_19429001_151C;SPAN=2126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:112 GQ:99 PL:[128.3, 0.0, 141.5] SR:28 DR:33 LR:-128.1 LO:128.2);ALT=G[chr22:19422257[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19429220	+	chr22	19434897	+	.	19	30	7216614_1	94.0	.	DISC_MAPQ=48;EVDNC=ASDIS;HOMSEQ=GCACCTG;MAPQ=60;MATEID=7216614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19428501_19453501_39C;SPAN=5677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:127 GQ:94.4 PL:[94.4, 0.0, 213.2] SR:30 DR:19 LR:-94.33 LO:96.89);ALT=G[chr22:19434897[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19463126	+	chr22	19466606	+	.	14	6	7216553_1	21.0	.	DISC_MAPQ=40;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7216553_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19453001_19478001_280C;SPAN=3480;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:127 GQ:21.8 PL:[21.8, 0.0, 285.8] SR:6 DR:14 LR:-21.71 LO:35.26);ALT=C[chr22:19466606[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19907171	+	chr22	19929270	+	.	15	0	7218913_1	37.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7218913_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:19907171(+)-22:19929270(-)__22_19894001_19919001D;SPAN=22099;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:46 GQ:37.1 PL:[37.1, 0.0, 73.4] SR:0 DR:15 LR:-37.05 LO:37.75);ALT=A[chr22:19929270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19929420	+	chr22	19948720	+	.	43	21	7218375_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7218375_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19918501_19943501_29C;SPAN=19300;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:21 DR:43 LR:-158.4 LO:158.4);ALT=G[chr22:19948720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19948812	+	chr22	19950048	+	.	42	72	7218265_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7218265_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19943001_19968001_172C;SPAN=1236;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:108 DP:119 GQ:32.1 PL:[353.1, 32.1, 0.0] SR:72 DR:42 LR:-353.2 LO:353.2);ALT=G[chr22:19950048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	19951815	+	chr22	19956057	+	TTTGG	10	5	7218272_1	14.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=TTTGG;MAPQ=60;MATEID=7218272_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_19943001_19968001_210C;SPAN=4242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:107 GQ:14 PL:[14.0, 0.0, 245.0] SR:5 DR:10 LR:-13.92 LO:26.38);ALT=T[chr22:19956057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20024378	+	chr22	20030875	+	.	3	5	7218603_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGG;MAPQ=60;MATEID=7218603_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_20016501_20041501_176C;SPAN=6497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:117 GQ:5.1 PL:[0.0, 5.1, 293.7] SR:5 DR:3 LR:5.29 LO:14.13);ALT=G[chr22:20030875[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20030967	+	chr22	20039987	+	.	0	11	7218637_1	9.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=7218637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_20016501_20041501_76C;SPAN=9020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:98 GQ:9.8 PL:[9.8, 0.0, 227.6] SR:11 DR:0 LR:-9.76 LO:21.91);ALT=G[chr22:20039987[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20105163	+	chr22	20109786	+	.	15	0	7219104_1	20.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7219104_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:20105163(+)-22:20109786(-)__22_20090001_20115001D;SPAN=4623;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:108 GQ:20.3 PL:[20.3, 0.0, 241.4] SR:0 DR:15 LR:-20.26 LO:31.37);ALT=C[chr22:20109786[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20105351	+	chr22	20106529	+	.	52	0	7219105_1	99.0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7219105_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:20105351(+)-22:20106529(-)__22_20090001_20115001D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:86 GQ:59.3 PL:[148.4, 0.0, 59.3] SR:0 DR:52 LR:-150.4 LO:150.4);ALT=G[chr22:20106529[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20151776	-	chr22	20152807	+	.	13	41	7219372_1	81.0	.	DISC_MAPQ=255;EVDNC=ASDIS;MAPQ=60;MATEID=7219372_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_22_20139001_20164001_235C;SPAN=1031;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:48 DP:286 GQ:81.1 PL:[81.1, 0.0, 612.5] SR:41 DR:13 LR:-80.96 LO:104.7);ALT=[chr22:20152807[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	20188935	-	chr22	48513210	+	GAGAGAAGGAAGGGAGGGAG	3	45	7219666_1	99.0	.	DISC_MAPQ=5;EVDNC=ASDIS;INSERTION=GAGAGAAGGAAGGGAGGGAG;MAPQ=26;MATEID=7219666_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_20188001_20213001_96C;SPAN=28324275;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:47 DP:30 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:45 DR:3 LR:-138.6 LO:138.6);ALT=[chr22:48513210[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	20862033	+	chr22	20891404	+	.	10	6	7222467_1	23.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=7222467_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_20849501_20874501_16C;SPAN=29371;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:62 GQ:23 PL:[23.0, 0.0, 125.3] SR:6 DR:10 LR:-22.81 LO:27.0);ALT=T[chr22:20891404[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	20950623	+	chr22	20953840	+	.	54	41	7222288_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7222288_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_20947501_20972501_293C;SPAN=3217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:82 DP:75 GQ:21.9 PL:[240.9, 21.9, 0.0] SR:41 DR:54 LR:-241.0 LO:241.0);ALT=C[chr22:20953840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	21213636	+	chr22	21224623	+	.	8	17	7224339_1	36.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7224339_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_21217001_21242001_295C;SPAN=10987;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:74 GQ:36.2 PL:[36.2, 0.0, 141.8] SR:17 DR:8 LR:-36.07 LO:39.69);ALT=G[chr22:21224623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	22652609	+	chr22	22658305	+	.	13	0	7231873_1	17.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7231873_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:22652609(+)-22:22658305(-)__22_22638001_22663001D;SPAN=5696;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:96 GQ:17 PL:[17.0, 0.0, 215.0] SR:0 DR:13 LR:-16.9 LO:27.04);ALT=G[chr22:22658305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	23478432	+	chr22	23479635	+	.	24	0	7234468_1	59.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7234468_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:23478432(+)-22:23479635(-)__22_23471001_23496001D;SPAN=1203;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:75 GQ:59 PL:[59.0, 0.0, 121.7] SR:0 DR:24 LR:-58.91 LO:60.15);ALT=C[chr22:23479635[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	23917275	+	chr22	23922172	+	.	0	12	7236132_1	6.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=34;MATEID=7236132_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_23912001_23937001_405C;SPAN=4897;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:122 GQ:6.8 PL:[6.8, 0.0, 287.3] SR:12 DR:0 LR:-6.559 LO:23.18);ALT=G[chr22:23922172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24108465	+	chr22	24109560	+	.	5	15	7236743_1	35.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=7236743_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_24108001_24133001_123C;SPAN=1095;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:101 GQ:35.6 PL:[35.6, 0.0, 207.2] SR:15 DR:5 LR:-35.36 LO:42.49);ALT=G[chr22:24109560[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24108516	+	chr22	24110032	+	.	10	0	7236947_1	20.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7236947_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:24108516(+)-22:24110032(-)__22_24083501_24108501D;SPAN=1516;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:46 GQ:20.6 PL:[20.6, 0.0, 89.9] SR:0 DR:10 LR:-20.55 LO:23.07);ALT=G[chr22:24110032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24129451	+	chr22	24133941	+	.	0	43	7237243_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=7237243_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24132501_24157501_376C;SPAN=4490;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:57 GQ:11 PL:[126.5, 0.0, 11.0] SR:43 DR:0 LR:-132.1 LO:132.1);ALT=T[chr22:24133941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24135876	+	chr22	24143125	+	.	2	5	7237257_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTCAGG;MAPQ=60;MATEID=7237257_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24132501_24157501_122C;SPAN=7249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:115 GQ:7.8 PL:[0.0, 7.8, 293.7] SR:5 DR:2 LR:8.049 LO:12.0);ALT=G[chr22:24143125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24195941	+	chr22	24198506	+	.	44	51	7237519_1	99.0	.	DISC_MAPQ=50;EVDNC=ASDIS;HOMSEQ=GAAAAAAA;MAPQ=60;MATEID=7237519_2;MATENM=1;NM=2;NUMPARTS=2;SCTG=c_22_24181501_24206501_422C;SPAN=2565;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:80 DP:72 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:51 DR:44 LR:-237.7 LO:237.7);ALT=A[chr22:24198506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24254525	-	chr22	24256334	+	.	14	0	7237445_1	30.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7237445_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:24254525(-)-22:24256334(-)__22_24230501_24255501D;SPAN=1809;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:59 GQ:30.2 PL:[30.2, 0.0, 112.7] SR:0 DR:14 LR:-30.23 LO:32.92);ALT=[chr22:24256334[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	24276436	+	chr22	24279226	+	.	102	97	7238239_1	99.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=CG;MAPQ=60;MATEID=7238239_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_24255001_24280001_53C;SPAN=2790;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:170 DP:40 GQ:46 PL:[505.0, 46.0, 0.0] SR:97 DR:102 LR:-505.0 LO:505.0);ALT=G[chr22:24279226[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24552045	+	chr22	24560367	+	.	9	5	7238623_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7238623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24549001_24574001_331C;SPAN=8322;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:79 GQ:18.2 PL:[18.2, 0.0, 173.3] SR:5 DR:9 LR:-18.21 LO:25.61);ALT=G[chr22:24560367[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24561595	+	chr22	24562605	+	.	3	3	7238647_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7238647_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24549001_24574001_126C;SPAN=1010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:102 GQ:10.8 PL:[0.0, 10.8, 267.3] SR:3 DR:3 LR:11.13 LO:8.092);ALT=G[chr22:24562605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24616558	+	chr22	24620963	+	.	8	0	7239064_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7239064_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:24616558(+)-22:24620963(-)__22_24598001_24623001D;SPAN=4405;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:109 GQ:3 PL:[0.0, 3.0, 270.6] SR:0 DR:8 LR:3.123 LO:14.39);ALT=A[chr22:24620963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24952039	+	chr22	24953624	+	.	97	14	7240580_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7240580_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24941001_24966001_110C;SPAN=1585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:112 GQ:30 PL:[330.0, 30.0, 0.0] SR:14 DR:97 LR:-330.1 LO:330.1);ALT=G[chr22:24953624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24952066	+	chr22	24963945	+	.	54	0	7240581_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7240581_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:24952066(+)-22:24963945(-)__22_24941001_24966001D;SPAN=11879;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:54 DP:116 GQ:99 PL:[146.9, 0.0, 133.7] SR:0 DR:54 LR:-146.9 LO:146.9);ALT=G[chr22:24963945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24953768	+	chr22	24963948	+	.	0	96	7240589_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CCAG;MAPQ=60;MATEID=7240589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_24941001_24966001_184C;SPAN=10180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:96 DP:158 GQ:99 PL:[274.1, 0.0, 109.1] SR:96 DR:0 LR:-278.0 LO:278.0);ALT=G[chr22:24963948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	24964144	+	chr22	24967882	+	.	6	16	7240629_1	60.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7240629_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_24941001_24966001_307C;SPAN=3738;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:44 GQ:44.3 PL:[60.8, 0.0, 44.3] SR:16 DR:6 LR:-60.81 LO:60.81);ALT=G[chr22:24967882[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	25177789	-	chr22	25179545	+	.	8	0	7241768_1	1.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7241768_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:25177789(-)-22:25179545(-)__22_25161501_25186501D;SPAN=1756;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:93 GQ:1.4 PL:[1.4, 0.0, 222.5] SR:0 DR:8 LR:-1.212 LO:14.96);ALT=[chr22:25179545[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	25455261	+	chr22	25456439	-	.	8	0	7242825_1	8.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7242825_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:25455261(+)-22:25456439(+)__22_25455501_25480501D;SPAN=1178;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:67 GQ:8.3 PL:[8.3, 0.0, 153.5] SR:0 DR:8 LR:-8.256 LO:16.17);ALT=C]chr22:25456439];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr22	28293882	+	chr22	28306952	+	.	0	8	7253317_1	11.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7253317_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_28297501_28322501_8C;SPAN=13070;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:54 GQ:11.9 PL:[11.9, 0.0, 117.5] SR:8 DR:0 LR:-11.78 LO:16.98);ALT=T[chr22:28306952[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	28307099	+	chr22	28315160	+	CCTGAACAGAACATGGCAAAACCACACGG	16	4	7253349_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=CCTGAACAGAACATGGCAAAACCACACGG;MAPQ=60;MATEID=7253349_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_28297501_28322501_233C;SPAN=8061;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:147 GQ:16.4 PL:[16.4, 0.0, 339.8] SR:4 DR:16 LR:-16.29 LO:34.1);ALT=T[chr22:28315160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	28315575	+	chr22	28320333	+	.	16	0	7253368_1	23.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7253368_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:28315575(+)-22:28320333(-)__22_28297501_28322501D;SPAN=4758;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:110 GQ:23 PL:[23.0, 0.0, 244.1] SR:0 DR:16 LR:-23.01 LO:33.81);ALT=A[chr22:28320333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	28315575	+	chr22	28318004	+	.	22	0	7253367_1	47.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7253367_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:28315575(+)-22:28318004(-)__22_28297501_28322501D;SPAN=2429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:93 GQ:47.6 PL:[47.6, 0.0, 176.3] SR:0 DR:22 LR:-47.43 LO:51.69);ALT=A[chr22:28318004[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	28318166	+	chr22	28320334	+	.	4	13	7253374_1	24.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7253374_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_28297501_28322501_138C;SPAN=2168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:118 GQ:24.2 PL:[24.2, 0.0, 261.8] SR:13 DR:4 LR:-24.15 LO:35.85);ALT=G[chr22:28320334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	29193195	+	chr22	29195045	+	.	0	17	7256386_1	21.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7256386_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_29179501_29204501_415C;SPAN=1850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:128 GQ:21.5 PL:[21.5, 0.0, 288.8] SR:17 DR:0 LR:-21.44 LO:35.2);ALT=T[chr22:29195045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	29193240	+	chr22	29196304	+	.	10	0	7256387_1	0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7256387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:29193240(+)-22:29196304(-)__22_29179501_29204501D;SPAN=3064;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:151 GQ:7.6 PL:[0.0, 7.6, 379.5] SR:0 DR:10 LR:7.9 LO:17.52);ALT=G[chr22:29196304[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	29195143	+	chr22	29196285	+	.	55	81	7256402_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7256402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_29179501_29204501_262C;SPAN=1142;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:100 DP:162 GQ:99 PL:[286.4, 0.0, 104.9] SR:81 DR:55 LR:-290.7 LO:290.7);ALT=T[chr22:29196285[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	29966522	+	chr22	29976974	+	.	24	4	7260068_1	53.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7260068_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_29963501_29988501_255C;SPAN=10452;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:122 GQ:53 PL:[53.0, 0.0, 241.1] SR:4 DR:24 LR:-52.77 LO:59.74);ALT=C[chr22:29976974[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30136722	+	chr22	30144407	+	TCAGTAGAAACTTCCTGCAGGGCCGCTTGTTCTGCTCATCCAGCAAGATGGCAGCTGCAT	0	21	7260465_1	36.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TCAGTAGAAACTTCCTGCAGGGCCGCTTGTTCTGCTCATCCAGCAAGATGGCAGCTGCAT;MAPQ=60;MATEID=7260465_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_30135001_30160001_183C;SPAN=7685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:120 GQ:36.8 PL:[36.8, 0.0, 254.6] SR:21 DR:0 LR:-36.81 LO:46.23);ALT=G[chr22:30144407[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30144593	+	chr22	30162808	+	.	14	0	7260676_1	31.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7260676_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:30144593(+)-22:30162808(-)__22_30159501_30184501D;SPAN=18215;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:54 GQ:31.7 PL:[31.7, 0.0, 97.7] SR:0 DR:14 LR:-31.58 LO:33.55);ALT=T[chr22:30162808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30163537	+	chr22	30165666	+	.	138	112	7260691_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7260691_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30159501_30184501_288C;SPAN=2129;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:208 DP:226 GQ:61 PL:[670.0, 61.0, 0.0] SR:112 DR:138 LR:-670.1 LO:670.1);ALT=G[chr22:30165666[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30230566	+	chr22	30234165	+	.	11	0	7261270_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7261270_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:30230566(+)-22:30234165(-)__22_30233001_30258001D;SPAN=3599;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:70 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:0 DR:11 LR:-17.35 LO:23.65);ALT=A[chr22:30234165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30279348	+	chr22	30353024	+	.	5	10	7261367_1	21.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7261367_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30331001_30356001_230C;SPAN=73676;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:55 GQ:21.5 PL:[21.5, 0.0, 110.6] SR:10 DR:5 LR:-21.41 LO:24.93);ALT=G[chr22:30353024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30742512	+	chr22	30748940	+	.	0	9	7262913_1	14.0	.	EVDNC=ASSMB;HOMSEQ=CTGG;MAPQ=60;MATEID=7262913_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30747501_30772501_45C;SPAN=6428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:57 GQ:14.3 PL:[14.3, 0.0, 123.2] SR:9 DR:0 LR:-14.27 LO:19.37);ALT=G[chr22:30748940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30749065	+	chr22	30752719	+	.	0	21	7262918_1	39.0	.	EVDNC=ASSMB;HOMSEQ=CTGT;MAPQ=60;MATEID=7262918_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30747501_30772501_451C;SPAN=3654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:111 GQ:39.5 PL:[39.5, 0.0, 227.6] SR:21 DR:0 LR:-39.25 LO:47.02);ALT=T[chr22:30752719[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30984163	+	chr22	30985177	+	.	0	5	7263905_1	0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7263905_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30968001_30993001_179C;SPAN=1014;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:102 GQ:10.8 PL:[0.0, 10.8, 267.3] SR:5 DR:0 LR:11.13 LO:8.092);ALT=T[chr22:30985177[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	30984195	+	chr22	30987796	+	.	8	0	7263906_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7263906_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:30984195(+)-22:30987796(-)__22_30968001_30993001D;SPAN=3601;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:0 DR:8 LR:1.497 LO:14.59);ALT=T[chr22:30987796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	31003382	+	chr22	31006857	+	.	7	9	7264545_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7264545_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_30992501_31017501_118C;SPAN=3475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:115 GQ:11.9 PL:[11.9, 0.0, 266.0] SR:9 DR:7 LR:-11.76 LO:25.94);ALT=G[chr22:31006857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	31796733	+	chr22	31799013	+	.	0	11	7267126_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AGGTTT;MAPQ=60;MATEID=7267126_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_31776501_31801501_163C;SPAN=2280;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:108 GQ:7.1 PL:[7.1, 0.0, 254.6] SR:11 DR:0 LR:-7.051 LO:21.42);ALT=T[chr22:31799013[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32340810	+	chr22	32352125	+	.	15	37	7269891_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTGA;MAPQ=60;MATEID=7269891_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_32340001_32365001_135C;SPAN=11315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:46 DP:103 GQ:99 PL:[124.1, 0.0, 124.1] SR:37 DR:15 LR:-123.9 LO:123.9);ALT=A[chr22:32352125[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32802748	+	chr22	32808049	+	ATGAACAATTCCAGGCAGGGCTGCCACATTGCCAATCTGTTTCATGGCTGGCAGGAAGCCACCAACACCACCACCTCGACAGGCATTCCTTAATTCCTCAAACATCAATTTCTCCAGAGCATCATTCACATAGAAAACACCTTCA	0	25	7271716_1	68.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=ATGAACAATTCCAGGCAGGGCTGCCACATTGCCAATCTGTTTCATGGCTGGCAGGAAGCCACCAACACCACCACCTCGACAGGCATTCCTTAATTCCTCAAACATCAATTTCTCCAGAGCATCATTCACATAGAAAACACCTTCA;MAPQ=60;MATEID=7271716_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_22_32781001_32806001_437C;SPAN=5301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:50 GQ:52.4 PL:[68.9, 0.0, 52.4] SR:25 DR:0 LR:-69.1 LO:69.1);ALT=G[chr22:32808049[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32804869	+	chr22	32808135	+	.	16	0	7271891_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7271891_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:32804869(+)-22:32808135(-)__22_32805501_32830501D;SPAN=3266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:72 GQ:33.5 PL:[33.5, 0.0, 139.1] SR:0 DR:16 LR:-33.31 LO:37.09);ALT=G[chr22:32808135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32871094	+	chr22	32874963	+	.	16	0	7272193_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7272193_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:32871094(+)-22:32874963(-)__22_32854501_32879501D;SPAN=3869;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:94 GQ:27.5 PL:[27.5, 0.0, 199.1] SR:0 DR:16 LR:-27.35 LO:35.01);ALT=G[chr22:32874963[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	32875262	+	chr22	32879883	+	.	4	6	7272227_1	13.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7272227_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_32879001_32904001_104C;SPAN=4621;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:59 GQ:13.7 PL:[13.7, 0.0, 129.2] SR:6 DR:4 LR:-13.72 LO:19.22);ALT=G[chr22:32879883[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	33759249	+	chr22	33838399	+	AACTACT	0	18	7276054_1	51.0	.	EVDNC=ASSMB;INSERTION=AACTACT;MAPQ=60;MATEID=7276054_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_33834501_33859501_242C;SPAN=79150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:29 GQ:18.5 PL:[51.5, 0.0, 18.5] SR:18 DR:0 LR:-52.4 LO:52.4);ALT=A[chr22:33838399[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	35653575	+	chr22	35659068	+	.	15	0	7282500_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7282500_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:35653575(+)-22:35659068(-)__22_35647501_35672501D;SPAN=5493;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:89 GQ:25.4 PL:[25.4, 0.0, 190.4] SR:0 DR:15 LR:-25.4 LO:32.75);ALT=A[chr22:35659068[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	35796599	+	chr22	35799197	+	.	0	11	7283058_1	8.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=7283058_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_35794501_35819501_121C;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:102 GQ:8.9 PL:[8.9, 0.0, 236.6] SR:11 DR:0 LR:-8.677 LO:21.71);ALT=G[chr22:35799197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36613001	+	chr22	36614319	+	.	0	47	7286330_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TT;MAPQ=60;MATEID=7286330_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_36603001_36628001_365C;SPAN=1318;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:47 DP:72 GQ:36.8 PL:[135.8, 0.0, 36.8] SR:47 DR:0 LR:-138.6 LO:138.6);ALT=T[chr22:36614319[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36685347	+	chr22	36688032	+	.	6	5	7286927_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTGG;MAPQ=60;MATEID=7286927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36676501_36701501_20C;SPAN=2685;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:103 GQ:1.2 PL:[0.0, 1.2, 250.8] SR:5 DR:6 LR:1.497 LO:14.59);ALT=G[chr22:36688032[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36690345	+	chr22	36691549	+	CGCTTCGTCTGCTCCAGCTGCTCCGCCAGCTCCTCCACGGCCTGTGAGTGCTTCTGCCTCATCTCCTGGATCTGGGCCTCGTGGGTCTTGGCCTCCTCCTCCAGGGTCTTCTTCAGGATGTTCACCTCCTGCTCACGTTTTG	6	15	7286950_1	30.0	.	DISC_MAPQ=52;EVDNC=TSI_G;HOMSEQ=ACCTG;INSERTION=CGCTTCGTCTGCTCCAGCTGCTCCGCCAGCTCCTCCACGGCCTGTGAGTGCTTCTGCCTCATCTCCTGGATCTGGGCCTCGTGGGTCTTGGCCTCCTCCTCCAGGGTCTTCTTCAGGATGTTCACCTCCTGCTCACGTTTTG;MAPQ=60;MATEID=7286950_2;MATENM=1;NM=0;NUMPARTS=3;SCTG=c_22_36676501_36701501_236C;SPAN=1204;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:94 GQ:30.8 PL:[30.8, 0.0, 195.8] SR:15 DR:6 LR:-30.65 LO:37.69);ALT=C[chr22:36691549[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36695090	+	chr22	36696172	+	.	4	11	7286977_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7286977_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36676501_36701501_463C;SPAN=1082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:115 GQ:15.2 PL:[15.2, 0.0, 262.7] SR:11 DR:4 LR:-15.06 LO:28.42);ALT=T[chr22:36696172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36702654	+	chr22	36705327	+	.	5	5	7286601_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7286601_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36701001_36726001_131C;SPAN=2673;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:128 GQ:4.8 PL:[0.0, 4.8, 320.1] SR:5 DR:5 LR:4.969 LO:16.01);ALT=C[chr22:36705327[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36705443	+	chr22	36708091	+	.	2	7	7286615_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CACCT;MAPQ=60;MATEID=7286615_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36701001_36726001_115C;SPAN=2648;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:115 GQ:4.5 PL:[0.0, 4.5, 287.1] SR:7 DR:2 LR:4.748 LO:14.2);ALT=T[chr22:36708091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36737571	+	chr22	36744949	+	.	8	6	7286832_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=7286832_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36725501_36750501_161C;SPAN=7378;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:109 GQ:6.8 PL:[6.8, 0.0, 257.6] SR:6 DR:8 LR:-6.78 LO:21.38);ALT=T[chr22:36744949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36745302	+	chr22	36783850	+	.	51	38	7287002_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=7287002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36774501_36799501_117C;SPAN=38548;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:70 DP:38 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:38 DR:51 LR:-208.0 LO:208.0);ALT=T[chr22:36783850[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36872903	+	chr22	36876619	+	.	0	20	7287479_1	35.0	.	EVDNC=ASSMB;HOMSEQ=CAC;MAPQ=60;MATEID=7287479_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36872501_36897501_173C;SPAN=3716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:114 GQ:35.3 PL:[35.3, 0.0, 239.9] SR:20 DR:0 LR:-35.13 LO:44.05);ALT=C[chr22:36876619[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36920779	+	chr22	36922044	+	TTGTGTACCTCTTATCTTGGTATGTGGCTCCTGTCCAGTCTGCA	5	108	7287918_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=ACCT;INSERTION=TTGTGTACCTCTTATCTTGGTATGTGGCTCCTGTCCAGTCTGCA;MAPQ=60;MATEID=7287918_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_36897001_36922001_121C;SPAN=1265;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:111 DP:91 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:108 DR:5 LR:-326.8 LO:326.8);ALT=T[chr22:36922044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36920837	+	chr22	36925120	+	.	38	0	7287919_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7287919_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36920837(+)-22:36925120(-)__22_36897001_36922001D;SPAN=4283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:38 DP:39 GQ:10.5 PL:[115.5, 10.5, 0.0] SR:0 DR:38 LR:-115.5 LO:115.5);ALT=A[chr22:36925120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36921808	+	chr22	36925122	+	.	51	0	7287926_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7287926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:36921808(+)-22:36925122(-)__22_36897001_36922001D;SPAN=3314;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:51 DP:54 GQ:14.4 PL:[158.4, 14.4, 0.0] SR:0 DR:51 LR:-158.4 LO:158.4);ALT=C[chr22:36925122[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	36922181	+	chr22	36925123	+	.	97	17	7287927_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7287927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_36897001_36922001_308C;SPAN=2942;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:103 DP:0 GQ:27.6 PL:[303.6, 27.6, 0.0] SR:17 DR:97 LR:-303.7 LO:303.7);ALT=G[chr22:36925123[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37143176	+	chr22	37147896	+	.	83	49	7288674_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AGTAGCT;MAPQ=60;MATEID=7288674_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37117501_37142501_166C;SPAN=4720;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:115 DP:0 GQ:30.9 PL:[339.9, 30.9, 0.0] SR:49 DR:83 LR:-340.0 LO:340.0);ALT=T[chr22:37147896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37154454	+	chr22	37158948	+	.	0	12	7288442_1	16.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7288442_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37142001_37167001_206C;SPAN=4494;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:87 GQ:16.1 PL:[16.1, 0.0, 194.3] SR:12 DR:0 LR:-16.04 LO:25.06);ALT=C[chr22:37158948[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37257225	+	chr22	37260960	+	.	9	0	7288941_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7288941_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37257225(+)-22:37260960(-)__22_37240001_37265001D;SPAN=3735;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:161 GQ:13.6 PL:[0.0, 13.6, 415.9] SR:0 DR:9 LR:13.91 LO:15.09);ALT=C[chr22:37260960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37257245	+	chr22	37260085	+	.	23	30	7288942_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7288942_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37240001_37265001_394C;SPAN=2840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:138 GQ:98 PL:[98.0, 0.0, 236.6] SR:30 DR:23 LR:-97.95 LO:101.1);ALT=G[chr22:37260085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37272137	+	chr22	37273668	+	.	3	5	7289085_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7289085_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37264501_37289501_304C;SPAN=1531;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:103 GQ:7.8 PL:[0.0, 7.8, 264.0] SR:5 DR:3 LR:8.099 LO:10.17);ALT=G[chr22:37273668[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37415952	+	chr22	37420230	+	.	31	0	7289659_1	77.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7289659_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37415952(+)-22:37420230(-)__22_37411501_37436501D;SPAN=4278;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:93 GQ:77.3 PL:[77.3, 0.0, 146.6] SR:0 DR:31 LR:-77.14 LO:78.38);ALT=G[chr22:37420230[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37622119	+	chr22	37627270	+	.	8	0	7290591_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7290591_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37622119(+)-22:37627270(-)__22_37607501_37632501D;SPAN=5151;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:110 GQ:3.3 PL:[0.0, 3.3, 273.9] SR:0 DR:8 LR:3.394 LO:14.36);ALT=T[chr22:37627270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37622844	+	chr22	37627271	+	.	13	12	7290595_1	41.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7290595_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37607501_37632501_280C;SPAN=4427;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:141 GQ:41.3 PL:[41.3, 0.0, 298.7] SR:12 DR:13 LR:-41.02 LO:52.52);ALT=C[chr22:37627271[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37627432	+	chr22	37628840	+	TGGCGCGGACGTTCTCATAAGAGGCTGGGCTGACGAGGGAGAAGCAGATGAGGAAGACGT	8	99	7290625_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=TGGCGCGGACGTTCTCATAAGAGGCTGGGCTGACGAGGGAGAAGCAGATGAGGAAGACGT;MAPQ=60;MATEID=7290625_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_37607501_37632501_97C;SPAN=1408;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:106 DP:176 GQ:99 PL:[302.3, 0.0, 124.1] SR:99 DR:8 LR:-306.2 LO:306.2);ALT=T[chr22:37628840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37627490	+	chr22	37640184	+	.	15	0	7290443_1	9.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7290443_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37627490(+)-22:37640184(-)__22_37632001_37657001D;SPAN=12694;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:148 GQ:9.5 PL:[9.5, 0.0, 349.4] SR:0 DR:15 LR:-9.418 LO:29.18);ALT=G[chr22:37640184[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37628082	+	chr22	37640178	+	.	53	0	7290446_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7290446_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37628082(+)-22:37640178(-)__22_37632001_37657001D;SPAN=12096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:53 DP:112 GQ:99 PL:[144.8, 0.0, 125.0] SR:0 DR:53 LR:-144.7 LO:144.7);ALT=T[chr22:37640178[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37637699	+	chr22	37640153	+	.	81	58	7290464_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=CC;MAPQ=60;MATEID=7290464_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CCC;SCTG=c_22_37632001_37657001_39C;SPAN=2454;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:157 GQ:99 PL:[277.7, 0.0, 102.8] SR:58 DR:81 LR:-282.0 LO:282.0);ALT=C[chr22:37640153[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37966743	+	chr22	37967856	+	.	0	72	7291698_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7291698_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_37950501_37975501_24C;SPAN=1113;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:72 DP:162 GQ:99 PL:[194.0, 0.0, 197.3] SR:72 DR:0 LR:-193.8 LO:193.8);ALT=C[chr22:37967856[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	37967989	+	chr22	37975965	+	.	73	0	7292182_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7292182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:37967989(+)-22:37975965(-)__22_37975001_38000001D;SPAN=7976;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:73 DP:98 GQ:23 PL:[214.4, 0.0, 23.0] SR:0 DR:73 LR:-223.4 LO:223.4);ALT=C[chr22:37975965[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38005133	+	chr22	38012927	+	.	13	0	7291972_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7291972_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:38005133(+)-22:38012927(-)__22_37999501_38024501D;SPAN=7794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:107 GQ:14 PL:[14.0, 0.0, 245.0] SR:0 DR:13 LR:-13.92 LO:26.38);ALT=T[chr22:38012927[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38035785	+	chr22	38037131	+	.	10	0	7291783_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7291783_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:38035785(+)-22:38037131(-)__22_38024001_38049001D;SPAN=1346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:70 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-14.05 LO:21.05);ALT=C[chr22:38037131[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38035853	+	chr22	38037378	+	CACCCCGGAGACCGCTGAGTTCCTGGGTGAGGACCTGCTG	13	26	7291785_1	79.0	.	DISC_MAPQ=58;EVDNC=TSI_G;HOMSEQ=CAGGTA;INSERTION=CACCCCGGAGACCGCTGAGTTCCTGGGTGAGGACCTGCTG;MAPQ=60;MATEID=7291785_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_38024001_38049001_207C;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:97 GQ:79.4 PL:[79.4, 0.0, 155.3] SR:26 DR:13 LR:-79.35 LO:80.72);ALT=G[chr22:38037378[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38046733	+	chr22	38049784	+	.	2	2	7291817_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGG;MAPQ=60;MATEID=7291817_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38024001_38049001_107C;SPAN=3051;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:2 DR:2 LR:4.677 LO:6.851);ALT=G[chr22:38049784[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38071719	+	chr22	38072993	+	.	30	59	7292138_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7292138_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38048501_38073501_271C;SPAN=1274;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:79 DP:264 GQ:99 PL:[189.4, 0.0, 450.2] SR:59 DR:30 LR:-189.3 LO:195.2);ALT=G[chr22:38072993[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38073072	+	chr22	38074488	+	.	17	127	7292462_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7292462_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38073001_38098001_250C;SPAN=1416;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:144 DP:826 GQ:99 PL:[251.8, 0.0, 1754.0] SR:127 DR:17 LR:-251.6 LO:316.7);ALT=G[chr22:38074488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38082483	+	chr22	38083916	+	.	21	7	7292504_1	45.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7292504_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38073001_38098001_90C;SPAN=1433;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:113 GQ:45.5 PL:[45.5, 0.0, 227.0] SR:7 DR:21 LR:-45.31 LO:52.32);ALT=G[chr22:38083916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38082503	+	chr22	38084855	+	.	8	0	7292506_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7292506_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:38082503(+)-22:38084855(-)__22_38073001_38098001D;SPAN=2352;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:125 GQ:7.2 PL:[0.0, 7.2, 316.8] SR:0 DR:8 LR:7.458 LO:13.9);ALT=G[chr22:38084855[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38087433	+	chr22	38089337	+	.	0	8	7292540_1	0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=7292540_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38073001_38098001_76C;SPAN=1904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:112 GQ:3.6 PL:[0.0, 3.6, 277.2] SR:8 DR:0 LR:3.936 LO:14.29);ALT=T[chr22:38089337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38245490	+	chr22	38247284	+	CGGCTTATGACCCCTACGCTTATCCCAGCGACTATGATATGCACA	126	42	7293202_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CAGG;INSERTION=CGGCTTATGACCCCTACGCTTATCCCAGCGACTATGATATGCACA;MAPQ=60;MATEID=7293202_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_38244501_38269501_180C;SPAN=1794;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:196 DP:191 GQ:52.9 PL:[580.9, 52.9, 0.0] SR:42 DR:126 LR:-580.9 LO:580.9);ALT=G[chr22:38247284[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38247497	+	chr22	38251570	+	.	0	59	7293211_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7293211_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38244501_38269501_46C;SPAN=4073;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:59 DP:121 GQ:99 PL:[162.2, 0.0, 129.2] SR:59 DR:0 LR:-162.1 LO:162.1);ALT=G[chr22:38251570[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38259352	+	chr22	38266180	+	.	5	4	7293261_1	0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7293261_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38244501_38269501_118C;SPAN=6828;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:118 GQ:5.4 PL:[0.0, 5.4, 297.0] SR:4 DR:5 LR:5.561 LO:14.1);ALT=G[chr22:38266180[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38282852	+	chr22	38284431	+	.	3	124	7293806_1	99.0	.	DISC_MAPQ=38;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=47;MATEID=7293806_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_22_38269001_38294001_379C;SPAN=1579;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:127 DP:170 GQ:39.7 PL:[373.1, 0.0, 39.7] SR:124 DR:3 LR:-388.9 LO:388.9);ALT=G[chr22:38284431[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38349814	+	chr22	38355351	+	TTTTGATGGCGACGACTTTGATGATGTGGAGGAGGATGAAGGGCTAGATGACTTGGAGAATGCCGAAG	41	42	7293627_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AGG;INSERTION=TTTTGATGGCGACGACTTTGATGATGTGGAGGAGGATGAAGGGCTAGATGACTTGGAGAATGCCGAAG;MAPQ=60;MATEID=7293627_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_38342501_38367501_184C;SPAN=5537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:63 DP:122 GQ:99 PL:[175.1, 0.0, 119.0] SR:42 DR:41 LR:-175.4 LO:175.4);ALT=A[chr22:38355351[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38349814	+	chr22	38352780	+	.	18	11	7293626_1	40.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=7293626_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=TTT;SCTG=c_22_38342501_38367501_184C;SPAN=2966;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:121 GQ:40.1 PL:[40.1, 0.0, 251.3] SR:11 DR:18 LR:-39.84 LO:48.84);ALT=A[chr22:38352780[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38355484	+	chr22	38363106	+	.	0	41	7293664_1	98.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7293664_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38342501_38367501_61C;SPAN=7622;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:136 GQ:98.6 PL:[98.6, 0.0, 230.6] SR:41 DR:0 LR:-98.5 LO:101.5);ALT=G[chr22:38363106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38598221	+	chr22	38609829	+	.	0	9	7294753_1	1.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=7294753_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38587501_38612501_93C;SPAN=11608;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:105 GQ:1.4 PL:[1.4, 0.0, 252.2] SR:9 DR:0 LR:-1.262 LO:16.82);ALT=T[chr22:38609829[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38888121	+	chr22	38889715	+	.	0	25	7296071_1	51.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7296071_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38881501_38906501_38C;SPAN=1594;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:116 GQ:51.2 PL:[51.2, 0.0, 229.4] SR:25 DR:0 LR:-51.1 LO:57.58);ALT=C[chr22:38889715[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38895504	+	chr22	38897135	+	.	0	8	7296099_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7296099_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38881501_38906501_328C;SPAN=1631;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:107 GQ:2.4 PL:[0.0, 2.4, 264.0] SR:8 DR:0 LR:2.581 LO:14.46);ALT=A[chr22:38897135[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	38897286	+	chr22	38901956	+	.	4	8	7296117_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7296117_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_38881501_38906501_443C;SPAN=4670;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:92 GQ:11.6 PL:[11.6, 0.0, 209.6] SR:8 DR:4 LR:-11.39 LO:22.24);ALT=C[chr22:38901956[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39178892	+	chr22	39190072	+	.	9	0	7297357_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7297357_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39178892(+)-22:39190072(-)__22_39175501_39200501D;SPAN=11180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:9 DP:125 GQ:3.9 PL:[0.0, 3.9, 310.2] SR:0 DR:9 LR:4.157 LO:16.11);ALT=A[chr22:39190072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39234361	-	chr22	39235548	+	.	9	0	7297451_1	0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=7297451_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39234361(-)-22:39235548(-)__22_39224501_39249501D;SPAN=1187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:107 GQ:0.8 PL:[0.8, 0.0, 258.2] SR:0 DR:9 LR:-0.7201 LO:16.74);ALT=[chr22:39235548[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	39294108	+	chr22	39298685	+	.	90	81	7297678_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TAAA;MAPQ=60;MATEID=7297678_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39298001_39323001_190C;SPAN=4577;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:135 DP:20 GQ:36.3 PL:[399.3, 36.3, 0.0] SR:81 DR:90 LR:-399.4 LO:399.4);ALT=A[chr22:39298685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39410384	+	chr22	39411596	+	.	18	6	7298476_1	36.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=TCAG;MAPQ=19;MATEID=7298476_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39396001_39421001_3C;SPAN=1212;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:108 GQ:36.8 PL:[36.8, 0.0, 224.9] SR:6 DR:18 LR:-36.76 LO:44.58);ALT=G[chr22:39411596[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39410386	+	chr22	39413766	+	.	9	0	7298477_1	3.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7298477_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39410386(+)-22:39413766(-)__22_39396001_39421001D;SPAN=3380;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:96 GQ:3.8 PL:[3.8, 0.0, 228.2] SR:0 DR:9 LR:-3.7 LO:17.19);ALT=T[chr22:39413766[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39411758	+	chr22	39413767	+	.	2	11	7298481_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCAGGT;MAPQ=60;MATEID=7298481_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39396001_39421001_101C;SPAN=2009;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:90 GQ:15.2 PL:[15.2, 0.0, 203.3] SR:11 DR:2 LR:-15.23 LO:24.87);ALT=T[chr22:39413767[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39540875	+	chr22	39568639	+	.	0	8	7299122_1	15.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7299122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39567501_39592501_144C;SPAN=27764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:41 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:8 DR:0 LR:-15.3 LO:18.03);ALT=G[chr22:39568639[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39711568	+	chr22	39713500	+	.	10	0	7299417_1	0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=7299417_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39711568(+)-22:39713500(-)__22_39690001_39715001D;SPAN=1932;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:10 DP:189 GQ:18.1 PL:[0.0, 18.1, 495.1] SR:0 DR:10 LR:18.19 LO:16.52);ALT=A[chr22:39713500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39746114	+	chr22	39770320	+	.	41	12	7299716_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7299716_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39763501_39788501_68C;SPAN=24206;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:65 GQ:25.4 PL:[131.0, 0.0, 25.4] SR:12 DR:41 LR:-134.8 LO:134.8);ALT=G[chr22:39770320[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39772202	+	chr22	39773602	+	.	0	7	7299740_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7299740_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39763501_39788501_225C;SPAN=1400;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:108 GQ:6 PL:[0.0, 6.0, 273.9] SR:7 DR:0 LR:6.153 LO:12.2);ALT=G[chr22:39773602[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39925682	+	chr22	39928690	+	.	14	0	7300475_1	14.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7300475_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39925682(+)-22:39928690(-)__22_39910501_39935501D;SPAN=3008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:116 GQ:14.9 PL:[14.9, 0.0, 265.7] SR:0 DR:14 LR:-14.79 LO:28.36);ALT=C[chr22:39928690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39925923	+	chr22	39928400	+	.	0	62	7300477_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7300477_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_39910501_39935501_275C;SPAN=2477;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:131 GQ:99 PL:[169.4, 0.0, 146.3] SR:62 DR:0 LR:-169.2 LO:169.2);ALT=C[chr22:39928400[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	39925974	+	chr22	39928691	+	.	62	0	7300478_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7300478_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:39925974(+)-22:39928691(-)__22_39910501_39935501D;SPAN=2717;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:62 DP:108 GQ:86.3 PL:[175.4, 0.0, 86.3] SR:0 DR:62 LR:-177.0 LO:177.0);ALT=A[chr22:39928691[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40742715	+	chr22	40745832	+	.	30	29	7303512_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GCAG;MAPQ=60;MATEID=7303512_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_40743501_40768501_15C;SPAN=3117;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:59 GQ:6 PL:[155.1, 6.0, 0.0] SR:29 DR:30 LR:-159.9 LO:159.9);ALT=G[chr22:40745832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40760371	+	chr22	40762437	+	.	2	6	7303583_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAGGT;MAPQ=60;MATEID=7303583_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_40743501_40768501_36C;SPAN=2066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:127 GQ:7.8 PL:[0.0, 7.8, 323.4] SR:6 DR:2 LR:7.999 LO:13.84);ALT=T[chr22:40762437[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40761062	+	chr22	40762436	+	.	0	24	7303586_1	45.0	.	EVDNC=ASSMB;HOMSEQ=GCAGGT;MAPQ=60;MATEID=7303586_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_40743501_40768501_171C;SPAN=1374;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:126 GQ:45.2 PL:[45.2, 0.0, 259.7] SR:24 DR:0 LR:-45.09 LO:53.82);ALT=T[chr22:40762436[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40798209	+	chr22	40800249	+	.	0	7	7303771_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7303771_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_40792501_40817501_447C;SPAN=2040;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:87 GQ:0.3 PL:[0.0, 0.3, 211.2] SR:7 DR:0 LR:0.4634 LO:12.88);ALT=G[chr22:40800249[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40831558	+	chr22	40859225	+	.	5	7	7303929_1	16.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7303929_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_40841501_40866501_37C;SPAN=27667;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:50 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:7 DR:5 LR:-16.16 LO:19.94);ALT=G[chr22:40859225[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	40948372	+	chr22	41032482	+	.	6	3	7304703_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7304703_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41013001_41038001_321C;SPAN=84110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:39 GQ:9.2 PL:[9.2, 0.0, 85.1] SR:3 DR:6 LR:-9.24 LO:12.84);ALT=C[chr22:41032482[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41253250	+	chr22	41264999	+	.	7	3	7305941_1	12.0	.	DISC_MAPQ=51;EVDNC=ASDIS;HOMSEQ=TCAGG;MAPQ=60;MATEID=7305941_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41233501_41258501_395C;SPAN=11749;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:3 DR:7 LR:-12.59 LO:17.19);ALT=G[chr22:41264999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347473	+	chr22	41351290	+	.	8	0	7306460_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7306460_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347473(+)-22:41351290(-)__22_41331501_41356501D;SPAN=3817;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:106 GQ:2.1 PL:[0.0, 2.1, 260.7] SR:0 DR:8 LR:2.31 LO:14.49);ALT=T[chr22:41351290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347480	+	chr22	41349557	+	.	0	33	7306461_1	76.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7306461_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41331501_41356501_256C;SPAN=2077;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:33 DP:121 GQ:76.4 PL:[76.4, 0.0, 215.0] SR:33 DR:0 LR:-76.15 LO:79.93);ALT=G[chr22:41349557[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347483	+	chr22	41363802	+	.	34	0	7306462_1	98.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7306462_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347483(+)-22:41363802(-)__22_41331501_41356501D;SPAN=16319;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:50 GQ:22.7 PL:[98.6, 0.0, 22.7] SR:0 DR:34 LR:-101.4 LO:101.4);ALT=T[chr22:41363802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347803	+	chr22	41349555	+	.	44	0	7306464_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7306464_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347803(+)-22:41349555(-)__22_41331501_41356501D;SPAN=1752;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:127 GQ:99 PL:[110.9, 0.0, 196.7] SR:0 DR:44 LR:-110.8 LO:112.2);ALT=G[chr22:41349555[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41347899	+	chr22	41360048	+	.	59	0	7306466_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7306466_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41347899(+)-22:41360048(-)__22_41331501_41356501D;SPAN=12149;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:69 GQ:8.7 PL:[184.8, 8.7, 0.0] SR:0 DR:59 LR:-189.4 LO:189.4);ALT=C[chr22:41360048[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41349637	+	chr22	41351291	+	.	0	8	7306474_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7306474_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41331501_41356501_179C;SPAN=1654;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:129 GQ:8.4 PL:[0.0, 8.4, 330.0] SR:8 DR:0 LR:8.541 LO:13.78);ALT=T[chr22:41351291[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41349638	+	chr22	41360051	+	.	0	116	7306475_1	99.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7306475_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41331501_41356501_335C;SPAN=10413;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:116 DP:73 GQ:31.2 PL:[343.2, 31.2, 0.0] SR:116 DR:0 LR:-343.3 LO:343.3);ALT=G[chr22:41360051[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41360121	+	chr22	41363803	+	.	0	128	7306116_1	99.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7306116_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41356001_41381001_341C;SPAN=3682;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:128 DP:173 GQ:42.4 PL:[375.8, 0.0, 42.4] SR:128 DR:0 LR:-390.9 LO:390.9);ALT=C[chr22:41363803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41363891	+	chr22	41368480	+	.	0	97	7306136_1	99.0	.	EVDNC=ASSMB;HOMSEQ=GTA;MAPQ=60;MATEID=7306136_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41356001_41381001_155C;SPAN=4589;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:97 DP:170 GQ:99 PL:[274.1, 0.0, 138.8] SR:97 DR:0 LR:-276.5 LO:276.5);ALT=A[chr22:41368480[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41601404	+	chr22	41605730	+	.	9	0	7307774_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7307774_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41601404(+)-22:41605730(-)__22_41576501_41601501D;SPAN=4326;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:69 GQ:11 PL:[11.0, 0.0, 156.2] SR:0 DR:9 LR:-11.02 LO:18.56);ALT=G[chr22:41605730[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41677087	+	chr22	41681990	+	.	0	7	7307935_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7307935_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41674501_41699501_370C;SPAN=4903;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:103 GQ:4.5 PL:[0.0, 4.5, 257.4] SR:7 DR:0 LR:4.798 LO:12.35);ALT=C[chr22:41681990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41856491	+	chr22	41863452	+	.	0	29	7309048_1	61.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7309048_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_41846001_41871001_331C;SPAN=6961;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:126 GQ:61.7 PL:[61.7, 0.0, 243.2] SR:29 DR:0 LR:-61.59 LO:67.74);ALT=T[chr22:41863452[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	41865224	+	chr22	41903793	+	.	10	0	7309093_1	20.0	.	DISC_MAPQ=51;EVDNC=DSCRD;IMPRECISE;MAPQ=51;MATEID=7309093_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:41865224(+)-22:41903793(-)__22_41846001_41871001D;SPAN=38569;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:48 GQ:20 PL:[20.0, 0.0, 95.9] SR:0 DR:10 LR:-20.01 LO:22.86);ALT=G[chr22:41903793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42022323	-	chr22	42023698	+	.	8	0	7309608_1	0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=7309608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42022323(-)-22:42023698(-)__22_42017501_42042501D;SPAN=1375;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:119 GQ:5.7 PL:[0.0, 5.7, 300.3] SR:0 DR:8 LR:5.832 LO:14.07);ALT=[chr22:42023698[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	42071200	+	chr22	42076248	+	.	0	91	7310092_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7310092_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42066501_42091501_161C;SPAN=5048;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:91 DP:148 GQ:98.6 PL:[260.3, 0.0, 98.6] SR:91 DR:0 LR:-264.3 LO:264.3);ALT=C[chr22:42076248[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42071233	+	chr22	42084796	+	.	61	0	7310094_1	99.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7310094_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42071233(+)-22:42084796(-)__22_42066501_42091501D;SPAN=13563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:61 DP:152 GQ:99 PL:[160.4, 0.0, 206.6] SR:0 DR:61 LR:-160.2 LO:160.5);ALT=T[chr22:42084796[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42071244	+	chr22	42078359	+	.	14	0	7310095_1	11.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7310095_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42071244(+)-22:42078359(-)__22_42066501_42091501D;SPAN=7115;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:131 GQ:11 PL:[11.0, 0.0, 304.7] SR:0 DR:14 LR:-10.72 LO:27.57);ALT=G[chr22:42078359[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42076369	+	chr22	42078360	+	.	20	5	7310126_1	34.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7310126_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42066501_42091501_52C;SPAN=1991;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:140 GQ:34.7 PL:[34.7, 0.0, 305.3] SR:5 DR:20 LR:-34.69 LO:47.3);ALT=C[chr22:42078360[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42076369	+	chr22	42084798	+	.	36	8	7310127_1	72.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7310127_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42066501_42091501_397C;SPAN=8429;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:170 GQ:72.8 PL:[72.8, 0.0, 340.1] SR:8 DR:36 LR:-72.78 LO:82.6);ALT=C[chr22:42084798[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42129934	+	chr22	42131118	-	.	10	0	7309892_1	5.0	.	DISC_MAPQ=47;EVDNC=DSCRD;IMPRECISE;MAPQ=47;MATEID=7309892_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42129934(+)-22:42131118(+)__22_42115501_42140501D;SPAN=1184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:103 GQ:5.3 PL:[5.3, 0.0, 242.9] SR:0 DR:10 LR:-5.105 LO:19.26);ALT=C]chr22:42131118];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr22	42229362	+	chr22	42262834	+	.	4	2	7310547_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7310547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42262501_42287501_290C;SPAN=33472;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:57 GQ:2.1 PL:[0.0, 2.1, 141.9] SR:2 DR:4 LR:2.239 LO:7.114);ALT=G[chr22:42262834[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42341311	+	chr22	42342421	+	TATTTGCTGTGAAGATTAACCACAAACACGATCAGGTCAATTCGGGGCCGATTCACACTGGAGGGCAAAGGGAGGGACTTTGCCAAGTGG	0	20	7310900_1	36.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=TATTTGCTGTGAAGATTAACCACAAACACGATCAGGTCAATTCGGGGCCGATTCACACTGGAGGGCAAAGGGAGGGACTTTGCCAAGTGG;MAPQ=60;MATEID=7310900_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_22_42336001_42361001_402C;SPAN=1110;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:111 GQ:36.2 PL:[36.2, 0.0, 230.9] SR:20 DR:0 LR:-35.95 LO:44.31);ALT=G[chr22:42342421[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42475958	+	chr22	42477929	+	.	40	84	7311743_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;MAPQ=60;MATEID=7311743_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42458501_42483501_304C;SPAN=1971;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:104 DP:159 GQ:85.7 PL:[300.2, 0.0, 85.7] SR:84 DR:40 LR:-306.8 LO:306.8);ALT=A[chr22:42477929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42478070	+	chr22	42479119	+	.	0	57	7311752_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACAGG;MAPQ=60;MATEID=7311752_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42458501_42483501_269C;SPAN=1049;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:57 DP:144 GQ:99 PL:[149.3, 0.0, 198.8] SR:57 DR:0 LR:-149.1 LO:149.6);ALT=G[chr22:42479119[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42483180	+	chr22	42486610	+	.	0	66	7311607_1	99.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7311607_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42483001_42508001_195C;SPAN=3430;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:66 DP:134 GQ:99 PL:[181.7, 0.0, 142.1] SR:66 DR:0 LR:-181.8 LO:181.8);ALT=C[chr22:42486610[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42912144	+	chr22	42914010	+	.	0	30	7313289_1	72.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7313289_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42899501_42924501_265C;SPAN=1866;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:98 GQ:72.5 PL:[72.5, 0.0, 164.9] SR:30 DR:0 LR:-72.48 LO:74.48);ALT=T[chr22:42914010[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42912195	+	chr22	42915739	+	.	21	0	7313290_1	43.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7313290_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42912195(+)-22:42915739(-)__22_42899501_42924501D;SPAN=3544;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:96 GQ:43.4 PL:[43.4, 0.0, 188.6] SR:0 DR:21 LR:-43.31 LO:48.52);ALT=G[chr22:42915739[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42914178	+	chr22	42915737	+	.	27	0	7313302_1	56.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7313302_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42914178(+)-22:42915737(-)__22_42899501_42924501D;SPAN=1559;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:122 GQ:56.3 PL:[56.3, 0.0, 237.8] SR:0 DR:27 LR:-56.07 LO:62.54);ALT=G[chr22:42915737[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42976379	+	chr22	42977949	+	.	8	0	7313387_1	0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=7313387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:42976379(+)-22:42977949(-)__22_42973001_42998001D;SPAN=1570;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:124 GQ:6.9 PL:[0.0, 6.9, 313.5] SR:0 DR:8 LR:7.187 LO:13.93);ALT=G[chr22:42977949[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	42999167	+	chr22	43010804	+	.	13	2	7313760_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=7313760_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_42997501_43022501_257C;SPAN=11637;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:94 GQ:17.6 PL:[17.6, 0.0, 209.0] SR:2 DR:13 LR:-17.45 LO:27.16);ALT=C[chr22:43010804[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43027042	+	chr22	43045298	+	.	17	0	7313856_1	38.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7313856_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43027042(+)-22:43045298(-)__22_43022001_43047001D;SPAN=18256;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:66 GQ:38.3 PL:[38.3, 0.0, 120.8] SR:0 DR:17 LR:-38.24 LO:40.68);ALT=T[chr22:43045298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43027458	+	chr22	43032721	+	.	0	65	7313858_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7313858_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43022001_43047001_81C;SPAN=5263;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:65 DP:137 GQ:99 PL:[177.5, 0.0, 154.4] SR:65 DR:0 LR:-177.5 LO:177.5);ALT=T[chr22:43032721[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43027507	+	chr22	43045300	+	.	41	0	7313859_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7313859_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43027507(+)-22:43045300(-)__22_43022001_43047001D;SPAN=17793;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:41 DP:54 GQ:8.6 PL:[120.8, 0.0, 8.6] SR:0 DR:41 LR:-126.2 LO:126.2);ALT=A[chr22:43045300[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43032853	+	chr22	43045301	+	.	50	7	7313877_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7313877_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43022001_43047001_196C;SPAN=12448;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:52 DP:85 GQ:56.3 PL:[148.7, 0.0, 56.3] SR:7 DR:50 LR:-150.8 LO:150.8);ALT=C[chr22:43045301[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43237023	+	chr22	43243520	+	.	0	9	7314947_1	17.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7314947_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43218001_43243001_416C;SPAN=6497;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:46 GQ:17.3 PL:[17.3, 0.0, 93.2] SR:9 DR:0 LR:-17.25 LO:20.3);ALT=C[chr22:43243520[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43243640	+	chr22	43253118	+	.	14	4	7314746_1	32.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=7314746_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43242501_43267501_154C;SPAN=9478;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:65 GQ:32 PL:[32.0, 0.0, 124.4] SR:4 DR:14 LR:-31.91 LO:35.06);ALT=T[chr22:43253118[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43308195	+	chr22	43411060	+	.	10	0	7315515_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7315515_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43308195(+)-22:43411060(-)__22_43389501_43414501D;SPAN=102865;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:42 GQ:21.8 PL:[21.8, 0.0, 77.9] SR:0 DR:10 LR:-21.63 LO:23.53);ALT=T[chr22:43411060[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43506839	+	chr22	43523697	+	.	21	0	7316070_1	61.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7316070_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43506839(+)-22:43523697(-)__22_43487501_43512501D;SPAN=16858;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:29 GQ:8.6 PL:[61.4, 0.0, 8.6] SR:0 DR:21 LR:-63.72 LO:63.72);ALT=C[chr22:43523697[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43506843	+	chr22	43520024	+	.	28	0	7316071_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7316071_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43506843(+)-22:43520024(-)__22_43487501_43512501D;SPAN=13181;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:28 LR:-89.12 LO:89.12);ALT=T[chr22:43520024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43520189	+	chr22	43523699	+	.	0	23	7315796_1	44.0	.	EVDNC=ASSMB;HOMSEQ=GCAG;MAPQ=60;MATEID=7315796_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43512001_43537001_106C;SPAN=3510;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:118 GQ:44 PL:[44.0, 0.0, 242.0] SR:23 DR:0 LR:-43.95 LO:51.84);ALT=G[chr22:43523699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43547662	+	chr22	43557055	+	.	45	0	7316166_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7316166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43547662(+)-22:43557055(-)__22_43536501_43561501D;SPAN=9393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:149 GQ:99 PL:[108.2, 0.0, 253.4] SR:0 DR:45 LR:-108.2 LO:111.4);ALT=G[chr22:43557055[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43547662	+	chr22	43555214	+	.	140	0	7316165_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7316165_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43547662(+)-22:43555214(-)__22_43536501_43561501D;SPAN=7552;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:140 DP:186 GQ:38.8 PL:[411.8, 0.0, 38.8] SR:0 DR:140 LR:-429.7 LO:429.7);ALT=G[chr22:43555214[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43555429	+	chr22	43557057	+	.	23	99	7316190_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGTA;MAPQ=60;MATEID=7316190_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43536501_43561501_168C;SPAN=1628;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:241 GQ:99 PL:[301.4, 0.0, 281.6] SR:99 DR:23 LR:-301.1 LO:301.1);ALT=A[chr22:43557057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43557197	+	chr22	43558808	+	.	12	39	7316197_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7316197_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_43536501_43561501_252C;SPAN=1611;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:129 GQ:99 PL:[130.1, 0.0, 182.9] SR:39 DR:12 LR:-130.1 LO:130.6);ALT=G[chr22:43558808[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	43749285	+	chr22	43750321	-	.	8	0	7316999_1	0	.	DISC_MAPQ=50;EVDNC=DSCRD;IMPRECISE;MAPQ=50;MATEID=7316999_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:43749285(+)-22:43750321(+)__22_43732501_43757501D;SPAN=1036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:122 GQ:6.3 PL:[0.0, 6.3, 306.9] SR:0 DR:8 LR:6.645 LO:13.98);ALT=T]chr22:43750321];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr22	44351478	+	chr22	44359165	+	.	23	9	7319390_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7319390_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44345001_44370001_410C;SPAN=7687;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:112 GQ:55.7 PL:[55.7, 0.0, 214.1] SR:9 DR:23 LR:-55.48 LO:60.85);ALT=G[chr22:44359165[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44351510	+	chr22	44360329	+	.	18	0	7319392_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7319392_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:44351510(+)-22:44360329(-)__22_44345001_44370001D;SPAN=8819;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:128 GQ:24.8 PL:[24.8, 0.0, 285.5] SR:0 DR:18 LR:-24.74 LO:37.75);ALT=G[chr22:44360329[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44359279	+	chr22	44360332	+	.	2	26	7319414_1	61.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GTG;MAPQ=60;MATEID=7319414_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44345001_44370001_19C;SPAN=1053;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:116 GQ:61.1 PL:[61.1, 0.0, 219.5] SR:26 DR:2 LR:-61.0 LO:66.08);ALT=G[chr22:44360332[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44360436	+	chr22	44364609	+	.	0	11	7319416_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AGGTA;MAPQ=60;MATEID=7319416_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44345001_44370001_345C;SPAN=4173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:107 GQ:7.4 PL:[7.4, 0.0, 251.6] SR:11 DR:0 LR:-7.322 LO:21.47);ALT=A[chr22:44364609[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44386287	+	chr22	44392216	+	.	0	24	7319623_1	50.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7319623_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44369501_44394501_347C;SPAN=5929;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:106 GQ:50.6 PL:[50.6, 0.0, 205.7] SR:24 DR:0 LR:-50.51 LO:55.87);ALT=G[chr22:44392216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44420276	+	chr22	44495931	+	.	14	0	7320209_1	35.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7320209_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:44420276(+)-22:44495931(-)__22_44492001_44517001D;SPAN=75655;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:41 GQ:35.3 PL:[35.3, 0.0, 61.7] SR:0 DR:14 LR:-35.11 LO:35.58);ALT=G[chr22:44495931[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44420331	+	chr22	44489807	+	.	39	22	7319655_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7319655_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44467501_44492501_36C;SPAN=69476;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:67 GQ:51.2 PL:[110.6, 0.0, 51.2] SR:22 DR:39 LR:-111.7 LO:111.7);ALT=G[chr22:44489807[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44496005	+	chr22	44514916	+	.	0	10	7320224_1	5.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=7320224_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44492001_44517001_73C;SPAN=18911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:102 GQ:5.6 PL:[5.6, 0.0, 239.9] SR:10 DR:0 LR:-5.376 LO:19.3);ALT=T[chr22:44514916[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44577728	+	chr22	44581685	+	.	8	0	7320170_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7320170_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:44577728(+)-22:44581685(-)__22_44565501_44590501D;SPAN=3957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:116 GQ:4.8 PL:[0.0, 4.8, 290.4] SR:0 DR:8 LR:5.019 LO:14.16);ALT=T[chr22:44581685[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44577798	+	chr22	44579197	+	.	20	32	7320171_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GG;MAPQ=60;MATEID=7320171_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44565501_44590501_410C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:43 DP:126 GQ:99 PL:[107.9, 0.0, 197.0] SR:32 DR:20 LR:-107.8 LO:109.3);ALT=G[chr22:44579197[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44579289	+	chr22	44581686	+	.	0	19	7320175_1	27.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7320175_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44565501_44590501_414C;SPAN=2397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:129 GQ:27.8 PL:[27.8, 0.0, 285.2] SR:19 DR:0 LR:-27.77 LO:40.26);ALT=G[chr22:44581686[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	44594602	+	chr22	44601636	+	.	0	7	7320625_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7320625_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_44590001_44615001_164C;SPAN=7034;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:102 GQ:4.2 PL:[0.0, 4.2, 254.1] SR:7 DR:0 LR:4.527 LO:12.38);ALT=G[chr22:44601636[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	45049189	+	chr22	45048157	+	.	31	0	7322063_1	69.0	.	DISC_MAPQ=21;EVDNC=DSCRD;IMPRECISE;MAPQ=21;MATEID=7322063_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:45048157(-)-22:45049189(+)__22_45031001_45056001D;SPAN=1032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:123 GQ:69.2 PL:[69.2, 0.0, 227.6] SR:0 DR:31 LR:-69.01 LO:73.83);ALT=]chr22:45049189]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	45504276	-	chr22	45505522	+	.	9	0	7323926_1	4.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7323926_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:45504276(-)-22:45505522(-)__22_45496501_45521501D;SPAN=1246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:93 GQ:4.7 PL:[4.7, 0.0, 219.2] SR:0 DR:9 LR:-4.513 LO:17.32);ALT=[chr22:45505522[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr22	45689195	+	chr22	45691441	+	.	5	5	7324763_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7324763_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_45668001_45693001_224C;SPAN=2246;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:7 DP:100 GQ:3.9 PL:[0.0, 3.9, 250.8] SR:5 DR:5 LR:3.985 LO:12.44);ALT=G[chr22:45691441[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	46068059	+	chr22	46085591	+	.	20	10	7326417_1	69.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7326417_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_46084501_46109501_180C;SPAN=17532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:47 GQ:43.4 PL:[69.8, 0.0, 43.4] SR:10 DR:20 LR:-70.1 LO:70.1);ALT=G[chr22:46085591[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	48793209	+	chr22	48792045	+	AAT	10	10	7336133_1	7.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AAT;MAPQ=60;MATEID=7336133_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_22_48779501_48804501_195C;SPAN=1164;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:118 GQ:7.7 PL:[7.7, 0.0, 278.3] SR:10 DR:10 LR:-7.643 LO:23.36);ALT=]chr22:48793209]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr22	50307493	+	chr22	50311911	+	.	8	2	7341386_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7341386_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_50298501_50323501_110C;SPAN=4418;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:95 GQ:0.8 PL:[0.8, 0.0, 228.5] SR:2 DR:8 LR:-0.6702 LO:14.89);ALT=T[chr22:50311911[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	50319205	+	chr22	50320902	+	.	2	12	7341432_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7341432_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_50298501_50323501_29C;SPAN=1697;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:97 GQ:16.7 PL:[16.7, 0.0, 218.0] SR:12 DR:2 LR:-16.63 LO:26.97);ALT=G[chr22:50320902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	50624455	+	chr22	50631472	+	.	37	0	7342490_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7342490_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:50624455(+)-22:50631472(-)__22_50617001_50642001D;SPAN=7017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:60 GQ:39.8 PL:[105.8, 0.0, 39.8] SR:0 DR:37 LR:-107.5 LO:107.5);ALT=C[chr22:50631472[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	50624464	+	chr22	50632713	+	.	24	0	7342491_1	64.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7342491_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=22:50624464(+)-22:50632713(-)__22_50617001_50642001D;SPAN=8249;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:56 GQ:64.1 PL:[64.1, 0.0, 70.7] SR:0 DR:24 LR:-64.05 LO:64.08);ALT=G[chr22:50632713[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr22	50965714	+	chr22	50968333	+	.	4	2	7343958_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7343958_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_22_50960001_50985001_401C;SPAN=2619;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:73 GQ:6.3 PL:[0.0, 6.3, 188.1] SR:2 DR:4 LR:6.574 LO:6.671);ALT=T[chr22:50968333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	14883691	+	chrX	14891105	+	.	9	0	7369390_1	14.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7369390_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:14883691(+)-23:14891105(-)__23_14871501_14896501D;SPAN=7414;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:55 GQ:14.9 PL:[14.9, 0.0, 117.2] SR:0 DR:9 LR:-14.81 LO:19.52);ALT=A[chrX:14891105[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	15756524	+	chrX	15768091	+	.	37	0	7370718_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7370718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:15756524(+)-23:15768091(-)__23_15753501_15778501D;SPAN=11567;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:37 DP:68 GQ:60.8 PL:[103.7, 0.0, 60.8] SR:0 DR:37 LR:-104.3 LO:104.3);ALT=A[chrX:15768091[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	15768288	+	chrX	15780904	+	.	0	10	7370739_1	23.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=7370739_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_15753501_15778501_196C;SPAN=12616;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:35 GQ:23.6 PL:[23.6, 0.0, 59.9] SR:10 DR:0 LR:-23.53 LO:24.46);ALT=T[chrX:15780904[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19362213	+	chrX	19367429	+	.	14	14	7376372_1	43.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=7376372_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_23_19355001_19380001_68C;SPAN=5216;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:14 DR:14 LR:-43.7 LO:44.82);ALT=G[chrX:19367429[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19362213	+	chrX	19368053	+	CAAGCAGAGTGCTGGTAGCATCCCGTAATTTTGCAAATGATGCTACATTTGAAATTA	9	23	7376373_1	73.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=CAAGCAGAGTGCTGGTAGCATCCCGTAATTTTGCAAATGATGCTACATTTGAAATTA;MAPQ=60;MATEID=7376373_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_19355001_19380001_68C;SPAN=5840;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:57 GQ:63.8 PL:[73.7, 0.0, 63.8] SR:23 DR:9 LR:-73.72 LO:73.72);ALT=G[chrX:19368053[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19560311	+	chrX	19564037	+	.	4	3	7376651_1	1.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CAC;MAPQ=60;MATEID=7376651_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=CACA;SCTG=c_23_19551001_19576001_202C;SPAN=3726;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:3 DR:4 LR:-1.062 LO:9.396);ALT=C[chrX:19564037[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19626165	+	chrX	19649981	+	.	5	15	7376914_1	59.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7376914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19649001_19674001_64C;SPAN=23816;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:20 DP:25 GQ:0 PL:[59.4, 0.0, 0.0] SR:15 DR:5 LR:-62.61 LO:62.61);ALT=T[chrX:19649981[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19650076	+	chrX	19663517	+	.	0	11	7376917_1	16.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7376917_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19649001_19674001_286C;SPAN=13441;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:74 GQ:16.4 PL:[16.4, 0.0, 161.6] SR:11 DR:0 LR:-16.26 LO:23.36);ALT=C[chrX:19663517[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19663595	+	chrX	19701941	+	.	11	5	7377006_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7377006_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19698001_19723001_62C;SPAN=38346;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:26 GQ:26 PL:[35.9, 0.0, 26.0] SR:5 DR:11 LR:-35.93 LO:35.93);ALT=T[chrX:19701941[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19702146	+	chrX	19713728	+	.	2	8	7377014_1	15.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AC;MAPQ=60;MATEID=7377014_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19698001_19723001_249C;SPAN=11582;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:53 GQ:15.5 PL:[15.5, 0.0, 111.2] SR:8 DR:2 LR:-15.35 LO:19.68);ALT=C[chrX:19713728[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19764559	+	chrX	19854242	+	.	3	4	7377280_1	16.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7377280_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19845001_19870001_251C;SPAN=89683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:24 GQ:16.7 PL:[16.7, 0.0, 39.8] SR:4 DR:3 LR:-16.6 LO:17.2);ALT=C[chrX:19854242[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	19854401	+	chrX	19905425	+	.	41	67	7377322_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7377322_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_19894001_19919001_262C;SPAN=51024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:28 GQ:22.8 PL:[250.8, 22.8, 0.0] SR:67 DR:41 LR:-250.9 LO:250.9);ALT=C[chrX:19905425[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	20174369	+	chrX	20179761	+	.	2	2	7377801_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=7377801_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_20163501_20188501_75C;SPAN=5392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:56 GQ:1.8 PL:[0.0, 1.8, 138.6] SR:2 DR:2 LR:1.968 LO:7.145);ALT=T[chrX:20179761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	46696639	+	chrX	46712909	+	.	7	7	7413853_1	22.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=7413853_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_46697001_46722001_7C;SPAN=16270;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:28 GQ:22.1 PL:[22.1, 0.0, 45.2] SR:7 DR:7 LR:-22.12 LO:22.58);ALT=T[chrX:46712909[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47002145	+	chrX	47003872	+	.	0	111	7414510_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=7414510_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_46991001_47016001_144C;SPAN=1727;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:111 DP:139 GQ:8.6 PL:[328.7, 0.0, 8.6] SR:111 DR:0 LR:-347.3 LO:347.3);ALT=T[chrX:47003872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47053423	+	chrX	47058201	+	.	0	10	7414354_1	18.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7414354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_47040001_47065001_192C;SPAN=4778;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:53 GQ:18.8 PL:[18.8, 0.0, 107.9] SR:10 DR:0 LR:-18.65 LO:22.38);ALT=G[chrX:47058201[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47072580	+	chrX	47073723	+	.	2	4	7414447_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7414447_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_47064501_47089501_93C;SPAN=1143;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:61 GQ:0.2 PL:[0.2, 0.0, 145.4] SR:4 DR:2 LR:0.0214 LO:9.242);ALT=G[chrX:47073723[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47104883	+	chrX	47106470	+	.	3	3	7414657_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=7414657_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_47089001_47114001_32C;SPAN=1587;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:54 GQ:1.2 PL:[0.0, 1.2, 132.0] SR:3 DR:3 LR:1.426 LO:7.211);ALT=T[chrX:47106470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47420689	+	chrX	47422623	+	.	8	0	7415494_1	8.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415494_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47420689(+)-23:47422623(-)__23_47407501_47432501D;SPAN=1934;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:68 GQ:8 PL:[8.0, 0.0, 156.5] SR:0 DR:8 LR:-7.985 LO:16.11);ALT=C[chrX:47422623[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47420691	+	chrX	47422305	+	.	10	0	7415495_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415495_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47420691(+)-23:47422305(-)__23_47407501_47432501D;SPAN=1614;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:71 GQ:14 PL:[14.0, 0.0, 155.9] SR:0 DR:10 LR:-13.77 LO:20.98);ALT=G[chrX:47422305[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47422728	+	chrX	47424195	+	.	0	6	7415501_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7415501_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_47407501_47432501_234C;SPAN=1467;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:72 GQ:0.5 PL:[0.5, 0.0, 172.1] SR:6 DR:0 LR:-0.2994 LO:11.14);ALT=G[chrX:47424195[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47441921	+	chrX	47444333	+	.	82	0	7415622_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7415622_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47441921(+)-23:47444333(-)__23_47432001_47457001D;SPAN=2412;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:82 DP:116 GQ:41.3 PL:[239.3, 0.0, 41.3] SR:0 DR:82 LR:-247.1 LO:247.1);ALT=G[chrX:47444333[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47441924	+	chrX	47444601	+	.	35	0	7415624_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415624_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47441924(+)-23:47444601(-)__23_47432001_47457001D;SPAN=2677;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:97 GQ:89.3 PL:[89.3, 0.0, 145.4] SR:0 DR:35 LR:-89.26 LO:90.01);ALT=T[chrX:47444601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47442935	+	chrX	47444334	+	.	7	108	7415627_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7415627_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_47432001_47457001_303C;SPAN=1399;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:115 DP:146 GQ:13.4 PL:[340.1, 0.0, 13.4] SR:108 DR:7 LR:-358.1 LO:358.1);ALT=G[chrX:47444334[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47483839	+	chrX	47485456	+	.	6	81	7415530_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7415530_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_47481001_47506001_222C;SPAN=1617;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:85 DP:88 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:81 DR:6 LR:-260.8 LO:260.8);ALT=C[chrX:47485456[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47487679	+	chrX	47488921	+	.	0	50	7415541_1	99.0	.	EVDNC=ASSMB;HOMSEQ=ACCTG;MAPQ=60;MATEID=7415541_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_47481001_47506001_19C;SPAN=1242;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:68 GQ:17.9 PL:[146.6, 0.0, 17.9] SR:50 DR:0 LR:-152.4 LO:152.4);ALT=G[chrX:47488921[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47487972	+	chrX	47488982	+	.	51	0	7415543_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7415543_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47487972(+)-23:47488982(-)__23_47481001_47506001D;SPAN=1010;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:94 GQ:83.6 PL:[143.0, 0.0, 83.6] SR:0 DR:51 LR:-143.7 LO:143.7);ALT=G[chrX:47488982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47511543	+	chrX	47516971	+	TCTGTGAGGAGAGAGCTCTTACGATCAATGAACTTGAGAGCTTCTGCCAGTGTCAACTCCAGGAAAAAACCATATCCCAGGGCCACATAGATGCGTGAAGTATCTGGG	0	225	7415818_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCTGTGAGGAGAGAGCTCTTACGATCAATGAACTTGAGAGCTTCTGCCAGTGTCAACTCCAGGAAAAAACCATATCCCAGGGCCACATAGATGCGTGAAGTATCTGGG;MAPQ=60;MATEID=7415818_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_47505501_47530501_216C;SPAN=5428;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:225 DP:155 GQ:60.7 PL:[666.7, 60.7, 0.0] SR:225 DR:0 LR:-666.8 LO:666.8);ALT=C[chrX:47516971[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47516740	+	chrX	47518290	+	.	16	0	7415827_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415827_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47516740(+)-23:47518290(-)__23_47505501_47530501D;SPAN=1550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:16 DP:102 GQ:25.4 PL:[25.4, 0.0, 220.1] SR:0 DR:16 LR:-25.18 LO:34.39);ALT=A[chrX:47518290[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47517076	+	chrX	47518512	+	.	9	0	7415833_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415833_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47517076(+)-23:47518512(-)__23_47505501_47530501D;SPAN=1436;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:90 GQ:5.3 PL:[5.3, 0.0, 213.2] SR:0 DR:9 LR:-5.326 LO:17.45);ALT=G[chrX:47518512[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	47517090	+	chrX	47518288	+	.	55	0	7415834_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7415834_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:47517090(+)-23:47518288(-)__23_47505501_47530501D;SPAN=1198;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:55 DP:97 GQ:79.4 PL:[155.3, 0.0, 79.4] SR:0 DR:55 LR:-156.6 LO:156.6);ALT=G[chrX:47518288[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48134218	+	chrX	48037219	+	.	14	0	7416735_1	38.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=7416735_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48037219(-)-23:48134218(+)__23_48118001_48143001D;SPAN=96999;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:30 GQ:34.7 PL:[38.0, 0.0, 34.7] SR:0 DR:14 LR:-38.09 LO:38.09);ALT=]chrX:48134218]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	48104326	+	chrX	52641761	+	.	8	0	7424166_1	14.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=7424166_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48104326(+)-23:52641761(-)__23_52626001_52651001D;SPAN=4537435;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:44 GQ:14.6 PL:[14.6, 0.0, 90.5] SR:0 DR:8 LR:-14.49 LO:17.76);ALT=G[chrX:52641761[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48140638	+	chrX	52641929	+	.	17	0	7424168_1	45.0	.	DISC_MAPQ=48;EVDNC=DSCRD;IMPRECISE;MAPQ=48;MATEID=7424168_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48140638(+)-23:52641929(-)__23_52626001_52651001D;SPAN=4501291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:39 GQ:45.5 PL:[45.5, 0.0, 48.8] SR:0 DR:17 LR:-45.55 LO:45.56);ALT=A[chrX:52641929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	52642052	+	chrX	48140756	+	.	9	0	7424169_1	20.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=7424169_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48140756(-)-23:52642052(+)__23_52626001_52651001D;SPAN=4501296;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:34 GQ:20.6 PL:[20.6, 0.0, 60.2] SR:0 DR:9 LR:-20.5 LO:21.66);ALT=]chrX:52642052]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	48326315	+	chrX	48327722	+	.	4	3	7417270_1	0	.	DISC_MAPQ=53;EVDNC=TSI_L;HOMSEQ=CCTG;MAPQ=60;MATEID=7417270_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_48314001_48339001_248C;SPAN=1407;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:60 GQ:0.2 PL:[0.2, 0.0, 145.4] SR:3 DR:4 LR:-0.2495 LO:9.28);ALT=G[chrX:48327722[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48334784	+	chrX	48336347	+	.	0	8	7417290_1	10.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=7417290_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48314001_48339001_37C;SPAN=1563;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:59 GQ:10.4 PL:[10.4, 0.0, 132.5] SR:8 DR:0 LR:-10.42 LO:16.64);ALT=G[chrX:48336347[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48380297	+	chrX	48382086	+	.	60	3	7417402_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GGT;MAPQ=60;MATEID=7417402_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48363001_48388001_60C;SPAN=1789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:60 DP:74 GQ:0 PL:[178.2, 0.0, 0.0] SR:3 DR:60 LR:-188.7 LO:188.7);ALT=T[chrX:48382086[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48432986	+	chrX	48434699	+	.	13	0	7417797_1	15.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7417797_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48432986(+)-23:48434699(-)__23_48412001_48437001D;SPAN=1713;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:0 DR:13 LR:-15.01 LO:26.61);ALT=C[chrX:48434699[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48433671	+	chrX	48434701	+	.	0	8	7417800_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7417800_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48412001_48437001_80C;SPAN=1030;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:170 GQ:19.6 PL:[0.0, 19.6, 452.2] SR:8 DR:0 LR:19.65 LO:12.8);ALT=G[chrX:48434701[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48455999	+	chrX	48457102	+	.	10	0	7417545_1	17.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7417545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48455999(+)-23:48457102(-)__23_48436501_48461501D;SPAN=1103;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:58 GQ:17.3 PL:[17.3, 0.0, 122.9] SR:0 DR:10 LR:-17.3 LO:21.94);ALT=G[chrX:48457102[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48542414	+	chrX	48543932	+	.	9	0	7417693_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7417693_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48542414(+)-23:48543932(-)__23_48534501_48559501D;SPAN=1518;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:65 GQ:12.2 PL:[12.2, 0.0, 144.2] SR:0 DR:9 LR:-12.1 LO:18.81);ALT=T[chrX:48543932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48547823	+	chrX	48549497	+	.	2	7	7417706_1	10.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7417706_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48534501_48559501_191C;SPAN=1674;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:61 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:7 DR:2 LR:-9.882 LO:16.52);ALT=G[chrX:48549497[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48751525	+	chrX	48755006	+	.	14	0	7418345_1	27.0	.	DISC_MAPQ=46;EVDNC=DSCRD;IMPRECISE;MAPQ=46;MATEID=7418345_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48751525(+)-23:48755006(-)__23_48730501_48755501D;SPAN=3481;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:71 GQ:27.2 PL:[27.2, 0.0, 142.7] SR:0 DR:14 LR:-26.98 LO:31.63);ALT=G[chrX:48755006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48752420	+	chrX	48755006	+	.	10	0	7418350_1	14.0	.	DISC_MAPQ=18;EVDNC=DSCRD;IMPRECISE;MAPQ=18;MATEID=7418350_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48752420(+)-23:48755006(-)__23_48730501_48755501D;SPAN=2586;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:67 GQ:14.9 PL:[14.9, 0.0, 146.9] SR:0 DR:10 LR:-14.86 LO:21.25);ALT=G[chrX:48755006[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48755369	+	chrX	48758465	+	.	23	0	7418360_1	67.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7418360_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48755369(+)-23:48758465(-)__23_48730501_48755501D;SPAN=3096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:31 GQ:5 PL:[67.7, 0.0, 5.0] SR:0 DR:23 LR:-70.29 LO:70.29);ALT=A[chrX:48758465[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48755859	+	chrX	48758466	+	.	0	26	7418260_1	68.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7418260_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48755001_48780001_169C;SPAN=2607;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:26 DP:64 GQ:68.6 PL:[68.6, 0.0, 85.1] SR:26 DR:0 LR:-68.49 LO:68.61);ALT=G[chrX:48758466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48847525	+	chrX	48849840	+	.	2	4	7418443_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=7418443_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_23_48828501_48853501_279C;SPAN=2315;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:64 GQ:0.6 PL:[0.0, 0.6, 155.1] SR:4 DR:2 LR:0.8342 LO:9.134);ALT=G[chrX:48849840[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48853832	+	chrX	48858597	+	.	10	0	7418576_1	16.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7418576_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:48853832(+)-23:48858597(-)__23_48853001_48878001D;SPAN=4765;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:60 GQ:16.7 PL:[16.7, 0.0, 128.9] SR:0 DR:10 LR:-16.75 LO:21.78);ALT=A[chrX:48858597[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	48930310	+	chrX	48931466	+	.	0	9	7419079_1	16.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=7419079_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_48926501_48951501_290C;SPAN=1156;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:51 GQ:16.1 PL:[16.1, 0.0, 105.2] SR:9 DR:0 LR:-15.89 LO:19.85);ALT=C[chrX:48931466[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49028443	+	chrX	49029476	+	.	102	154	7418806_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;MAPQ=60;MATEID=7418806_2;MATENM=0;NM=0;NUMPARTS=4;REPSEQ=TATTAT;SCTG=c_23_49024501_49049501_63C;SPAN=1033;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:225 DP:175 GQ:60.5 PL:[525.3, 60.5, 0.0] SR:154 DR:102 LR:-525.4 LO:525.4);ALT=T[chrX:49029476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49028443	+	chrX	49031020	+	ATATTATGCCTGGTGATCCTGATCTGCTTCAGTGCCTCCACACCAGGCTACTCCTCCCTGTCGGTGATTGAGATGATCCTTGCTGCTATTTTCTTTGTTGTCTACATGTGTGACCTGCACACCAAGATACCATTCATCAACTGGCCCTGGAGTGATTTCTTCCGAACCCTCATAGCGGCAATCCTCTACCTGATCACCTCCATTGTTGTCCTTGTTGAGAGAGGAAACCACTCCAAAATCGTCGCAGGGGTACTGGGCCTAATCGCTACGTGCCTCTTTGGCTATGATGCCTATGTCACCTTCCCCGTTCGGCAGCCAAGACATACAGCAGCCCCCACT	0	189	7418807_1	99.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=G;INSERTION=ATATTATGCCTGGTGATCCTGATCTGCTTCAGTGCCTCCACACCAGGCTACTCCTCCCTGTCGGTGATTGAGATGATCCTTGCTGCTATTTTCTTTGTTGTCTACATGTGTGACCTGCACACCAAGATACCATTCATCAACTGGCCCTGGAGTGATTTCTTCCGAACCCTCATAGCGGCAATCCTCTACCTGATCACCTCCATTGTTGTCCTTGTTGAGAGAGGAAACCACTCCAAAATCGTCGCAGGGGTACTGGGCCTAATCGCTACGTGCCTCTTTGGCTATGATGCCTATGTCACCTTCCCCGTTCGGCAGCCAAGACATACAGCAGCCCCCACT;MAPQ=60;MATEID=7418807_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_49024501_49049501_63C;SPAN=2577;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:189 DP:117 GQ:51.1 PL:[561.1, 51.1, 0.0] SR:189 DR:0 LR:-561.1 LO:561.1);ALT=T[chrX:49031020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49029881	+	chrX	49031019	+	.	12	0	7418813_1	25.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=7418813_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:49029881(+)-23:49031019(-)__23_49024501_49049501D;SPAN=1138;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=C[chrX:49031019[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	49092147	+	chrX	49093553	+	.	0	12	7418928_1	22.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7418928_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_49073501_49098501_13C;SPAN=1406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:64 GQ:22.4 PL:[22.4, 0.0, 131.3] SR:12 DR:0 LR:-22.27 LO:26.82);ALT=G[chrX:49093553[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	50870275	-	chrX	50871316	+	.	12	0	7421640_1	25.0	.	DISC_MAPQ=31;EVDNC=DSCRD;IMPRECISE;MAPQ=31;MATEID=7421640_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:50870275(-)-23:50871316(-)__23_50862001_50887001D;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:52 GQ:25.7 PL:[25.7, 0.0, 98.3] SR:0 DR:12 LR:-25.52 LO:28.05);ALT=[chrX:50871316[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	51279677	+	chrX	51966036	-	.	32	0	7423313_1	86.0	.	DISC_MAPQ=33;EVDNC=DSCRD;IMPRECISE;MAPQ=33;MATEID=7423313_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:51279677(+)-23:51966036(+)__23_51964501_51989501D;SPAN=686359;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:32 DP:72 GQ:86.3 PL:[86.3, 0.0, 86.3] SR:0 DR:32 LR:-86.13 LO:86.13);ALT=C]chrX:51966036];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	53442119	+	chrX	53449439	+	.	0	14	7425589_1	25.0	.	EVDNC=ASSMB;HOMSEQ=ACC;MAPQ=60;MATEID=7425589_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_53434501_53459501_60C;SPAN=7320;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:78 GQ:25.1 PL:[25.1, 0.0, 163.7] SR:14 DR:0 LR:-25.08 LO:30.99);ALT=C[chrX:53449439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	53459359	+	chrX	53460667	+	.	0	42	7425679_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AC;MAPQ=60;MATEID=7425679_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_53459001_53484001_138C;SPAN=1308;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:42 DP:70 GQ:50.3 PL:[119.6, 0.0, 50.3] SR:42 DR:0 LR:-121.2 LO:121.2);ALT=C[chrX:53460667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	53459404	+	chrX	53461264	+	.	44	0	7425680_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7425680_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:53459404(+)-23:53461264(-)__23_53459001_53484001D;SPAN=1860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:76 GQ:58.7 PL:[124.7, 0.0, 58.7] SR:0 DR:44 LR:-125.9 LO:125.9);ALT=C[chrX:53461264[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	54466927	+	chrX	54469831	+	.	18	0	7427615_1	39.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7427615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:54466927(+)-23:54469831(-)__23_54463501_54488501D;SPAN=2904;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:73 GQ:39.8 PL:[39.8, 0.0, 135.5] SR:0 DR:18 LR:-39.64 LO:42.67);ALT=G[chrX:54469831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	54466934	+	chrX	54470438	+	.	10	0	7427617_1	14.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7427617_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:54466934(+)-23:54470438(-)__23_54463501_54488501D;SPAN=3504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:68 GQ:14.6 PL:[14.6, 0.0, 149.9] SR:0 DR:10 LR:-14.59 LO:21.18);ALT=A[chrX:54470438[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	54467213	+	chrX	54470439	+	CTGACTTGGAGCTAGATGAGGTGGAAGACTTCCTTGGAGAGCTGTTGACCAACGAGTTTGATACAGTTGTGGAAGACGGGAGTCTGCCCC	0	35	7427621_1	98.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AGGTGAGC;INSERTION=CTGACTTGGAGCTAGATGAGGTGGAAGACTTCCTTGGAGAGCTGTTGACCAACGAGTTTGATACAGTTGTGGAAGACGGGAGTCTGCCCC;MAPQ=60;MATEID=7427621_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_54463501_54488501_254C;SPAN=3226;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:35 DP:62 GQ:49.4 PL:[98.9, 0.0, 49.4] SR:35 DR:0 LR:-99.53 LO:99.53);ALT=G[chrX:54470439[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	54751766	-	chrX	54752835	+	.	8	0	7428194_1	11.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7428194_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:54751766(-)-23:54752835(-)__23_54733001_54758001D;SPAN=1069;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:0 DR:8 LR:-11.51 LO:16.91);ALT=[chrX:54752835[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	54834898	+	chrX	54836151	+	.	12	0	7428273_1	25.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7428273_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:54834898(+)-23:54836151(-)__23_54831001_54856001D;SPAN=1253;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:53 GQ:25.4 PL:[25.4, 0.0, 101.3] SR:0 DR:12 LR:-25.25 LO:27.93);ALT=C[chrX:54836151[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70129274	-	chrX	70140010	+	.	42	0	7444682_1	99.0	.	DISC_MAPQ=52;EVDNC=DSCRD;IMPRECISE;MAPQ=52;MATEID=7444682_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:70129274(-)-23:70140010(-)__23_70119001_70144001D;SPAN=10736;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:39 GQ:11.1 PL:[122.1, 11.1, 0.0] SR:0 DR:42 LR:-122.1 LO:122.1);ALT=[chrX:70140010[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	70129420	+	chrX	70137257	-	.	2	26	7444683_1	79.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=7444683_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_70119001_70144001_29C;SPAN=7837;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:49 GQ:39.5 PL:[79.1, 0.0, 39.5] SR:26 DR:2 LR:-79.86 LO:79.86);ALT=T]chrX:70137257];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	70282800	+	chrX	70287992	+	.	0	9	7445002_1	14.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7445002_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_70266001_70291001_188C;SPAN=5192;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:55 GQ:14.9 PL:[14.9, 0.0, 117.2] SR:9 DR:0 LR:-14.81 LO:19.52);ALT=C[chrX:70287992[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70329240	+	chrX	70330354	+	AGTCCAGCTGTGGTCCCAGTCAGTCCGGTACTGCACCAAGTGCTCCAAACAGTGGTTCAAGAATCTGTTGTTCCAGTTCAGTTCTAGCTGGGATTCACTCAGTTTGTGAAGTGTTAGGTTCTCTGGAGCCCAGGGGATCA	0	9	7445235_1	16.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGTCCAGCTGTGGTCCCAGTCAGTCCGGTACTGCACCAAGTGCTCCAAACAGTGGTTCAAGAATCTGTTGTTCCAGTTCAGTTCTAGCTGGGATTCACTCAGTTTGTGAAGTGTTAGGTTCTCTGGAGCCCAGGGGATCA;MAPQ=60;MATEID=7445235_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_70315001_70340001_297C;SPAN=1114;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:9 DR:0 LR:-16.43 LO:20.02);ALT=C[chrX:70330354[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70503594	+	chrX	70510476	+	.	41	0	7445461_1	99.0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=7445461_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:70503594(+)-23:70510476(-)__23_70486501_70511501D;SPAN=6882;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:45 GQ:12 PL:[132.0, 12.0, 0.0] SR:0 DR:41 LR:-132.0 LO:132.0);ALT=T[chrX:70510476[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70753065	+	chrX	70756024	+	.	8	0	7446178_1	5.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7446178_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:70753065(+)-23:70756024(-)__23_70731501_70756501D;SPAN=2959;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:79 GQ:5 PL:[5.0, 0.0, 186.5] SR:0 DR:8 LR:-5.005 LO:15.56);ALT=A[chrX:70756024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	70787966	+	chrX	70793470	+	.	3	6	7446024_1	11.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=7446024_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_70780501_70805501_212C;SPAN=5504;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:57 GQ:11 PL:[11.0, 0.0, 126.5] SR:6 DR:3 LR:-10.97 LO:16.77);ALT=A[chrX:70793470[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	71493837	+	chrX	71494902	+	.	9	0	7447670_1	15.0	.	DISC_MAPQ=45;EVDNC=DSCRD;IMPRECISE;MAPQ=45;MATEID=7447670_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:71493837(+)-23:71494902(-)__23_71491001_71516001D;SPAN=1065;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:54 GQ:15.2 PL:[15.2, 0.0, 114.2] SR:0 DR:9 LR:-15.08 LO:19.6);ALT=G[chrX:71494902[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	71788736	+	chrX	71792500	+	CATCTGCTTATGCAGTGCATATGCTTCAATCAAAGAATGCACCATACTGG	0	10	7447909_1	17.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=CATCTGCTTATGCAGTGCATATGCTTCAATCAAAGAATGCACCATACTGG;MAPQ=60;MATEID=7447909_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_71785001_71810001_149C;SPAN=3764;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:56 GQ:17.9 PL:[17.9, 0.0, 116.9] SR:10 DR:0 LR:-17.84 LO:22.11);ALT=T[chrX:71792500[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	73164337	+	chrX	73166831	+	.	15	0	7449789_1	32.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7449789_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:73164337(+)-23:73166831(-)__23_73157001_73182001D;SPAN=2494;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:62 GQ:32.9 PL:[32.9, 0.0, 115.4] SR:0 DR:15 LR:-32.72 LO:35.42);ALT=C[chrX:73166831[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	74273422	+	chrX	74282163	+	GATCCAAGACAATGATTTCATCTGCATCAACCACTGTTGACAATCTGTGTGCAATGAAAATAGAAGTTCTGTGTTTGACCACATCCTTCATGGCACCAAGAATAGT	4	11	7451295_1	30.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=GATCCAAGACAATGATTTCATCTGCATCAACCACTGTTGACAATCTGTGTGCAATGAAAATAGAAGTTCTGTGTTTGACCACATCCTTCATGGCACCAAGAATAGT;MAPQ=60;MATEID=7451295_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_74259501_74284501_216C;SPAN=8741;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:58 GQ:30.5 PL:[30.5, 0.0, 109.7] SR:11 DR:4 LR:-30.5 LO:33.04);ALT=T[chrX:74282163[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	74332809	+	chrX	74334588	+	.	0	9	7451544_1	23.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7451544_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_74333001_74358001_22C;SPAN=1779;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:9 DR:0 LR:-23.21 LO:23.34);ALT=T[chrX:74334588[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	74332854	+	chrX	74376054	+	.	8	0	7451448_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7451448_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:74332854(+)-23:74376054(-)__23_74357501_74382501D;SPAN=43200;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:40 GQ:15.5 PL:[15.5, 0.0, 81.5] SR:0 DR:8 LR:-15.57 LO:18.13);ALT=C[chrX:74376054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	74334672	+	chrX	74375940	+	.	0	14	7451547_1	37.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7451547_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_74333001_74358001_225C;SPAN=41268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:32 GQ:37.7 PL:[37.7, 0.0, 37.7] SR:14 DR:0 LR:-37.54 LO:37.55);ALT=G[chrX:74375940[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	75393005	+	chrX	75395306	+	TTCCGGGGAGTTGGTGTCTGTGGCACATGCGCTTTCTCTCCCAGCAGAGTCGTATGGCAACGATCCTGACATTGAGATGGCTTGGGCCATGAGAGCAATGCAGCATGCTGAAGTCTATTACA	9	13	7452735_1	54.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TTCCGGGGAGTTGGTGTCTGTGGCACATGCGCTTTCTCTCCCAGCAGAGTCGTATGGCAACGATCCTGACATTGAGATGGCTTGGGCCATGAGAGCAATGCAGCATGCTGAAGTCTATTACA;MAPQ=60;MATEID=7452735_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_75386501_75411501_132C;SPAN=2301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:54 GQ:54.8 PL:[54.8, 0.0, 74.6] SR:13 DR:9 LR:-54.69 LO:54.89);ALT=T[chrX:75395306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77121417	+	chrX	77123867	+	.	70	27	7455196_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=CTCACGCCTGTAATCCCAGCACTTTGGGAGGC;MAPQ=60;MATEID=7455196_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_77101501_77126501_63C;SPAN=2450;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:91 DP:20 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:27 DR:70 LR:-267.4 LO:267.4);ALT=C[chrX:77123867[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77155090	+	chrX	77160681	+	TTCGAAGCATTCAGCAAACAATGGCAAGGCAGAGCCACCAGAAACGTACACCTGATTTTCATGACAAATACGGTAATGCTGTATTAGCTAGTGGAGCCACTTTCTGTATTGTTACATGGACATAT	28	203	7455259_1	99.0	.	DISC_MAPQ=57;EVDNC=TSI_G;HOMSEQ=GTA;INSERTION=TTCGAAGCATTCAGCAAACAATGGCAAGGCAGAGCCACCAGAAACGTACACCTGATTTTCATGACAAATACGGTAATGCTGTATTAGCTAGTGGAGCCACTTTCTGTATTGTTACATGGACATAT;MAPQ=60;MATEID=7455259_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_77150501_77175501_297C;SPAN=5591;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:221 DP:105 GQ:59.5 PL:[653.5, 59.5, 0.0] SR:203 DR:28 LR:-653.6 LO:653.6);ALT=G[chrX:77160681[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77155090	+	chrX	77158137	+	.	80	45	7455258_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AAG;MAPQ=60;MATEID=7455258_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_77150501_77175501_297C;SPAN=3047;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:86 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:45 DR:80 LR:-333.4 LO:333.4);ALT=G[chrX:77158137[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77359865	+	chrX	77369238	+	.	45	0	7455545_1	99.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7455545_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:77359865(+)-23:77369238(-)__23_77346501_77371501D;SPAN=9373;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:97 GQ:99 PL:[122.3, 0.0, 112.4] SR:0 DR:45 LR:-122.3 LO:122.3);ALT=G[chrX:77369238[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77378870	+	chrX	77380369	+	.	11	0	7455778_1	17.0	.	DISC_MAPQ=27;EVDNC=DSCRD;IMPRECISE;MAPQ=27;MATEID=7455778_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:77378870(+)-23:77380369(-)__23_77371001_77396001D;SPAN=1499;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:68 GQ:17.9 PL:[17.9, 0.0, 146.6] SR:0 DR:11 LR:-17.89 LO:23.8);ALT=T[chrX:77380369[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77529272	+	chrX	77538950	+	.	0	8	7455999_1	12.0	.	EVDNC=ASSMB;HOMSEQ=CCT;MAPQ=60;MATEID=7455999_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_77518001_77543001_196C;SPAN=9678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.59 LO:17.19);ALT=T[chrX:77538950[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	77539040	+	chrX	77582802	+	.	0	18	7456009_1	52.0	.	EVDNC=ASSMB;HOMSEQ=CTG;MAPQ=60;MATEID=7456009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_77518001_77543001_125C;SPAN=43762;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:26 GQ:9.5 PL:[52.4, 0.0, 9.5] SR:18 DR:0 LR:-53.93 LO:53.93);ALT=G[chrX:77582802[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	106871845	+	chrX	106882523	+	.	8	0	7492757_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7492757_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:106871845(+)-23:106882523(-)__23_106869001_106894001D;SPAN=10678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:56 GQ:11.3 PL:[11.3, 0.0, 123.5] SR:0 DR:8 LR:-11.24 LO:16.84);ALT=G[chrX:106882523[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	106890999	+	chrX	106893168	+	.	2	2	7492791_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTGA;MAPQ=60;MATEID=7492791_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_106869001_106894001_221C;SPAN=2169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:62 GQ:3.3 PL:[0.0, 3.3, 155.1] SR:2 DR:2 LR:3.593 LO:6.963);ALT=A[chrX:106893168[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	106957980	+	chrX	106959920	+	ATGGCCTGTTCGATCTTGTTGTCTATGGCCACCACGCTGGCTCCGGAGGCA	65	165	7492976_1	99.0	.	DISC_MAPQ=59;EVDNC=TSI_G;HOMSEQ=CTG;INSERTION=ATGGCCTGTTCGATCTTGTTGTCTATGGCCACCACGCTGGCTCCGGAGGCA;MAPQ=60;MATEID=7492976_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_106942501_106967501_92C;SPAN=1940;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:198 DP:123 GQ:53.5 PL:[587.5, 53.5, 0.0] SR:165 DR:65 LR:-587.5 LO:587.5);ALT=C[chrX:106959920[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	108780694	+	chrX	108784702	+	.	10	0	7495197_1	29.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7495197_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:108780694(+)-23:108784702(-)__23_108755501_108780501D;SPAN=4008;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:10 DP:0 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:0 DR:10 LR:-29.71 LO:29.71);ALT=T[chrX:108784702[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	114398129	+	chrX	114201840	+	TCTCATACC	0	28	7502543_1	89.0	.	EVDNC=ASSMB;INSERTION=TCTCATACC;MAPQ=60;MATEID=7502543_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_114390501_114415501_164C;SPAN=196289;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:28 DP:30 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:28 DR:0 LR:-89.12 LO:89.12);ALT=]chrX:114398129]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chrX	122840848	+	chrX	122866812	+	.	24	0	7515961_1	68.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7515961_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:122840848(+)-23:122866812(-)__23_122843001_122868001D;SPAN=25964;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:24 DP:39 GQ:25.7 PL:[68.6, 0.0, 25.7] SR:0 DR:24 LR:-69.71 LO:69.71);ALT=A[chrX:122866812[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	123156522	+	chrX	123159690	+	.	0	7	7516652_1	12.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=7516652_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_123137001_123162001_37C;SPAN=3168;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:39 GQ:12.5 PL:[12.5, 0.0, 81.8] SR:7 DR:0 LR:-12.54 LO:15.5);ALT=G[chrX:123159690[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	123179218	+	chrX	123181202	+	.	3	3	7516684_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=7516684_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_123161501_123186501_153C;SPAN=1984;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:3 DR:3 LR:-1.062 LO:9.396);ALT=G[chrX:123181202[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	123480631	+	chrX	123499611	+	.	3	4	7517213_1	9.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GT;MAPQ=60;MATEID=7517213_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_123455501_123480501_8C;SPAN=18980;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:4 DP:0 GQ:0.9 PL:[9.9, 0.9, 0.0] SR:4 DR:3 LR:-9.903 LO:9.903);ALT=T[chrX:123499611[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	123480631	+	chrX	123504024	+	ATCACGGTTACATTTATACATACCGAGTGTCCCAGACAGAAACAGGTTCTTGGAGTGCTG	0	7	7517147_1	5.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=ATCACGGTTACATTTATACATACCGAGTGTCCCAGACAGAAACAGGTTCTTGGAGTGCTG;MAPQ=60;MATEID=7517147_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_123480001_123505001_6C;SPAN=23393;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:64 GQ:5.9 PL:[5.9, 0.0, 147.8] SR:7 DR:0 LR:-5.768 LO:13.86);ALT=T[chrX:123504024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	133507497	+	chrX	133511601	+	.	12	3	7530318_1	27.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7530318_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_133500501_133525501_119C;SPAN=4104;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:56 GQ:27.8 PL:[27.8, 0.0, 107.0] SR:3 DR:12 LR:-27.74 LO:30.42);ALT=G[chrX:133511601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	133594368	+	chrX	133607388	+	.	50	11	7530656_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=G;MAPQ=60;MATEID=7530656_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_133574001_133599001_157C;SPAN=13020;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:52 DP:30 GQ:13.8 PL:[151.8, 13.8, 0.0] SR:11 DR:50 LR:-151.8 LO:151.8);ALT=G[chrX:133607388[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	133594407	+	chrX	133609208	+	.	77	0	7530657_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7530657_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:133594407(+)-23:133609208(-)__23_133574001_133599001D;SPAN=14801;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:77 DP:17 GQ:20.7 PL:[227.7, 20.7, 0.0] SR:0 DR:77 LR:-227.8 LO:227.8);ALT=C[chrX:133609208[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135229817	+	chrX	135288563	+	.	29	0	7533858_1	86.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7533858_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:135229817(+)-23:135288563(-)__23_135264501_135289501D;SPAN=58746;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:36 GQ:0.2 PL:[86.0, 0.0, 0.2] SR:0 DR:29 LR:-91.0 LO:91.0);ALT=G[chrX:135288563[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135229898	+	chrX	135252064	+	.	12	0	7533703_1	33.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7533703_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:135229898(+)-23:135252064(-)__23_135240001_135265001D;SPAN=22166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:24 GQ:23.3 PL:[33.2, 0.0, 23.3] SR:0 DR:12 LR:-33.17 LO:33.17);ALT=G[chrX:135252064[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135326955	+	chrX	135328224	+	.	0	4	7534095_1	0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7534095_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_23_135313501_135338501_6C;SPAN=1269;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:50 GQ:0.3 PL:[0.0, 0.3, 122.1] SR:4 DR:0 LR:0.3422 LO:7.35);ALT=C[chrX:135328224[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135328501	+	chrX	135333448	+	.	14	7	7534097_1	45.0	.	DISC_MAPQ=53;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=7534097_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_135313501_135338501_280C;SPAN=4947;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:52 GQ:45.5 PL:[45.5, 0.0, 78.5] SR:7 DR:14 LR:-45.33 LO:45.88);ALT=C[chrX:135333448[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135579600	+	chrX	135581755	+	AGGAAACATGAGCGGCACCAACTTGGATGGGAACGATGAGTTTGATGAGCAGTTGCGAATGCAAGAATTGTACGGAGACGGCAAGGATGGTGACACCCAGACCGATGCCGGCGGAGAACCCGATTCTCTCGGGCAGCAGCCGACGGACACTCCCTACGAGTGGGACCTGGACAAAAAGGCTTGGTTCCCCA	0	11	7534268_1	22.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=AGGAAACATGAGCGGCACCAACTTGGATGGGAACGATGAGTTTGATGAGCAGTTGCGAATGCAAGAATTGTACGGAGACGGCAAGGATGGTGACACCCAGACCGATGCCGGCGGAGAACCCGATTCTCTCGGGCAGCAGCCGACGGACACTCCCTACGAGTGGGACCTGGACAAAAAGGCTTGGTTCCCCA;MAPQ=60;MATEID=7534268_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_135558501_135583501_197C;SPAN=2155;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:51 GQ:22.7 PL:[22.7, 0.0, 98.6] SR:11 DR:0 LR:-22.49 LO:25.34);ALT=T[chrX:135581755[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135829751	+	chrX	135862877	+	TTCCACTTGGAGGGTTGCACATCCTTTCAGGAAGTCATTGATGTTGTTGATGCAGTCAGCTTCAGTTTGGGGATCCAGACAAAA	0	24	7534758_1	72.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CT;INSERTION=TTCCACTTGGAGGGTTGCACATCCTTTCAGGAAGTCATTGATGTTGTTGATGCAGTCAGCTTCAGTTTGGGGATCCAGACAAAA;MAPQ=60;MATEID=7534758_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_135852501_135877501_167C;SPAN=33126;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:24 DP:25 GQ:6.6 PL:[72.6, 6.6, 0.0] SR:24 DR:0 LR:-72.62 LO:72.62);ALT=T[chrX:135862877[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	135861705	+	chrX	135862982	+	.	11	0	7534773_1	22.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7534773_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:135861705(+)-23:135862982(-)__23_135852501_135877501D;SPAN=1277;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:53 GQ:22.1 PL:[22.1, 0.0, 104.6] SR:0 DR:11 LR:-21.95 LO:25.13);ALT=A[chrX:135862982[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	148564752	+	chrX	148568455	+	.	3	2	7552162_1	9.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=7552162_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_148568001_148593001_281C;SPAN=3703;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:27 GQ:9.2 PL:[9.2, 0.0, 55.4] SR:2 DR:3 LR:-9.19 LO:11.14);ALT=G[chrX:148568455[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	148735758	+	chrX	148830979	-	.	41	0	7552645_1	99.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7552645_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:148735758(+)-23:148830979(+)__23_148813001_148838001D;SPAN=95221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:24 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:0 DR:41 LR:-118.8 LO:118.8);ALT=T]chrX:148830979];VARTYPE=BND:INV-hh;JOINTYPE=hh
chrX	149983411	+	chrX	149984477	+	.	0	8	7554165_1	12.0	.	EVDNC=ASSMB;HOMSEQ=TACCT;MAPQ=60;MATEID=7554165_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_149964501_149989501_228C;SPAN=1066;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:51 GQ:12.8 PL:[12.8, 0.0, 108.5] SR:8 DR:0 LR:-12.59 LO:17.19);ALT=T[chrX:149984477[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	149999797	+	chrX	150067020	+	.	9	0	7554329_1	26.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7554329_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:149999797(+)-23:150067020(-)__23_150062501_150087501D;SPAN=67223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:13 GQ:3.2 PL:[26.3, 0.0, 3.2] SR:0 DR:9 LR:-26.96 LO:26.96);ALT=T[chrX:150067020[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	150244965	-	chrX	150246916	+	TGAGGAGCCCTGACTGCACCTAGACAGGCATGGATCTCAAC	4	7	7554729_1	3.0	.	DISC_MAPQ=55;EVDNC=TSI_L;HOMSEQ=AAGTGCT;INSERTION=TGAGGAGCCCTGACTGCACCTAGACAGGCATGGATCTCAAC;MAPQ=15;MATEID=7554729_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_150234001_150259001_89C;SPAN=1951;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:73 GQ:3.5 PL:[3.5, 0.0, 171.8] SR:7 DR:4 LR:-3.33 LO:13.44);ALT=[chrX:150246916[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chrX	150293942	+	chrX	150295716	+	.	39	34	7554681_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=GAA;MAPQ=60;MATEID=7554681_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_150283001_150308001_38C;SPAN=1774;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:59 DP:15 GQ:15.9 PL:[174.9, 15.9, 0.0] SR:34 DR:39 LR:-174.9 LO:174.9);ALT=A[chrX:150295716[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	150565794	+	chrX	150573385	+	.	15	0	7555027_1	36.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7555027_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:150565794(+)-23:150573385(-)__23_150552501_150577501D;SPAN=7591;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:49 GQ:36.2 PL:[36.2, 0.0, 82.4] SR:0 DR:15 LR:-36.24 LO:37.24);ALT=A[chrX:150573385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	150565833	+	chrX	150572100	+	.	35	19	7555028_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CAG;MAPQ=60;MATEID=7555028_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_150552501_150577501_214C;SPAN=6267;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:46 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:19 DR:35 LR:-148.5 LO:148.5);ALT=G[chrX:150572100[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	150572213	+	chrX	150573386	+	.	0	40	7555037_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7555037_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_150552501_150577501_251C;SPAN=1173;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:69 GQ:53.9 PL:[113.3, 0.0, 53.9] SR:40 DR:0 LR:-114.5 LO:114.5);ALT=G[chrX:150573386[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
