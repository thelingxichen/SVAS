chr6	6163630	+	chr6	6164671	-	.	9	0	4002299_1	0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4002299_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6163630(+)-6:6164671(+)__6_6149501_6174501D;SPAN=1041;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:143 GQ:8.7 PL:[0.0, 8.7, 363.0] SR:0 DR:9 LR:9.033 LO:15.57);ALT=T]chr6:6164671];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	6312664	+	chr6	9434113	-	.	36	141	4004107_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=ACTTTGG;MAPQ=60;MATEID=4004107_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_6_6296501_6321501_491C;SPAN=3121449;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:153 DP:39 GQ:41.2 PL:[452.2, 41.2, 0.0] SR:141 DR:36 LR:-452.2 LO:452.2);ALT=G]chr6:9434113];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	6312782	-	chr6	9434001	+	.	33	0	4004109_1	95.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=32;MATEID=4004109_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=6:6312782(-)-6:9434001(-)__6_6296501_6321501D;SPAN=3121219;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:33 DP:10 GQ:8.7 PL:[95.7, 8.7, 0.0] SR:0 DR:33 LR:-95.72 LO:95.72);ALT=[chr6:9434001[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr6	48952287	+	chr6	7442113	+	.	18	86	4009120_1	99.0	.	DISC_MAPQ=32;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4009120_2;MATENM=1;NM=7;NUMPARTS=2;SCTG=c_6_7423501_7448501_9C;SPAN=41510174;SUBN=4;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:91 DP:35 GQ:24.3 PL:[267.3, 24.3, 0.0] SR:86 DR:18 LR:-267.4 LO:267.4);ALT=]chr6:48952287]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr11	64154407	+	chr6	8439300	+	.	0	29	4012921_1	85.0	.	EVDNC=ASSMB;HOMSEQ=CCTTCCTTCCTTCCTTTCTT;MAPQ=60;MATEID=4012921_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_6_8428001_8453001_14C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:29 DP:17 GQ:7.8 PL:[85.8, 7.8, 0.0] SR:29 DR:0 LR:-85.82 LO:85.82);ALT=]chr11:64154407]C;VARTYPE=BND:TRX-th;JOINTYPE=th
chr11	63446610	+	chr11	63447746	-	.	8	0	6849764_1	0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=6849764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63446610(+)-11:63447746(+)__11_63430501_63455501D;SPAN=1136;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:133 GQ:9.3 PL:[0.0, 9.3, 339.9] SR:0 DR:8 LR:9.625 LO:13.68);ALT=A]chr11:63447746];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	63561696	+	chr11	63563025	-	.	8	0	6850927_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=6850927_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:63561696(+)-11:63563025(+)__11_63553001_63578001D;SPAN=1329;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:147 GQ:13.3 PL:[0.0, 13.3, 382.8] SR:0 DR:8 LR:13.42 LO:13.32);ALT=T]chr11:63563025];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr11	64047134	-	chr11	64048200	+	.	15	0	6852995_1	14.0	.	DISC_MAPQ=40;EVDNC=DSCRD;IMPRECISE;MAPQ=40;MATEID=6852995_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=11:64047134(-)-11:64048200(-)__11_64043001_64068001D;SPAN=1066;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:15 DP:128 GQ:14.9 PL:[14.9, 0.0, 295.4] SR:0 DR:15 LR:-14.84 LO:30.18);ALT=[chr11:64048200[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
