chr16	81010072	+	chr16	81015411	+	TGTA	3	3	6260514_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TGTA;MAPQ=60;MATEID=6260514_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_80997001_81022001_61C;SPAN=5339;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:69 GQ:1.1 PL:[1.1, 0.0, 166.1] SR:3 DR:3 LR:-1.112 LO:11.25);ALT=A[chr16:81015411[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	81015482	+	chr16	81030919	+	.	0	19	6260524_1	54.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6260524_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_80997001_81022001_240C;SPAN=15437;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:30 GQ:18.2 PL:[54.5, 0.0, 18.2] SR:19 DR:0 LR:-55.59 LO:55.59);ALT=G[chr16:81030919[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	81015531	+	chr16	81040392	+	.	9	0	6260525_1	23.0	.	DISC_MAPQ=55;EVDNC=DSCRD;IMPRECISE;MAPQ=55;MATEID=6260525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=16:81015531(+)-16:81040392(-)__16_80997001_81022001D;SPAN=24861;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:24 GQ:23.3 PL:[23.3, 0.0, 33.2] SR:0 DR:9 LR:-23.21 LO:23.34);ALT=G[chr16:81040392[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	81031035	+	chr16	81040337	+	.	42	22	6260430_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=60;MATEID=6260430_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_16_81021501_81046501_277C;SPAN=9302;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:72 GQ:26.9 PL:[145.7, 0.0, 26.9] SR:22 DR:42 LR:-149.9 LO:149.9);ALT=C[chr16:81040337[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr16	81053882	+	chr16	81056357	+	.	0	13	6260321_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=6260321_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_16_81046001_81071001_68C;SPAN=2475;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:47 GQ:30.2 PL:[30.2, 0.0, 83.0] SR:13 DR:0 LR:-30.18 LO:31.58);ALT=G[chr16:81056357[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
