chr7	85853700	+	chr7	85844668	+	GTC	22	19	3434852_1	98.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=GTC;MAPQ=60;MATEID=3434852_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_7_85848001_85873001_144C;SPAN=9032;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:34 DP:51 GQ:22.7 PL:[98.6, 0.0, 22.7] SR:19 DR:22 LR:-100.8 LO:100.8);ALT=]chr7:85853700]A;VARTYPE=BND:DUP-th;JOINTYPE=th
