chr3	133377996	+	chr3	133379888	+	.	0	8	1664217_1	4.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=1664217_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_133378001_133403001_16C;SPAN=1892;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:82 GQ:4.4 PL:[4.4, 0.0, 192.5] SR:8 DR:0 LR:-4.192 LO:15.42);ALT=T[chr3:133379888[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	133503782	+	chr3	133505083	+	.	45	32	1664430_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AACAATACTATTTTTT;MAPQ=60;MATEID=1664430_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_133500501_133525501_38C;SPAN=1301;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:62 DP:62 GQ:16.5 PL:[181.5, 16.5, 0.0] SR:32 DR:45 LR:-181.5 LO:181.5);ALT=T[chr3:133505083[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	133534570	+	chr3	133535720	+	.	0	5	1664624_1	0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=1664624_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_133525001_133550001_102C;SPAN=1150;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:91 GQ:7.8 PL:[0.0, 7.8, 234.3] SR:5 DR:0 LR:8.149 LO:8.345);ALT=G[chr3:133535720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	134197558	+	chr3	134201648	+	.	0	18	1667354_1	29.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=1667354_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_134186501_134211501_251C;SPAN=4090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:111 GQ:29.6 PL:[29.6, 0.0, 237.5] SR:18 DR:0 LR:-29.35 LO:38.97);ALT=C[chr3:134201648[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	134197606	+	chr3	134204793	+	.	22	0	1667355_1	43.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=1667355_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:134197606(+)-3:134204793(-)__3_134186501_134211501D;SPAN=7187;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:107 GQ:43.7 PL:[43.7, 0.0, 215.3] SR:0 DR:22 LR:-43.63 LO:50.16);ALT=C[chr3:134204793[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
