chr1	211500263	+	chr1	211526580	+	.	11	0	528432_1	21.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=528432_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:211500263(+)-1:211526580(-)__1_211508501_211533501D;SPAN=26317;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:56 GQ:21.2 PL:[21.2, 0.0, 113.6] SR:0 DR:11 LR:-21.14 LO:24.83);ALT=C[chr1:211526580[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	211556267	+	chr1	211564958	+	.	7	7	528833_1	19.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=528833_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_211557501_211582501_184C;SPAN=8691;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:51 GQ:19.4 PL:[19.4, 0.0, 101.9] SR:7 DR:7 LR:-19.19 LO:22.57);ALT=A[chr1:211564958[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212471153	+	chr1	212472617	+	.	99	52	532013_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AAGATGAAGTGAATTGTT;MAPQ=60;MATEID=532013_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212464001_212489001_39C;SPAN=1464;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:121 DP:40 GQ:32.4 PL:[356.4, 32.4, 0.0] SR:52 DR:99 LR:-356.5 LO:356.5);ALT=T[chr1:212472617[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212583910	+	chr1	212588140	+	.	8	0	532608_1	11.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=532608_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:212583910(+)-1:212588140(-)__1_212562001_212587001D;SPAN=4230;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:0 DR:8 LR:-11.51 LO:16.91);ALT=C[chr1:212588140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212606388	+	chr1	212615903	+	.	40	0	532695_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=532695_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:212606388(+)-1:212615903(-)__1_212611001_212636001D;SPAN=9515;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:40 DP:62 GQ:32.9 PL:[115.4, 0.0, 32.9] SR:0 DR:40 LR:-117.6 LO:117.6);ALT=C[chr1:212615903[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212606462	+	chr1	212617679	+	.	24	4	532696_1	67.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=532696_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212611001_212636001_34C;SPAN=11217;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:57 GQ:67.1 PL:[67.1, 0.0, 70.4] SR:4 DR:24 LR:-67.08 LO:67.09);ALT=G[chr1:212617679[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212617784	+	chr1	212619172	+	.	0	30	532742_1	67.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=532742_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212611001_212636001_266C;SPAN=1388;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:116 GQ:67.7 PL:[67.7, 0.0, 212.9] SR:30 DR:0 LR:-67.6 LO:71.85);ALT=T[chr1:212619172[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212782272	+	chr1	212788358	+	.	46	50	533281_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=533281_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212758001_212783001_218C;SPAN=6086;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:78 DP:90 GQ:14.4 PL:[247.5, 14.4, 0.0] SR:50 DR:46 LR:-251.9 LO:251.9);ALT=G[chr1:212788358[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212788605	+	chr1	212791467	+	.	8	12	533401_1	32.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGT;MAPQ=60;MATEID=533401_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_212782501_212807501_191C;SPAN=2862;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:101 GQ:32.3 PL:[32.3, 0.0, 210.5] SR:12 DR:8 LR:-32.05 LO:39.78);ALT=T[chr1:212791467[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212957836	+	chr1	212964872	+	CATAAAACAATTATCTGAAGCTTCCTGCCATGCTTGCCCATTAATGCTGATATTCTCTTGCACAGCTGATTCAAAAGT	0	15	533846_1	21.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=CATAAAACAATTATCTGAAGCTTCCTGCCATGCTTGCCCATTAATGCTGATATTCTCTTGCACAGCTGATTCAAAAGT;MAPQ=60;MATEID=533846_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_1_212954001_212979001_296C;SPAN=7036;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:104 GQ:21.5 PL:[21.5, 0.0, 229.4] SR:15 DR:0 LR:-21.34 LO:31.64);ALT=C[chr1:212964872[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	212983252	-	chr1	212985112	+	.	8	0	534028_1	0	.	DISC_MAPQ=38;EVDNC=DSCRD;IMPRECISE;MAPQ=38;MATEID=534028_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:212983252(-)-1:212985112(-)__1_212978501_213003501D;SPAN=1860;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:8 DP:108 GQ:2.7 PL:[0.0, 2.7, 267.3] SR:0 DR:8 LR:2.852 LO:14.42);ALT=[chr1:212985112[G;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr1	213224767	+	chr1	213251034	+	.	8	0	535129_1	7.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=535129_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:213224767(+)-1:213251034(-)__1_213223501_213248501D;SPAN=26267;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:0 DR:8 LR:-7.443 LO:16.0);ALT=G[chr1:213251034[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
