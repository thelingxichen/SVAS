chr13	89110977	-	chr13	89112603	+	ATATTATATTATAATATAA	18	44	8206899_1	99.0	.	DISC_MAPQ=10;EVDNC=ASDIS;INSERTION=ATATTATATTATAATATAA;MAPQ=60;MATEID=8206899_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_13_89106501_89131501_192C;SPAN=1626;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:52 DP:87 GQ:62.3 PL:[148.1, 0.0, 62.3] SR:44 DR:18 LR:-149.9 LO:149.9);ALT=[chr13:89112603[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr13	89645968	+	chr13	89650857	+	.	15	11	8209043_1	47.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=8209043_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_89621001_89646001_12C;SPAN=4889;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:20 DP:71 GQ:47 PL:[47.0, 0.0, 122.9] SR:11 DR:15 LR:-46.78 LO:48.78);ALT=T[chr13:89650857[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
