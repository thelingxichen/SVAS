chr1	100598833	+	chr1	100602435	+	.	8	0	250525_1	13.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=250525_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=1:100598833(+)-1:100602435(-)__1_100597001_100622001D;SPAN=3602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:49 GQ:13.1 PL:[13.1, 0.0, 105.5] SR:0 DR:8 LR:-13.13 LO:17.35);ALT=G[chr1:100602435[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr1	100732181	+	chr1	100733706	+	.	0	8	250970_1	7.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=250970_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_1_100719501_100744501_115C;SPAN=1525;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:70 GQ:7.4 PL:[7.4, 0.0, 162.5] SR:8 DR:0 LR:-7.443 LO:16.0);ALT=G[chr1:100733706[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
