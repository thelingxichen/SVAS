chr15	74800751	-	chr15	74802028	+	.	8	0	8983731_1	0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=8983731_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=15:74800751(-)-15:74802028(-)__15_74798501_74823501D;SPAN=1277;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:177 GQ:21.4 PL:[0.0, 21.4, 472.0] SR:0 DR:8 LR:21.55 LO:12.66);ALT=[chr15:74802028[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr15	75170356	-	chr15	75171566	+	.	8	4	8986122_1	3.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=ATTTTTTGTATTTTTAGTA;MAPQ=60;MATEID=8986122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_15_75166001_75191001_176C;SPAN=1210;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:121 GQ:3.8 PL:[3.8, 0.0, 287.6] SR:4 DR:8 LR:-3.529 LO:20.85);ALT=[chr15:75171566[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
