chr5	118604602	+	chr5	118728511	+	.	15	6	2564631_1	47.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2564631_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_118727001_118752001_280C;SPAN=123909;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:32 GQ:27.8 PL:[47.6, 0.0, 27.8] SR:6 DR:15 LR:-47.65 LO:47.65);ALT=A[chr5:118728511[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	118788306	+	chr5	118809601	+	.	14	0	2564711_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=2564711_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:118788306(+)-5:118809601(-)__5_118800501_118825501D;SPAN=21295;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:29 GQ:31.7 PL:[38.3, 0.0, 31.7] SR:0 DR:14 LR:-38.39 LO:38.39);ALT=A[chr5:118809601[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	118788329	+	chr5	118792008	+	.	6	5	2564799_1	6.0	.	DISC_MAPQ=59;EVDNC=TSI_L;HOMSEQ=AGG;MAPQ=60;MATEID=2564799_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_5_118776001_118801001_218C;SPAN=3679;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:48 GQ:6.8 PL:[6.8, 0.0, 109.1] SR:5 DR:6 LR:-6.802 LO:12.25);ALT=G[chr5:118792008[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	118814716	+	chr5	118824885	+	.	3	2	2564733_1	0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2564733_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_118800501_118825501_151C;SPAN=10169;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:61 GQ:0.2 PL:[0.2, 0.0, 145.4] SR:2 DR:3 LR:0.0214 LO:9.242);ALT=G[chr5:118824885[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	118861719	+	chr5	118862825	+	.	2	4	2564773_1	2.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGG;MAPQ=60;MATEID=2564773_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_118849501_118874501_193C;SPAN=1106;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:51 GQ:2.9 PL:[2.9, 0.0, 118.4] SR:4 DR:2 LR:-2.688 LO:9.65);ALT=G[chr5:118862825[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
