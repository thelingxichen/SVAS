chr5	153414575	+	chr5	153418413	+	.	8	0	2617054_1	12.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2617054_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:153414575(+)-5:153418413(-)__5_153394501_153419501D;SPAN=3838;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:0 DR:8 LR:-12.05 LO:17.05);ALT=T[chr5:153418413[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	154320741	+	chr5	154330379	+	.	14	0	2618763_1	40.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2618763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:154320741(+)-5:154330379(-)__5_154301001_154326001D;SPAN=9638;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:20 GQ:7.7 PL:[40.7, 0.0, 7.7] SR:0 DR:14 LR:-42.07 LO:42.07);ALT=T[chr5:154330379[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	154320745	+	chr5	154335929	+	.	13	0	2618764_1	37.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2618764_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:154320745(+)-5:154335929(-)__5_154301001_154326001D;SPAN=15184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:21 GQ:11 PL:[37.4, 0.0, 11.0] SR:0 DR:13 LR:-37.82 LO:37.82);ALT=A[chr5:154335929[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	154320859	+	chr5	154336693	+	.	8	0	2618766_1	20.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=2618766_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=5:154320859(+)-5:154336693(-)__5_154301001_154326001D;SPAN=15834;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:24 GQ:20 PL:[20.0, 0.0, 36.5] SR:0 DR:8 LR:-19.91 LO:20.23);ALT=C[chr5:154336693[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	154339609	+	chr5	154346243	+	.	0	8	2618717_1	11.0	.	EVDNC=ASSMB;HOMSEQ=TAG;MAPQ=60;MATEID=2618717_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_154325501_154350501_160C;SPAN=6634;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:55 GQ:11.6 PL:[11.6, 0.0, 120.5] SR:8 DR:0 LR:-11.51 LO:16.91);ALT=G[chr5:154346243[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	62029870	+	chr5	155039561	+	TGGGGAATTGGTTCCATATGAACTTTAAAG	18	84	2872260_1	99.0	.	DISC_MAPQ=0;EVDNC=ASDIS;INSERTION=TGGGGAATTGGTTCCATATGAACTTTAAAG;MAPQ=60;MATEID=2872260_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_6_62009501_62034501_169C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:25 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:84 DR:18 LR:-254.2 LO:254.2);ALT=]chr6:62029870]T;VARTYPE=BND:TRX-th;JOINTYPE=th
chr5	155656242	-	chrX	119488901	+	.	3	11	7511753_1	29.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=ATACATACATATATATATATA;MAPQ=42;MATEID=7511753_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_23_119486501_119511501_20C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:11 DP:7 GQ:2.7 PL:[29.7, 2.7, 0.0] SR:11 DR:3 LR:-29.71 LO:29.71);ALT=[chrX:119488901[A;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr6	62200437	+	chr6	62206527	+	.	45	22	2873056_1	99.0	.	DISC_MAPQ=57;EVDNC=ASDIS;HOMSEQ=AGATGAATGCACACATCACAAAG;MAPQ=60;MATEID=2873056_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_62205501_62230501_262C;SPAN=6090;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:63 DP:30 GQ:16.8 PL:[184.8, 16.8, 0.0] SR:22 DR:45 LR:-184.8 LO:184.8);ALT=G[chr6:62206527[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	117861699	+	chrX	117874978	+	.	9	0	7508763_1	24.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7508763_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:117861699(+)-23:117874978(-)__23_117845001_117870001D;SPAN=13279;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:19 GQ:21.2 PL:[24.5, 0.0, 21.2] SR:0 DR:9 LR:-24.57 LO:24.57);ALT=A[chrX:117874978[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118602603	+	chrX	118603621	+	.	98	0	7510061_1	99.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7510061_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:118602603(+)-23:118603621(-)__23_118580001_118605001D;SPAN=1018;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:98 DP:96 GQ:26.4 PL:[290.4, 26.4, 0.0] SR:0 DR:98 LR:-290.5 LO:290.5);ALT=T[chrX:118603621[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118708664	+	chrX	118715468	+	.	10	0	7510120_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7510120_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:118708664(+)-23:118715468(-)__23_118702501_118727501D;SPAN=6804;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:65 GQ:15.5 PL:[15.5, 0.0, 140.9] SR:0 DR:10 LR:-15.4 LO:21.4);ALT=C[chrX:118715468[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118708945	+	chrX	118715469	+	CCTGAAGGGACCCCGTTTGAGGAT	0	29	7510122_1	78.0	.	EVDNC=ASSMB;INSERTION=CCTGAAGGGACCCCGTTTGAGGAT;MAPQ=60;MATEID=7510122_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118702501_118727501_66C;SPAN=6524;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:65 GQ:78.2 PL:[78.2, 0.0, 78.2] SR:29 DR:0 LR:-78.12 LO:78.12);ALT=G[chrX:118715469[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118715559	+	chrX	118717088	+	TCTATGCAGATGGTAGTATATGTCTGGACATACTTCAGAACCGTTGGAGTCCAACCTATGATGTGTCTTCCATTCTAACATCCATAC	0	15	7510129_1	35.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=AG;INSERTION=TCTATGCAGATGGTAGTATATGTCTGGACATACTTCAGAACCGTTGGAGTCCAACCTATGATGTGTCTTCCATTCTAACATCCATAC;MAPQ=60;MATEID=7510129_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118702501_118727501_32C;SPAN=1529;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:54 GQ:35 PL:[35.0, 0.0, 94.4] SR:15 DR:0 LR:-34.89 LO:36.48);ALT=G[chrX:118717088[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118754015	+	chrX	118759298	+	.	10	8	7510492_1	43.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7510492_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GG;SCTG=c_23_118751501_118776501_145C;SPAN=5283;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:8 DR:10 LR:-43.7 LO:44.82);ALT=C[chrX:118759298[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118754015	+	chrX	118763281	+	AGGACCCTGGGTCTCATGCAGCATGCAGCAAACAGCAGAGTTAA	19	10	7510493_1	60.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AGGACCCTGGGTCTCATGCAGCATGCAGCAAACAGCAGAGTTAA;MAPQ=60;MATEID=7510493_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118751501_118776501_145C;SPAN=9266;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:58 GQ:60.2 PL:[60.2, 0.0, 80.0] SR:10 DR:19 LR:-60.21 LO:60.37);ALT=C[chrX:118763281[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118763473	+	chrX	118767323	+	.	8	11	7510520_1	44.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7510520_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118751501_118776501_306C;SPAN=3850;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:66 GQ:44.9 PL:[44.9, 0.0, 114.2] SR:11 DR:8 LR:-44.84 LO:46.56);ALT=T[chrX:118767323[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118767458	+	chrX	118770990	+	.	10	11	7510527_1	44.0	.	DISC_MAPQ=50;EVDNC=TSI_L;HOMSEQ=CTG;MAPQ=60;MATEID=7510527_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118751501_118776501_318C;SPAN=3532;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:55 GQ:44.6 PL:[44.6, 0.0, 87.5] SR:11 DR:10 LR:-44.52 LO:45.33);ALT=G[chrX:118770990[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118767458	+	chrX	118774655	+	AAGGGTTTGCTGTCAGGGTCGGTGTCCTTGAAGCCCATCTCCTCCAGCTTACAGCGGCGATACAGCTCATAGTGCCGGGTGTGGGTCTGCTCCCGCAGATCCTCCATGTTGACCCGAATCAGCATCTCCCGCAGCTTCACAAAGTCGCAGTGGGCCTCGTTTTCAA	3	43	7510528_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=AAGGGTTTGCTGTCAGGGTCGGTGTCCTTGAAGCCCATCTCCTCCAGCTTACAGCGGCGATACAGCTCATAGTGCCGGGTGTGGGTCTGCTCCCGCAGATCCTCCATGTTGACCCGAATCAGCATCTCCCGCAGCTTCACAAAGTCGCAGTGGGCCTCGTTTTCAA;MAPQ=60;MATEID=7510528_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118751501_118776501_318C;SPAN=7197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:45 DP:69 GQ:37.4 PL:[129.8, 0.0, 37.4] SR:43 DR:3 LR:-132.7 LO:132.7);ALT=G[chrX:118774655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118771159	+	chrX	118774655	+	.	6	38	7510538_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7510538_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118751501_118776501_318C;SPAN=3496;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:44 DP:79 GQ:67.7 PL:[123.8, 0.0, 67.7] SR:38 DR:6 LR:-124.7 LO:124.7);ALT=C[chrX:118774655[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118774751	+	chrX	118783899	+	.	0	14	7510544_1	38.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=7510544_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118751501_118776501_212C;SPAN=9148;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:30 GQ:34.7 PL:[38.0, 0.0, 34.7] SR:14 DR:0 LR:-38.09 LO:38.09);ALT=C[chrX:118783899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118787005	+	chrX	118797445	+	.	5	9	7510341_1	31.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=7510341_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118776001_118801001_150C;SPAN=10440;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:42 GQ:31.7 PL:[31.7, 0.0, 68.0] SR:9 DR:5 LR:-31.53 LO:32.35);ALT=T[chrX:118797445[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118797641	+	chrX	118809516	+	.	0	88	7510432_1	99.0	.	EVDNC=ASSMB;HOMSEQ=CC;MAPQ=60;MATEID=7510432_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118800501_118825501_248C;SPAN=11875;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:88 DP:58 GQ:23.7 PL:[260.7, 23.7, 0.0] SR:88 DR:0 LR:-260.8 LO:260.8);ALT=C[chrX:118809516[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118797689	+	chrX	118827042	+	.	65	0	7510364_1	99.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7510364_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:118797689(+)-23:118827042(-)__23_118825001_118850001D;SPAN=29353;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:65 DP:36 GQ:17.4 PL:[191.4, 17.4, 0.0] SR:0 DR:65 LR:-191.4 LO:191.4);ALT=A[chrX:118827042[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118809632	+	chrX	118827038	+	.	82	19	7510456_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=7510456_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118800501_118825501_238C;SPAN=17406;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:92 DP:27 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:19 DR:82 LR:-270.7 LO:270.7);ALT=C[chrX:118827038[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118969040	+	chrX	118971718	+	.	15	0	7510899_1	38.0	.	DISC_MAPQ=59;EVDNC=DSCRD;IMPRECISE;MAPQ=59;MATEID=7510899_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:118969040(+)-23:118971718(-)__23_118947501_118972501D;SPAN=2678;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:43 GQ:38 PL:[38.0, 0.0, 64.4] SR:0 DR:15 LR:-37.87 LO:38.3);ALT=T[chrX:118971718[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	118985566	+	chrX	118986733	+	CGTATCATTAGAAAAAAACTCAAAATAATCATGCTCAGGCATAGGTTGAAGATGTTCCTGAAGCTGCTCCTTGGTCAAAGTGGGAGGTAATCTTCGAATTAC	0	28	7510829_1	74.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CACCTT;INSERTION=CGTATCATTAGAAAAAAACTCAAAATAATCATGCTCAGGCATAGGTTGAAGATGTTCCTGAAGCTGCTCCTTGGTCAAAGTGGGAGGTAATCTTCGAATTAC;MAPQ=60;MATEID=7510829_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_118972001_118997001_194C;SPAN=1167;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:68 GQ:74 PL:[74.0, 0.0, 90.5] SR:28 DR:0 LR:-74.01 LO:74.1);ALT=T[chrX:118986733[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119005977	+	chrX	119007268	+	A	0	109	7511141_1	99.0	.	EVDNC=ASSMB;INSERTION=A;MAPQ=60;MATEID=7511141_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118996501_119021501_121C;SPAN=1291;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:109 DP:142 GQ:21.2 PL:[321.5, 0.0, 21.2] SR:109 DR:0 LR:-336.6 LO:336.6);ALT=G[chrX:119007268[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119005991	+	chrX	119010473	+	.	22	0	7511142_1	48.0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=7511142_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:119005991(+)-23:119010473(-)__23_118996501_119021501D;SPAN=4482;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:88 GQ:48.8 PL:[48.8, 0.0, 164.3] SR:0 DR:22 LR:-48.78 LO:52.31);ALT=G[chrX:119010473[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119007357	+	chrX	119010475	+	.	0	130	7511145_1	99.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=7511145_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_118996501_119021501_52C;SPAN=3118;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:130 DP:160 GQ:2.8 PL:[385.7, 0.0, 2.8] SR:130 DR:0 LR:-409.2 LO:409.2);ALT=G[chrX:119010475[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119070396	+	chrX	119077182	+	TCTGAAGTAGAAGCTGAAGTAGTGCTTTTCTTTGGCTCTTCATCCTCCACTGGTGTATGTTCATCAGAATCTGGTTCAGGATTCTTTGGAGAAAGTCCCCATACTTCAGGAGCTCCCAATTCTCCAATTCTCTCTCTCTCACTTAATCT	0	20	7511060_1	50.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=C;INSERTION=TCTGAAGTAGAAGCTGAAGTAGTGCTTTTCTTTGGCTCTTCATCCTCCACTGGTGTATGTTCATCAGAATCTGGTTCAGGATTCTTTGGAGAAAGTCCCCATACTTCAGGAGCTCCCAATTCTCCAATTCTCTCTCTCTCACTTAATCT;MAPQ=60;MATEID=7511060_2;MATENM=0;NM=0;NUMPARTS=4;SCTG=c_23_119070001_119095001_197C;SPAN=6786;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:58 GQ:50.3 PL:[50.3, 0.0, 89.9] SR:20 DR:0 LR:-50.31 LO:50.93);ALT=T[chrX:119077182[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119575750	+	chrX	119580160	+	GGAGCCATTAACCAAATACATGCTGATGTTCACTTCCTTCAGATAAAATCGGTTTTCATTTTT	6	8	7511905_1	23.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=C;INSERTION=GGAGCCATTAACCAAATACATGCTGATGTTCACTTCCTTCAGATAAAATCGGTTTTCATTTTT;MAPQ=60;MATEID=7511905_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_119560001_119585001_142C;SPAN=4410;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:58 GQ:23.9 PL:[23.9, 0.0, 116.3] SR:8 DR:6 LR:-23.9 LO:27.4);ALT=C[chrX:119580160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119576518	+	chrX	119580160	+	.	2	4	7511908_1	3.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=C;MAPQ=60;MATEID=7511908_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_119560001_119585001_142C;SPAN=3642;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:49 GQ:3.2 PL:[3.2, 0.0, 115.4] SR:4 DR:2 LR:-3.23 LO:9.742);ALT=C[chrX:119580160[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119580285	+	chrX	119581694	+	.	3	5	7511914_1	6.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCTT;MAPQ=60;MATEID=7511914_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_119560001_119585001_165C;SPAN=1409;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:60 GQ:6.8 PL:[6.8, 0.0, 138.8] SR:5 DR:3 LR:-6.852 LO:14.07);ALT=T[chrX:119581694[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119589425	+	chrX	119602960	+	ATAAGTTTTATTTGTAGTTTCATAGCGAACTGTGAAATTCATCTGCCATTTTGCATAAAGGCAAGTGGCATTTTCTGAATCTGTCAAATTAAGTTCCAATGCATAAGACCGCACAGCT	0	31	7511928_1	83.0	.	DISC_MAPQ=255;EVDNC=TSI_G;HOMSEQ=CC;INSERTION=ATAAGTTTTATTTGTAGTTTCATAGCGAACTGTGAAATTCATCTGCCATTTTGCATAAAGGCAAGTGGCATTTTCTGAATCTGTCAAATTAAGTTCCAATGCATAAGACCGCACAGCT;MAPQ=60;MATEID=7511928_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_23_119584501_119609501_84C;SPAN=13535;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:31 DP:71 GQ:83.3 PL:[83.3, 0.0, 86.6] SR:31 DR:0 LR:-83.1 LO:83.11);ALT=T[chrX:119602960[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119589425	+	chrX	119590506	+	.	4	7	7511927_1	18.0	.	DISC_MAPQ=60;EVDNC=TSI_L;MAPQ=60;MATEID=7511927_2;MATENM=1;NM=0;NUMPARTS=3;REPSEQ=TTTT;SCTG=c_23_119584501_119609501_84C;SPAN=1081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:41 GQ:18.8 PL:[18.8, 0.0, 78.2] SR:7 DR:4 LR:-18.6 LO:20.81);ALT=T[chrX:119590506[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119590674	+	chrX	119603061	+	.	18	0	7511935_1	43.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=7511935_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:119590674(+)-23:119603061(-)__23_119584501_119609501D;SPAN=12387;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:58 GQ:43.7 PL:[43.7, 0.0, 96.5] SR:0 DR:18 LR:-43.7 LO:44.82);ALT=T[chrX:119603061[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chrX	119738149	+	chrX	119739932	+	.	13	0	7512365_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=7512365_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=23:119738149(+)-23:119739932(-)__23_119731501_119756501D;SPAN=1783;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:58 GQ:27.2 PL:[27.2, 0.0, 113.0] SR:0 DR:13 LR:-27.2 LO:30.19);ALT=G[chrX:119739932[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
