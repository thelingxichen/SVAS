chr6	143610134	+	chr6	143611280	-	.	2	4	3056409_1	0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=TCTT;MAPQ=60;MATEID=3056409_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_143594501_143619501_190C;SPAN=1146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:66 GQ:4.5 PL:[0.0, 4.5, 168.3] SR:4 DR:2 LR:4.677 LO:6.851);ALT=A]chr6:143611280];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr6	144471841	+	chr6	144507757	+	.	0	12	3058662_1	30.0	.	EVDNC=ASSMB;HOMSEQ=CAGG;MAPQ=60;MATEID=3058662_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_144501001_144526001_174C;SPAN=35916;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:34 GQ:30.5 PL:[30.5, 0.0, 50.3] SR:12 DR:0 LR:-30.4 LO:30.71);ALT=G[chr6:144507757[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr6	144606960	+	chr6	144612871	+	.	5	4	3058916_1	5.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AGGTA;MAPQ=60;MATEID=3058916_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_6_144599001_144624001_226C;SPAN=5911;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:65 GQ:5.6 PL:[5.6, 0.0, 150.8] SR:4 DR:5 LR:-5.497 LO:13.81);ALT=A[chr6:144612871[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
