chr10	134533815	+	chr10	134532717	+	.	9	0	4725156_1	16.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=4725156_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134532717(-)-10:134533815(+)__10_134529501_134554501D;SPAN=1098;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:49 GQ:16.4 PL:[16.4, 0.0, 102.2] SR:0 DR:9 LR:-16.43 LO:20.02);ALT=]chr10:134533815]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	134825456	+	chr10	134824111	+	.	71	0	4725568_1	99.0	.	DISC_MAPQ=30;EVDNC=DSCRD;IMPRECISE;MAPQ=30;MATEID=4725568_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:134824111(-)-10:134825456(+)__10_134823501_134848501D;SPAN=1345;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:71 DP:68 GQ:18.9 PL:[207.9, 18.9, 0.0] SR:0 DR:71 LR:-208.0 LO:208.0);ALT=]chr10:134825456]G;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	135089092	+	chr10	135090276	+	.	4	2	4726082_1	4.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4726082_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_135068501_135093501_40C;SPAN=1184;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:32 GQ:4.7 PL:[4.7, 0.0, 70.7] SR:2 DR:4 LR:-4.534 LO:8.169);ALT=C[chr10:135090276[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135093408	+	chr10	135094776	+	.	0	5	4725991_1	2.0	.	EVDNC=ASSMB;HOMSEQ=CCTG;MAPQ=60;MATEID=4725991_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_135093001_135118001_71C;SPAN=1368;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:53 GQ:2.3 PL:[2.3, 0.0, 124.4] SR:5 DR:0 LR:-2.146 LO:9.562);ALT=G[chr10:135094776[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135103475	+	chr10	135106003	+	.	2	5	4726008_1	10.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=CT;MAPQ=60;MATEID=4726008_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_135093001_135118001_111C;SPAN=2528;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:46 GQ:10.7 PL:[10.7, 0.0, 99.8] SR:5 DR:2 LR:-10.64 LO:14.94);ALT=T[chr10:135106003[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135104817	+	chr10	135105899	+	.	19	0	4726011_1	59.0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=4726011_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:135104817(+)-10:135105899(-)__10_135093001_135118001D;SPAN=1082;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:19 DP:20 GQ:5.4 PL:[59.4, 5.4, 0.0] SR:0 DR:19 LR:-59.41 LO:59.41);ALT=C[chr10:135105899[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135113619	+	chr10	135116294	+	.	3	7	4726026_1	18.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=4726026_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_135093001_135118001_13C;SPAN=2675;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:55 GQ:18.2 PL:[18.2, 0.0, 113.9] SR:7 DR:3 LR:-18.11 LO:22.2);ALT=T[chr10:135116294[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135116501	+	chr10	135122322	+	.	30	0	4726101_1	89.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4726101_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:135116501(+)-10:135122322(-)__10_135117501_135142501D;SPAN=5821;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:30 DP:24 GQ:8.1 PL:[89.1, 8.1, 0.0] SR:0 DR:30 LR:-89.12 LO:89.12);ALT=A[chr10:135122322[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135170292	+	chr10	135171458	+	.	13	0	4726164_1	31.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4726164_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:135170292(+)-10:135171458(-)__10_135166501_135191501D;SPAN=1166;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:43 GQ:31.4 PL:[31.4, 0.0, 71.0] SR:0 DR:13 LR:-31.26 LO:32.19);ALT=G[chr10:135171458[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135183582	+	chr10	135186791	+	.	9	0	4726182_1	11.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4726182_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:135183582(+)-10:135186791(-)__10_135166501_135191501D;SPAN=3209;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:67 GQ:11.6 PL:[11.6, 0.0, 150.2] SR:0 DR:9 LR:-11.56 LO:18.68);ALT=C[chr10:135186791[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135184262	+	chr10	135186747	+	.	100	22	4726183_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CACC;MAPQ=60;MATEID=4726183_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_135166501_135191501_260C;SPAN=2485;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:106 DP:68 GQ:28.5 PL:[313.5, 28.5, 0.0] SR:22 DR:100 LR:-313.6 LO:313.6);ALT=C[chr10:135186747[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135207837	+	chr10	135209216	+	.	20	17	4726308_1	63.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=GG;MAPQ=60;MATEID=4726308_2;MATENM=0;NM=0;NUMPARTS=3;REPSEQ=GGG;SCTG=c_10_135191001_135216001_71C;SPAN=1379;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:72 GQ:63.2 PL:[63.2, 0.0, 109.4] SR:17 DR:20 LR:-63.02 LO:63.76);ALT=G[chr10:135209216[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	135207837	+	chr10	135209667	+	GCTGAAGAAGATGCAGAGCAGCCTGAAGCTGGTGGACTGTATCATCGAGGTCCACGATGCCCGG	26	43	4726309_1	99.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=AT;INSERTION=GCTGAAGAAGATGCAGAGCAGCCTGAAGCTGGTGGACTGTATCATCGAGGTCCACGATGCCCGG;MAPQ=60;MATEID=4726309_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_135191001_135216001_71C;SPAN=1830;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:50 DP:71 GQ:23.9 PL:[146.0, 0.0, 23.9] SR:43 DR:26 LR:-150.5 LO:150.5);ALT=G[chr10:135209667[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
