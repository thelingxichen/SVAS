chr4	167669322	+	chr4	167670545	+	.	27	0	2322004_1	75.0	.	DISC_MAPQ=17;EVDNC=DSCRD;IMPRECISE;MAPQ=17;MATEID=2322004_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:167669322(+)-4:167670545(-)__4_167653501_167678501D;SPAN=1223;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:52 GQ:48.8 PL:[75.2, 0.0, 48.8] SR:0 DR:27 LR:-75.28 LO:75.28);ALT=T[chr4:167670545[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	167677048	+	chr4	167683072	+	.	32	16	2322258_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AAGAGATTTGGG;MAPQ=60;MATEID=2322258_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_167678001_167703001_231C;SPAN=6024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:41 DP:33 GQ:10.8 PL:[118.8, 10.8, 0.0] SR:16 DR:32 LR:-118.8 LO:118.8);ALT=G[chr4:167683072[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
