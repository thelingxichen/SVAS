chr10	108030321	+	chr10	108032542	+	.	58	48	4684082_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CTCC;MAPQ=60;MATEID=4684082_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_10_108020501_108045501_127C;SPAN=2221;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:86 DP:21 GQ:23.1 PL:[254.1, 23.1, 0.0] SR:48 DR:58 LR:-254.2 LO:254.2);ALT=C[chr10:108032542[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
