chr7	152281703	+	chr7	152284306	+	.	82	76	5333607_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=CACATGTTTTA;MAPQ=60;MATEID=5333607_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_7_152267501_152292501_401C;SPAN=2603;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:132 DP:40 GQ:35.4 PL:[389.4, 35.4, 0.0] SR:76 DR:82 LR:-389.5 LO:389.5);ALT=A[chr7:152284306[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
