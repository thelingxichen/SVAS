chr2	153103158	-	chr2	153104501	+	.	8	0	1429463_1	0	.	DISC_MAPQ=43;EVDNC=ASDIS;HOMSEQ=TCCTGCCTCAGCCTCCCGAGTAGCTGGGATTACAGG;MAPQ=60;MATEID=1429463_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_153100501_153125501_320C;SPAN=1343;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:138 GQ:10.8 PL:[0.0, 10.8, 356.4] SR:0 DR:8 LR:10.98 LO:13.54);ALT=[chr2:153104501[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
