chr14	31146164	-	chr14	31175535	+	GCA	56	60	8417160_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=GCA;MAPQ=60;MATEID=8417160_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_31139501_31164501_324C;SPAN=29371;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:94 DP:88 GQ:25.2 PL:[277.2, 25.2, 0.0] SR:60 DR:56 LR:-277.3 LO:277.3);ALT=[chr14:31175535[T;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	31165547	+	chr14	31181017	-	TATATATATGCA	25	36	8416614_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TATATATATGCA;MAPQ=60;MATEID=8416614_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_14_31164001_31189001_216C;SPAN=15470;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:57 DP:135 GQ:99 PL:[151.7, 0.0, 174.8] SR:36 DR:25 LR:-151.6 LO:151.7);ALT=T]chr14:31181017];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr14	31746949	-	chr14	31747963	+	.	2	4	8419795_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCCAAAGTGCTGGGATTACAGGCAT;MAPQ=44;MATEID=8419795_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_14_31727501_31752501_323C;SPAN=1014;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:6 DP:146 GQ:19.6 PL:[0.0, 19.6, 392.7] SR:4 DR:2 LR:19.75 LO:9.244);ALT=[chr14:31747963[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr14	32106180	+	chr14	32112024	+	TTTTCTTTTCTTCTCTGTTAG	24	48	8421978_1	72.0	.	DISC_MAPQ=9;EVDNC=ASDIS;INSERTION=TTTTCTTTTCTTCTCTGTTAG;MAPQ=0;MATEID=8421978_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=TTTCTTTTCT;SCTG=c_14_32095001_32120001_29C;SECONDARY;SPAN=5844;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:70 DP:93 GQ:6.5 PL:[72.8, 6.5, 0.0] SR:48 DR:24 LR:-73.62 LO:73.62);ALT=T[chr14:32112024[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
