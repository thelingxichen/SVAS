chr12	2904412	+	chr12	2906302	+	.	0	15	5070198_1	33.0	.	EVDNC=ASSMB;HOMSEQ=AGGT;MAPQ=60;MATEID=5070198_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_12_2891001_2916001_159C;SPAN=1890;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:15 DP:58 GQ:33.8 PL:[33.8, 0.0, 106.4] SR:15 DR:0 LR:-33.8 LO:35.92);ALT=T[chr12:2906302[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr12	2921962	+	chr12	2926385	+	.	13	0	5070726_1	15.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=5070726_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=12:2921962(+)-12:2926385(-)__12_2915501_2940501D;SPAN=4423;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:103 GQ:15.2 PL:[15.2, 0.0, 233.0] SR:0 DR:13 LR:-15.01 LO:26.61);ALT=G[chr12:2926385[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
