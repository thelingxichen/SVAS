chr10	96957656	-	chr10	99459897	+	.	11	0	4669479_1	21.0	.	DISC_MAPQ=15;EVDNC=DSCRD;IMPRECISE;MAPQ=15;MATEID=4669479_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:96957656(-)-10:99459897(-)__10_99445501_99470501D;SPAN=2502241;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:55 GQ:21.5 PL:[21.5, 0.0, 110.6] SR:0 DR:11 LR:-21.41 LO:24.93);ALT=[chr10:99459897[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr10	97028620	+	chr10	97050577	+	.	10	5	4665348_1	30.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=4665348_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_97044501_97069501_7C;SPAN=21957;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:45 GQ:30.8 PL:[30.8, 0.0, 77.0] SR:5 DR:10 LR:-30.72 LO:31.88);ALT=C[chr10:97050577[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	97031542	+	chr10	97050575	+	.	113	78	4665351_1	99.0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=ACC;MAPQ=3;MATEID=4665351_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_97044501_97069501_4C;SPAN=19033;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:156 DP:41 GQ:42.1 PL:[462.1, 42.1, 0.0] SR:78 DR:113 LR:-462.1 LO:462.1);ALT=C[chr10:97050575[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	97208025	+	chr10	97206786	+	.	61	51	4665597_1	99.0	.	DISC_MAPQ=55;EVDNC=ASDIS;HOMSEQ=TGCTC;MAPQ=60;MATEID=4665597_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_97191501_97216501_66C;SPAN=1239;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:96 DP:60 GQ:25.8 PL:[283.8, 25.8, 0.0] SR:51 DR:61 LR:-283.9 LO:283.9);ALT=]chr10:97208025]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr10	97402963	+	chr10	97413047	+	.	0	9	4665927_1	21.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=4665927_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_97387501_97412501_160C;SPAN=10084;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:29 GQ:21.8 PL:[21.8, 0.0, 48.2] SR:9 DR:0 LR:-21.85 LO:22.41);ALT=T[chr10:97413047[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	98469743	+	chr10	98480138	+	.	35	8	4667528_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCTG;MAPQ=60;MATEID=4667528_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_98465501_98490501_252C;SPAN=10395;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:36 DP:51 GQ:16.1 PL:[105.2, 0.0, 16.1] SR:8 DR:35 LR:-108.4 LO:108.4);ALT=G[chr10:98480138[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	99034873	+	chr10	99037398	+	.	62	40	4668584_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=TAAAGCACTG;MAPQ=60;MATEID=4668584_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_99029001_99054001_58C;SPAN=2525;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:81 DP:29 GQ:21.6 PL:[237.6, 21.6, 0.0] SR:40 DR:62 LR:-237.7 LO:237.7);ALT=G[chr10:99037398[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	99201060	+	chr10	99205488	+	.	15	0	4669004_1	42.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4669004_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:99201060(+)-10:99205488(-)__10_99176001_99201001D;SPAN=4428;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:15 DP:5 GQ:3.9 PL:[42.9, 3.9, 0.0] SR:0 DR:15 LR:-42.91 LO:42.91);ALT=T[chr10:99205488[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	99203112	+	chr10	99205710	+	.	22	0	4668886_1	55.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4668886_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:99203112(+)-10:99205710(-)__10_99200501_99225501D;SPAN=2598;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:22 DP:64 GQ:55.4 PL:[55.4, 0.0, 98.3] SR:0 DR:22 LR:-55.28 LO:55.99);ALT=T[chr10:99205710[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	99497078	+	chr10	99498235	+	A	13	11	4669434_1	34.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=A;MAPQ=60;MATEID=4669434_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_99494501_99519501_99C;SPAN=1157;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:80 GQ:34.4 PL:[34.4, 0.0, 159.8] SR:11 DR:13 LR:-34.44 LO:39.04);ALT=G[chr10:99498235[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	100202999	+	chr10	100205057	+	.	2	38	4670705_1	99.0	.	DISC_MAPQ=3;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4670705_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_100205001_100230001_61C;SPAN=2058;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:40 DP:43 GQ:11.4 PL:[125.4, 11.4, 0.0] SR:38 DR:2 LR:-125.4 LO:125.4);ALT=T[chr10:100205057[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	100203052	+	chr10	100206589	+	.	32	0	4670706_1	92.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=4670706_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:100203052(+)-10:100206589(-)__10_100205001_100230001D;SPAN=3537;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:32 DP:25 GQ:8.4 PL:[92.4, 8.4, 0.0] SR:0 DR:32 LR:-92.42 LO:92.42);ALT=C[chr10:100206589[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	100205172	+	chr10	100206564	+	.	30	5	4670707_1	84.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=4670707_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_100205001_100230001_20C;SPAN=1392;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:30 DP:54 GQ:44.9 PL:[84.5, 0.0, 44.9] SR:5 DR:30 LR:-84.98 LO:84.98);ALT=T[chr10:100206564[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
