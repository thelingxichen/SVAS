chr5	46270656	+	chr5	46275837	+	.	0	108	3410418_1	99.0	.	EVDNC=ASSMB;HOMSEQ=TTCT;MAPQ=55;MATEID=3410418_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_46256001_46281001_188C;SPAN=5181;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:108 DP:36 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:108 DR:0 LR:-320.2 LO:320.2);ALT=T[chr5:46275837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
