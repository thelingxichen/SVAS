chr6	55554099	+	chr6	55555112	+	.	22	22	2861140_1	99.0	.	DISC_MAPQ=16;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=2861140_2;MATENM=0;NM=0;NUMPARTS=2;REPSEQ=ATAT;SCTG=c_6_55541501_55566501_6C;SECONDARY;SPAN=1013;SUBN=7;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:55 GQ:18.2 PL:[113.9, 0.0, 18.2] SR:22 DR:22 LR:-117.6 LO:117.6);ALT=A[chr6:55555112[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
