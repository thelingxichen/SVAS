chr2	215728763	+	chr2	215730832	+	.	57	46	1678253_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=TA;MAPQ=60;MATEID=1678253_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_2_215722501_215747501_220C;SPAN=2069;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:89 DP:78 GQ:24 PL:[264.0, 24.0, 0.0] SR:46 DR:57 LR:-264.1 LO:264.1);ALT=A[chr2:215730832[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
