chr4	137144956	+	chr4	137212822	+	.	70	56	2938836_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AT;MAPQ=60;MATEID=2938836_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_4_137200001_137225001_295C;SPAN=67866;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:100 DP:40 GQ:27 PL:[297.0, 27.0, 0.0] SR:56 DR:70 LR:-297.1 LO:297.1);ALT=T[chr4:137212822[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
