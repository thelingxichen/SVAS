chr11	40355317	+	chr11	40356557	-	.	3	2	4834459_1	0	.	DISC_MAPQ=44;EVDNC=ASDIS;HOMSEQ=ACAAAATCCCATGTATTTAT;MAPQ=60;MATEID=4834459_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_40351501_40376501_202C;SPAN=1240;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:4 DP:74 GQ:6.6 PL:[0.0, 6.6, 191.4] SR:2 DR:3 LR:6.844 LO:6.647);ALT=T]chr11:40356557];VARTYPE=BND:INV-hh;JOINTYPE=hh
