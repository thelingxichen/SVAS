chr3	60132754	+	chr3	60204543	+	.	29	22	1439921_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=1439921_2;MATENM=32;NM=0;NUMPARTS=2;SCTG=c_3_60196501_60221501_265C;SPAN=71789;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:47 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:22 DR:29 LR:-137.9 LO:137.9);ALT=T[chr3:60204543[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60341327	+	chr3	60466724	+	.	3	3	1440637_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTTG;MAPQ=60;MATEID=1440637_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_60466001_60491001_251C;SPAN=125397;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:5 DP:58 GQ:0.8 PL:[0.8, 0.0, 139.4] SR:3 DR:3 LR:-0.7914 LO:9.357);ALT=G[chr3:60466724[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	60872125	+	chr3	61013213	+	.	23	24	1442356_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=GC;MAPQ=60;MATEID=1442356_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_61005001_61030001_309C;SPAN=141088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:42 DP:47 GQ:12.6 PL:[138.6, 12.6, 0.0] SR:24 DR:23 LR:-137.9 LO:137.9);ALT=C[chr3:61013213[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	61027818	+	chr3	61237015	+	.	9	0	1443062_1	10.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=1443062_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:61027818(+)-3:61237015(-)__3_61225501_61250501D;SPAN=209197;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:71 GQ:10.7 PL:[10.7, 0.0, 159.2] SR:0 DR:9 LR:-10.47 LO:18.44);ALT=A[chr3:61237015[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
