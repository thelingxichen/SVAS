chr10	1053069	+	chr10	1054896	+	.	0	9	4492540_1	21.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4492540_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_1053501_1078501_86C;SECONDARY;SPAN=1827;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:32 GQ:21.2 PL:[21.2, 0.0, 54.2] SR:9 DR:0 LR:-21.04 LO:21.94);ALT=G[chr10:1054896[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	1090087	+	chr10	1094803	+	.	9	0	4492710_1	10.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4492710_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:1090087(+)-10:1094803(-)__10_1078001_1103001D;SPAN=4716;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:72 GQ:10.4 PL:[10.4, 0.0, 162.2] SR:0 DR:9 LR:-10.2 LO:18.38);ALT=A[chr10:1094803[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	1092494	+	chr10	1093539	+	.	14	0	4492718_1	32.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=4492718_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:1092494(+)-10:1093539(-)__10_1078001_1103001D;SPAN=1045;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:14 DP:51 GQ:32.6 PL:[32.6, 0.0, 88.7] SR:0 DR:14 LR:-32.4 LO:33.96);ALT=C[chr10:1093539[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	1102908	+	chr10	1118054	+	.	12	5	4492734_1	35.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=4492734_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_1078001_1103001_206C;SPAN=15146;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:27 GQ:29 PL:[35.6, 0.0, 29.0] SR:5 DR:12 LR:-35.62 LO:35.62);ALT=G[chr10:1118054[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
