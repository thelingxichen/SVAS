chr5	88100620	+	chr5	88119548	+	.	13	9	2524400_1	55.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TCACCT;MAPQ=60;MATEID=2524400_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_88077501_88102501_179C;SPAN=18928;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:19 DP:28 GQ:12.2 PL:[55.1, 0.0, 12.2] SR:9 DR:13 LR:-56.61 LO:56.61);ALT=T[chr5:88119548[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	88119747	+	chr5	88178772	+	.	0	27	2524533_1	68.0	.	EVDNC=ASSMB;MAPQ=60;MATEID=2524533_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_88175501_88200501_211C;SPAN=59025;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:27 DP:76 GQ:68.6 PL:[68.6, 0.0, 114.8] SR:27 DR:0 LR:-68.54 LO:69.2);ALT=G[chr5:88178772[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
