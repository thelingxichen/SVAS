chr1	222374165	+	chr1	222380540	+	TA	71	34	835227_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;INSERTION=TA;MAPQ=60;MATEID=835227_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_1_222362001_222387001_124C;SPAN=6375;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:92 DP:16 GQ:24.6 PL:[270.6, 24.6, 0.0] SR:34 DR:71 LR:-270.7 LO:270.7);ALT=C[chr1:222380540[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
