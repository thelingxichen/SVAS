chr13	103249555	+	chr13	103257140	+	.	0	12	5626700_1	16.0	.	EVDNC=ASSMB;HOMSEQ=CAGGT;MAPQ=60;MATEID=5626700_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_103243001_103268001_60C;SPAN=7585;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:12 DP:86 GQ:16.4 PL:[16.4, 0.0, 191.3] SR:12 DR:0 LR:-16.31 LO:25.12);ALT=T[chr13:103257140[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	103295727	+	chr13	103296907	+	.	0	5	5626912_1	0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=5626912_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_103292001_103317001_203C;SPAN=1180;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:81 GQ:5.1 PL:[0.0, 5.1, 204.6] SR:5 DR:0 LR:5.44 LO:8.605);ALT=G[chr13:103296907[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	103421940	+	chr13	103426028	+	.	13	0	5627201_1	24.0	.	DISC_MAPQ=57;EVDNC=DSCRD;IMPRECISE;MAPQ=57;MATEID=5627201_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:103421940(+)-13:103426028(-)__13_103414501_103439501D;SPAN=4088;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:13 DP:69 GQ:24.2 PL:[24.2, 0.0, 143.0] SR:0 DR:13 LR:-24.22 LO:29.08);ALT=A[chr13:103426028[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	103504645	+	chr13	103506106	+	.	0	9	5627489_1	7.0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=5627489_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_103488001_103513001_345C;SPAN=1461;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:84 GQ:7.1 PL:[7.1, 0.0, 195.2] SR:9 DR:0 LR:-6.951 LO:17.74);ALT=T[chr13:103506106[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
