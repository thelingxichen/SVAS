chr9	2837402	+	chr9	2838426	+	.	0	6	4126606_1	8.0	.	EVDNC=ASSMB;HOMSEQ=C;MAPQ=60;MATEID=4126606_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_9_2817501_2842501_216C;SPAN=1024;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:43 GQ:8.3 PL:[8.3, 0.0, 94.1] SR:6 DR:0 LR:-8.156 LO:12.56);ALT=C[chr9:2838426[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr9	2837442	+	chr9	2844044	+	.	11	0	4126615_1	27.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4126615_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=9:2837442(+)-9:2844044(-)__9_2842001_2867001D;SPAN=6602;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:34 GQ:27.2 PL:[27.2, 0.0, 53.6] SR:0 DR:11 LR:-27.1 LO:27.63);ALT=C[chr9:2844044[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
