chr10	89096648	+	chr10	89101999	+	.	26	12	4652951_1	80.0	.	DISC_MAPQ=22;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=52;MATEID=4652951_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_89082001_89107001_124C;SPAN=5351;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:29 DP:55 GQ:51.2 PL:[80.9, 0.0, 51.2] SR:12 DR:26 LR:-81.15 LO:81.15);ALT=T[chr10:89101999[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	89700299	+	chr10	89712341	+	GAGATTATACTTTGTGTA	0	49	4653957_1	99.0	.	EVDNC=ASSMB;INSERTION=GAGATTATACTTTGTGTA;MAPQ=60;MATEID=4653957_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_89694501_89719501_123C;SPAN=12042;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:49 DP:19 GQ:13.2 PL:[145.2, 13.2, 0.0] SR:49 DR:0 LR:-145.2 LO:145.2);ALT=A[chr10:89712341[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	90695125	+	chr10	90697818	+	.	0	8	4655269_1	10.0	.	EVDNC=ASSMB;HOMSEQ=CT;MAPQ=60;MATEID=4655269_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_90674501_90699501_216C;SPAN=2693;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:60 GQ:10.1 PL:[10.1, 0.0, 135.5] SR:8 DR:0 LR:-10.15 LO:16.58);ALT=T[chr10:90697818[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	90983589	+	chr10	90984848	+	.	5	7	4655768_1	14.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CCT;MAPQ=60;MATEID=4655768_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_90968501_90993501_146C;SPAN=1259;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:56 GQ:14.6 PL:[14.6, 0.0, 120.2] SR:7 DR:5 LR:-14.54 LO:19.45);ALT=T[chr10:90984848[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	91005599	+	chr10	91011493	+	.	21	0	4655716_1	54.0	.	DISC_MAPQ=60;EVDNC=DSCRD;IMPRECISE;MAPQ=60;MATEID=4655716_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:91005599(+)-10:91011493(-)__10_90993001_91018001D;SPAN=5894;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:21 DP:56 GQ:54.2 PL:[54.2, 0.0, 80.6] SR:0 DR:21 LR:-54.15 LO:54.46);ALT=G[chr10:91011493[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	91007409	+	chr10	91011494	+	.	20	7	4655719_1	63.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTG;MAPQ=60;MATEID=4655719_2;MATENM=0;NM=1;NUMPARTS=2;SCTG=c_10_90993001_91018001_129C;SPAN=4085;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:23 DP:47 GQ:50 PL:[63.2, 0.0, 50.0] SR:7 DR:20 LR:-63.26 LO:63.26);ALT=G[chr10:91011494[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	91461437	+	chr10	91465045	+	.	5	2	4656486_1	1.0	.	DISC_MAPQ=60;EVDNC=TSI_L;HOMSEQ=TTGCAG;MAPQ=60;MATEID=4656486_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_10_91458501_91483501_171C;SPAN=3608;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:6 DP:69 GQ:1.1 PL:[1.1, 0.0, 166.1] SR:2 DR:5 LR:-1.112 LO:11.25);ALT=G[chr10:91465045[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr10	91465199	+	chr10	91468922	+	.	0	9	4656497_1	20.0	.	EVDNC=ASSMB;HOMSEQ=AGG;MAPQ=60;MATEID=4656497_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_91458501_91483501_95C;SPAN=3723;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:36 GQ:20 PL:[20.0, 0.0, 66.2] SR:9 DR:0 LR:-19.96 LO:21.4);ALT=G[chr10:91468922[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
