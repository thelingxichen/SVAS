chr2	192401671	+	chr2	192436215	-	.	33	76	1584835_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=CT;MAPQ=60;MATEID=1584835_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_192398501_192423501_139C;SPAN=34544;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:87 DP:51 GQ:23.4 PL:[257.4, 23.4, 0.0] SR:76 DR:33 LR:-257.5 LO:257.5);ALT=T]chr2:192436215];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr2	192436160	-	chr2	192486430	+	GAAAAAACCCCACAAAATT	19	73	1584895_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;INSERTION=GAAAAAACCCCACAAAATT;MAPQ=60;MATEID=1584895_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_192472001_192497001_14C;SPAN=50270;SUBN=6;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:79 DP:32 GQ:21.3 PL:[234.3, 21.3, 0.0] SR:73 DR:19 LR:-234.4 LO:234.4);ALT=[chr2:192486430[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
