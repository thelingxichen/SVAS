chr2	16407988	+	chr2	16406393	+	CAGGCCC	39	27	923545_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;INSERTION=CAGGCCC;MAPQ=60;MATEID=923545_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_2_16390501_16415501_147C;SPAN=1595;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:54 DP:79 GQ:34.7 PL:[156.8, 0.0, 34.7] SR:27 DR:39 LR:-161.2 LO:161.2);ALT=]chr2:16407988]A;VARTYPE=BND:DUP-th;JOINTYPE=th
chr2	16406433	-	chr2	16407765	+	GAGAGTAGACCCTGAGCCACGTGGGCTTCTAGCAGTTCCCTGGGCCTGCTGGCACCAAGATGGGCTCCC	21	61	923549_1	99.0	.	DISC_MAPQ=33;EVDNC=TSI_L;INSERTION=GAGAGTAGACCCTGAGCCACGTGGGCTTCTAGCAGTTCCCTGGGCCTGCTGGCACCAAGATGGGCTCCC;MAPQ=60;MATEID=923549_2;MATENM=11;NM=3;NUMPARTS=3;REPSEQ=AGAG;SCTG=c_2_16390501_16415501_51C;SPAN=1332;SUBN=3;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:74 DP:85 GQ:16.2 PL:[237.6, 16.2, 0.0] SR:61 DR:21 LR:-239.5 LO:239.5);ALT=[chr2:16407765[C;VARTYPE=BND:INV-tt;JOINTYPE=tt
