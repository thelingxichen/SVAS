chr18	14865661	+	chr18	14864580	+	.	10	0	6552028_1	16.0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6552028_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:14864580(-)-18:14865661(+)__18_14847001_14872001D;SPAN=1081;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:10 DP:62 GQ:16.4 PL:[16.4, 0.0, 131.9] SR:0 DR:10 LR:-16.21 LO:21.62);ALT=]chr18:14865661]T;VARTYPE=BND:DUP-th;JOINTYPE=th
chr18	15194713	+	chr18	15193030	+	.	28	0	6552832_1	76.0	.	DISC_MAPQ=44;EVDNC=DSCRD;IMPRECISE;MAPQ=44;MATEID=6552832_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=18:15193030(-)-18:15194713(+)__18_15190001_15215001D;SPAN=1683;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:28 DP:59 GQ:66.5 PL:[76.4, 0.0, 66.5] SR:0 DR:28 LR:-76.48 LO:76.48);ALT=]chr18:15194713]T;VARTYPE=BND:DUP-th;JOINTYPE=th
