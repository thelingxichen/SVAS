chr3	146385190	+	chr3	146394862	+	.	53	27	2387940_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;HOMSEQ=CA;MAPQ=60;MATEID=2387940_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_3_146387501_146412501_20C;SPAN=9672;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:67 DP:76 GQ:17.1 PL:[217.8, 17.1, 0.0] SR:27 DR:53 LR:-218.2 LO:218.2);ALT=A[chr3:146394862[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	146395165	+	chr3	146390405	+	ATTGGGGAG	0	45	2387947_1	99.0	.	EVDNC=ASSMB;INSERTION=ATTGGGGAG;MAPQ=60;MATEID=2387947_2;MATENM=0;NM=3;NUMPARTS=2;SCTG=c_3_146387501_146412501_5C;SPAN=4760;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:45 DP:126 GQ:99 PL:[114.5, 0.0, 190.4] SR:45 DR:0 LR:-114.4 LO:115.5);ALT=]chr3:146395165]A;VARTYPE=BND:DUP-th;JOINTYPE=th
