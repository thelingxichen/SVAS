chr4	110618960	+	chr4	110624510	+	.	18	0	2143661_1	29.0	.	DISC_MAPQ=56;EVDNC=DSCRD;IMPRECISE;MAPQ=56;MATEID=2143661_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:110618960(+)-4:110624510(-)__4_110617501_110642501D;SPAN=5550;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:18 DP:110 GQ:29.6 PL:[29.6, 0.0, 237.5] SR:0 DR:18 LR:-29.62 LO:39.05);ALT=T[chr4:110624510[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr4	110743646	+	chr4	110745120	+	.	0	6	2144108_1	0	.	EVDNC=ASSMB;HOMSEQ=GGT;MAPQ=60;MATEID=2144108_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_110740001_110765001_159C;SPAN=1474;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:6 DP:122 GQ:12.9 PL:[0.0, 12.9, 320.1] SR:6 DR:0 LR:13.25 LO:9.719);ALT=T[chr4:110745120[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
