chr13	77566407	+	chr13	77570036	+	CGCTTTGACTTCCGTCCAAAACCTGATCCTTATTGTCAAGCTAAGTATACTTTCTGTCCAACTGGCTCACCTATCCCAGTTATGGAGGGTGATGATGACATTGAAGTTTTTCGATTACAAGCCCCAGTATGGGAATTTAAATATGGAGACCTCCTGGGACACTT	7	18	5561911_1	54.0	.	DISC_MAPQ=60;EVDNC=TSI_G;HOMSEQ=G;INSERTION=CGCTTTGACTTCCGTCCAAAACCTGATCCTTATTGTCAAGCTAAGTATACTTTCTGTCCAACTGGCTCACCTATCCCAGTTATGGAGGGTGATGATGACATTGAAGTTTTTCGATTACAAGCCCCAGTATGGGAATTTAAATATGGAGACCTCCTGGGACACTT;MAPQ=60;MATEID=5561911_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_77542501_77567501_72C;SPAN=3629;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:20 DP:44 GQ:50.9 PL:[54.2, 0.0, 50.9] SR:18 DR:7 LR:-54.1 LO:54.1);ALT=G[chr13:77570036[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	77566407	+	chr13	77569198	+	.	23	7	5561910_1	70.0	.	DISC_MAPQ=58;EVDNC=TSI_L;HOMSEQ=G;MAPQ=60;MATEID=5561910_2;MATENM=0;NM=0;NUMPARTS=3;SCTG=c_13_77542501_77567501_72C;SPAN=2791;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:25 DP:44 GQ:34.4 PL:[70.7, 0.0, 34.4] SR:7 DR:23 LR:-71.2 LO:71.2);ALT=G[chr13:77569198[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	77844675	+	chr13	77847605	+	.	5	6	5562568_1	4.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=ACCT;MAPQ=60;MATEID=5562568_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_77836501_77861501_125C;SPAN=2930;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:7 DP:70 GQ:4.1 PL:[4.1, 0.0, 165.8] SR:6 DR:5 LR:-4.142 LO:13.57);ALT=T[chr13:77847605[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	78764969	+	chr13	78767837	+	.	34	29	5565009_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=C;MAPQ=60;MATEID=5565009_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_13_78767501_78792501_113C;SPAN=2868;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:53 DP:36 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:29 DR:34 LR:-155.1 LO:155.1);ALT=C[chr13:78767837[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	78997624	+	chr13	78998720	+	.	38	25	5565570_1	99.0	.	DISC_MAPQ=47;EVDNC=ASDIS;HOMSEQ=AACATGGTGAAACCC;MAPQ=60;MATEID=5565570_2;MATENM=1;NM=1;NUMPARTS=2;SCTG=c_13_78988001_79013001_355C;SPAN=1096;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:51 DP:68 GQ:14.6 PL:[149.9, 0.0, 14.6] SR:25 DR:38 LR:-156.4 LO:156.4);ALT=C[chr13:78998720[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr13	79747137	-	chr13	79748295	+	.	9	0	5567511_1	18.0	.	DISC_MAPQ=53;EVDNC=DSCRD;IMPRECISE;MAPQ=53;MATEID=5567511_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=13:79747137(-)-13:79748295(-)__13_79723001_79748001D;SPAN=1158;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:42 GQ:18.5 PL:[18.5, 0.0, 81.2] SR:0 DR:9 LR:-18.33 LO:20.7);ALT=[chr13:79748295[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
