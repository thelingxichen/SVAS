chr16	84501438	+	chr16	84504116	+	CAGCTGCCCCAGGATGGACC	0	46	9445019_1	99.0	.	EVDNC=ASSMB;INSERTION=CAGCTGCCCCAGGATGGACC;MAPQ=60;MATEID=9445019_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_16_84500501_84525501_175C;SPAN=2678;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:46 DP:22 GQ:12.3 PL:[135.3, 12.3, 0.0] SR:46 DR:0 LR:-135.3 LO:135.3);ALT=C[chr16:84504116[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
