chr3	196318448	+	chr11	45399421	-	.	29	41	6780345_1	99.0	.	DISC_MAPQ=56;EVDNC=ASDIS;HOMSEQ=GTGCCTGTAATCCCAGCTACT;MAPQ=44;MATEID=6780345_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_45398501_45423501_120C;SPAN=-1;SUBN=5;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:68 DP:75 GQ:20.1 PL:[221.1, 20.1, 0.0] SR:41 DR:29 LR:-221.2 LO:221.2);ALT=T]chr11:45399421];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr3	196318494	-	chr11	45399307	+	.	29	55	2595197_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;HOMSEQ=CTCTGTCACCCAGGCTGGAGTGCAATGGCGCGATCTCGGCTCACTGCAA;MAPQ=60;MATEID=2595197_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_3_196318501_196343501_116C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:83 DP:23 GQ:22.2 PL:[244.2, 22.2, 0.0] SR:55 DR:29 LR:-244.3 LO:244.3);ALT=[chr11:45399307[T;VARTYPE=BND:TRX-tt;JOINTYPE=tt
chr3	196530024	+	chr15	21937518	-	.	8	0	8769422_1	0	.	DISC_MAPQ=22;EVDNC=DSCRD;IMPRECISE;MAPQ=22;MATEID=8769422_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:196530024(+)-15:21937518(+)__15_21927501_21952501D;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:307 GQ:56.6 PL:[0.0, 56.6, 858.2] SR:0 DR:8 LR:56.77 LO:10.73);ALT=T]chr15:21937518];VARTYPE=BND:TRX-hh;JOINTYPE=hh
chr11	45429849	+	chr11	45431614	+	.	56	36	6780297_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=GCC;MAPQ=60;MATEID=6780297_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_11_45423001_45448001_360C;SPAN=1765;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:84 DP:72 GQ:22.5 PL:[247.5, 22.5, 0.0] SR:36 DR:56 LR:-247.6 LO:247.6);ALT=C[chr11:45431614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr15	22336853	+	chr15	22344094	+	A	209	79	8772818_1	99.0	.	DISC_MAPQ=255;EVDNC=ASDIS;INSERTION=A;MAPQ=47;MATEID=8772818_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_15_22344001_22369001_297C;SPAN=7241;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:241 DP:39 GQ:64.9 PL:[712.9, 64.9, 0.0] SR:79 DR:209 LR:-713.0 LO:713.0);ALT=T[chr15:22344094[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
