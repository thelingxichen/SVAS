chr4	58621414	+	chr4	59443105	-	.	21	0	2727993_1	59.0	.	DISC_MAPQ=42;EVDNC=DSCRD;IMPRECISE;MAPQ=42;MATEID=2727993_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:58621414(+)-4:59443105(+)__4_59437001_59462001D;SPAN=821691;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:21 DP:37 GQ:29.6 PL:[59.3, 0.0, 29.6] SR:0 DR:21 LR:-59.79 LO:59.79);ALT=A]chr4:59443105];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr4	58621621	-	chr4	59442908	+	.	14	0	2727994_1	29.0	.	DISC_MAPQ=16;EVDNC=DSCRD;IMPRECISE;MAPQ=16;MATEID=2727994_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=4:58621621(-)-4:59442908(-)__4_59437001_59462001D;SPAN=821287;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:14 DP:61 GQ:29.9 PL:[29.9, 0.0, 115.7] SR:0 DR:14 LR:-29.69 LO:32.68);ALT=[chr4:59442908[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr4	58887276	+	chr4	58888335	+	TCTAGAGACTTT	80	56	2727325_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCTAGAGACTTT;MAPQ=60;MATEID=2727325_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_58873501_58898501_82C;SPAN=1059;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:108 DP:50 GQ:29.1 PL:[320.1, 29.1, 0.0] SR:56 DR:80 LR:-320.2 LO:320.2);ALT=A[chr4:58888335[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
