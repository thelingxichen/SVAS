chrX	33831103	+	chrX	22263700	+	.	4	4	11063848_1	1.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CTTCT;MAPQ=60;MATEID=11063848_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_23_33810001_33835001_123C;SPAN=11567403;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:5 DP:57 GQ:1.1 PL:[1.1, 0.0, 136.4] SR:4 DR:4 LR:-1.062 LO:9.396);ALT=]chrX:33831103]C;VARTYPE=BND:DUP-th;JOINTYPE=th
