chr2	33091738	+	chr2	33095624	+	.	31	25	744505_1	99.0	.	DISC_MAPQ=54;EVDNC=ASDIS;HOMSEQ=ATGGAATATTT;MAPQ=60;MATEID=744505_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_33075001_33100001_45C;SPAN=3886;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:50 DP:23 GQ:13.5 PL:[148.5, 13.5, 0.0] SR:25 DR:31 LR:-148.5 LO:148.5);ALT=T[chr2:33095624[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	33224462	+	chr2	33227293	+	.	53	37	744309_1	99.0	.	DISC_MAPQ=58;EVDNC=ASDIS;MAPQ=60;MATEID=744309_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_33222001_33247001_79C;SPAN=2831;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:76 DP:44 GQ:20.4 PL:[224.4, 20.4, 0.0] SR:37 DR:53 LR:-224.5 LO:224.5);ALT=A[chr2:33227293[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	33334387	+	chr2	33335653	+	TCACTCCAGCCTCAA	4	3	744569_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=TCACTCCAGCCTCAA;MAPQ=60;MATEID=744569_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_33320001_33345001_253C;SPAN=1266;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/0 AD:5 DP:71 GQ:2.4 PL:[0.0, 2.4, 174.9] SR:3 DR:4 LR:2.731 LO:8.9);ALT=T[chr2:33335653[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	33740273	+	chr2	33741608	+	.	0	9	745760_1	9.0	.	EVDNC=ASSMB;HOMSEQ=G;MAPQ=60;MATEID=745760_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_2_33736501_33761501_342C;SPAN=1335;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:9 DP:76 GQ:9.2 PL:[9.2, 0.0, 174.2] SR:9 DR:0 LR:-9.119 LO:18.15);ALT=G[chr2:33741608[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	34695829	+	chr2	34736568	+	GTAGGGGT	82	60	747955_1	99.0	.	DISC_MAPQ=45;EVDNC=ASDIS;INSERTION=GTAGGGGT;MAPQ=60;MATEID=747955_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_34716501_34741501_7C;SPAN=40739;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:113 DP:18 GQ:30.3 PL:[333.3, 30.3, 0.0] SR:60 DR:82 LR:-333.4 LO:333.4);ALT=T[chr2:34736568[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr2	34965729	+	chr2	34967270	+	AACAG	32	15	748654_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;INSERTION=AACAG;MAPQ=60;MATEID=748654_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_2_34961501_34986501_279C;SPAN=1541;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:39 DP:53 GQ:12.2 PL:[114.5, 0.0, 12.2] SR:15 DR:32 LR:-118.9 LO:118.9);ALT=A[chr2:34967270[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
