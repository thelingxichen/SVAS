chr15	20581504	+	chr15	20589614	+	.	75	35	5887925_1	99.0	.	DISC_MAPQ=30;EVDNC=ASDIS;HOMSEQ=AATACTATGCAGCCATAAGAAAGGATGAGTTCATGTCCTTTG;MAPQ=60;MATEID=5887925_2;MATENM=0;NM=2;NUMPARTS=2;SCTG=c_15_20580001_20605001_372C;SPAN=8110;SUBN=1;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:1/1 AD:101 DP:91 GQ:27 PL:[297.0, 27.0, 0.0] SR:35 DR:75 LR:-297.1 LO:297.1);ALT=G[chr15:20589614[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
