chr4	24578302	+	chr4	24585945	+	.	10	10	1923264_1	39.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=CC;MAPQ=60;MATEID=1923264_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_24573501_24598501_17C;SPAN=7643;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:17 DP:62 GQ:39.5 PL:[39.5, 0.0, 108.8] SR:10 DR:10 LR:-39.32 LO:41.22);ALT=C[chr4:24585945[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
