chr7	52397548	+	chr7	52171280	+	.	11	0	3308848_1	20.0	.	DISC_MAPQ=29;EVDNC=DSCRD;IMPRECISE;MAPQ=29;MATEID=3308848_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:52171280(-)-7:52397548(+)__7_52381001_52406001D;SPAN=226268;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:11 DP:57 GQ:20.9 PL:[20.9, 0.0, 116.6] SR:0 DR:11 LR:-20.87 LO:24.74);ALT=]chr7:52397548]A;VARTYPE=BND:DUP-th;JOINTYPE=th
