chr5	167915741	+	chr5	167919662	+	.	0	8	2637751_1	12.0	.	EVDNC=ASSMB;HOMSEQ=AG;MAPQ=60;MATEID=2637751_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_167898501_167923501_168C;SPAN=3921;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:8 DP:53 GQ:12.2 PL:[12.2, 0.0, 114.5] SR:8 DR:0 LR:-12.05 LO:17.05);ALT=G[chr5:167919662[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr5	167945068	+	chr5	167946085	+	.	0	4	2637803_1	2.0	.	EVDNC=ASSMB;HOMSEQ=GG;MAPQ=60;MATEID=2637803_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_5_167923001_167948001_45C;SPAN=1017;SVTYPE=BND;TOOL=svaba;GENOTYPE=colo829(GT:0/1 AD:4 DP:41 GQ:2.3 PL:[2.3, 0.0, 94.7] SR:4 DR:0 LR:-2.096 LO:7.711);ALT=G[chr5:167946085[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
