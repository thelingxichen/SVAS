chr10	1487730	+	chr10	1486195	+	.	86	1	6061979_1	99.0	.	DISC_MAPQ=52;EVDNC=ASDIS;HOMSEQ=TCTGTCCAT;MAPQ=2;MATEID=6061979_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_10_1470001_1495001_55C;SPAN=1535;SUBN=2;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:86 DP:107 GQ:4.1 PL:[254.9, 0.0, 4.1] SR:1 DR:86 LR:-269.6 LO:269.6);ALT=]chr10:1487730]T;VARTYPE=BND:DUP-th;JOINTYPE=th
