chr10	109273966	+	chr10	109277346	-	.	4	5	6510506_1	0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=6510506_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_109270001_109295001_417C;SPAN=3380;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:136 GQ:10.2 PL:[0.0, 10.2, 349.8] SR:5 DR:4 LR:10.44 LO:13.6);ALT=A]chr10:109277346];VARTYPE=BND:INV-hh;JOINTYPE=hh
chr10	109273971	+	chr10	109277262	+	.	0	8	6510507_1	0	.	EVDNC=ASSMB;MAPQ=60;MATEID=6510507_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_10_109270001_109295001_217C;SPAN=3291;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:8 DP:136 GQ:10.2 PL:[0.0, 10.2, 349.8] SR:8 DR:0 LR:10.44 LO:13.6);ALT=A[chr10:109277262[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
