chr10	46961047	+	chr10	46963026	-	.	9	0	6236297_1	0	.	DISC_MAPQ=25;EVDNC=DSCRD;IMPRECISE;MAPQ=25;MATEID=6236297_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=10:46961047(+)-10:46963026(+)__10_46942001_46967001D;SPAN=1979;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:9 DP:317 GQ:56 PL:[0.0, 56.0, 881.3] SR:0 DR:9 LR:56.17 LO:12.41);ALT=T]chr10:46963026];VARTYPE=BND:INV-hh;JOINTYPE=hh
