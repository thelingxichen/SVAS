chr7	47104654	+	chr7	47102859	+	.	11	0	4776515_1	0	.	DISC_MAPQ=58;EVDNC=DSCRD;IMPRECISE;MAPQ=58;MATEID=4776515_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=7:47102859(-)-7:47104654(+)__7_47089001_47114001D;SPAN=1795;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:11 DP:161 GQ:7 PL:[0.0, 7.0, 402.6] SR:0 DR:11 LR:7.308 LO:19.43);ALT=]chr7:47104654]T;VARTYPE=BND:DUP-th;JOINTYPE=th
