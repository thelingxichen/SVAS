chr4	22523077	+	chr4	22437123	+	.	69	64	2653893_1	99.0	.	DISC_MAPQ=59;EVDNC=ASDIS;HOMSEQ=AG;MAPQ=60;MATEID=2653893_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_4_22515501_22540501_118C;SPAN=85954;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:111 DP:41 GQ:29.7 PL:[326.7, 29.7, 0.0] SR:64 DR:69 LR:-326.8 LO:326.8);ALT=]chr4:22523077]A;VARTYPE=BND:DUP-th;JOINTYPE=th
