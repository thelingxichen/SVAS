chr3	113577328	-	chr3	113579541	+	.	10	0	2250387_1	0	.	DISC_MAPQ=54;EVDNC=DSCRD;IMPRECISE;MAPQ=54;MATEID=2250387_2;MATENM=-1;NM=-1;NUMPARTS=0;SCTG=3:113577328(-)-3:113579541(-)__3_113557501_113582501D;SPAN=2213;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/0 AD:10 DP:196 GQ:19.9 PL:[0.0, 19.9, 514.9] SR:0 DR:10 LR:20.09 LO:16.36);ALT=[chr3:113579541[A;VARTYPE=BND:INV-tt;JOINTYPE=tt
chr3	114146389	+	chr3	114279002	+	.	7	7	2252629_1	17.0	.	DISC_MAPQ=60;EVDNC=ASDIS;MAPQ=60;MATEID=2252629_2;MATENM=0;NM=0;NUMPARTS=2;SCTG=c_3_114145501_114170501_158C;SPAN=132613;SUBN=8;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:0/1 AD:11 DP:71 GQ:17.3 PL:[17.3, 0.0, 152.6] SR:7 DR:7 LR:-17.08 LO:23.58);ALT=G[chr3:114279002[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
chr3	114472276	+	chr13	58340088	-	.	14	45	2253783_1	99.0	.	DISC_MAPQ=42;EVDNC=ASDIS;HOMSEQ=TATATATATACACACACGTATATATATATATATA;MAPQ=60;MATEID=2253783_2;MATENM=1;NM=0;NUMPARTS=2;SCTG=c_3_114464001_114489001_30C;SPAN=-1;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:53 DP:43 GQ:14.1 PL:[155.1, 14.1, 0.0] SR:45 DR:14 LR:-155.1 LO:155.1);ALT=A]chr13:58340088];VARTYPE=BND:TRX-hh;JOINTYPE=hh
