chr1	116229486	+	chr1	116232841	+	.	48	60	465957_1	99.0	.	DISC_MAPQ=60;EVDNC=ASDIS;HOMSEQ=TTG;MAPQ=60;MATEID=465957_2;MATENM=2;NM=0;NUMPARTS=2;SCTG=c_1_116228001_116253001_152C;SPAN=3355;SVTYPE=BND;TOOL=svaba;GENOTYPE=mkn45(GT:1/1 AD:93 DP:24 GQ:24.9 PL:[273.9, 24.9, 0.0] SR:60 DR:48 LR:-274.0 LO:274.0);ALT=G[chr1:116232841[;VARTYPE=BND:DEL-ht;JOINTYPE=ht
